* NGSPICE file created from phoeniX.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 Q CLK D gnd vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

.subckt phoeniX vdd gnd CLK reset instruction_memory_interface_data[0] instruction_memory_interface_data[1]
+ instruction_memory_interface_data[2] instruction_memory_interface_data[3] instruction_memory_interface_data[4]
+ instruction_memory_interface_data[5] instruction_memory_interface_data[6] instruction_memory_interface_data[7]
+ instruction_memory_interface_data[8] instruction_memory_interface_data[9] instruction_memory_interface_data[10]
+ instruction_memory_interface_data[11] instruction_memory_interface_data[12] instruction_memory_interface_data[13]
+ instruction_memory_interface_data[14] instruction_memory_interface_data[15] instruction_memory_interface_data[16]
+ instruction_memory_interface_data[17] instruction_memory_interface_data[18] instruction_memory_interface_data[19]
+ instruction_memory_interface_data[20] instruction_memory_interface_data[21] instruction_memory_interface_data[22]
+ instruction_memory_interface_data[23] instruction_memory_interface_data[24] instruction_memory_interface_data[25]
+ instruction_memory_interface_data[26] instruction_memory_interface_data[27] instruction_memory_interface_data[28]
+ instruction_memory_interface_data[29] instruction_memory_interface_data[30] instruction_memory_interface_data[31]
+ data_memory_interface_data[0] data_memory_interface_data[1] data_memory_interface_data[2]
+ data_memory_interface_data[3] data_memory_interface_data[4] data_memory_interface_data[5]
+ data_memory_interface_data[6] data_memory_interface_data[7] data_memory_interface_data[8]
+ data_memory_interface_data[9] data_memory_interface_data[10] data_memory_interface_data[11]
+ data_memory_interface_data[12] data_memory_interface_data[13] data_memory_interface_data[14]
+ data_memory_interface_data[15] data_memory_interface_data[16] data_memory_interface_data[17]
+ data_memory_interface_data[18] data_memory_interface_data[19] data_memory_interface_data[20]
+ data_memory_interface_data[21] data_memory_interface_data[22] data_memory_interface_data[23]
+ data_memory_interface_data[24] data_memory_interface_data[25] data_memory_interface_data[26]
+ data_memory_interface_data[27] data_memory_interface_data[28] data_memory_interface_data[29]
+ data_memory_interface_data[30] data_memory_interface_data[31] instruction_memory_interface_enable
+ instruction_memory_interface_state instruction_memory_interface_address[0] instruction_memory_interface_address[1]
+ instruction_memory_interface_address[2] instruction_memory_interface_address[3]
+ instruction_memory_interface_address[4] instruction_memory_interface_address[5]
+ instruction_memory_interface_address[6] instruction_memory_interface_address[7]
+ instruction_memory_interface_address[8] instruction_memory_interface_address[9]
+ instruction_memory_interface_address[10] instruction_memory_interface_address[11]
+ instruction_memory_interface_address[12] instruction_memory_interface_address[13]
+ instruction_memory_interface_address[14] instruction_memory_interface_address[15]
+ instruction_memory_interface_address[16] instruction_memory_interface_address[17]
+ instruction_memory_interface_address[18] instruction_memory_interface_address[19]
+ instruction_memory_interface_address[20] instruction_memory_interface_address[21]
+ instruction_memory_interface_address[22] instruction_memory_interface_address[23]
+ instruction_memory_interface_address[24] instruction_memory_interface_address[25]
+ instruction_memory_interface_address[26] instruction_memory_interface_address[27]
+ instruction_memory_interface_address[28] instruction_memory_interface_address[29]
+ instruction_memory_interface_address[30] instruction_memory_interface_address[31]
+ instruction_memory_interface_frame_mask[0] instruction_memory_interface_frame_mask[1]
+ instruction_memory_interface_frame_mask[2] instruction_memory_interface_frame_mask[3]
+ data_memory_interface_enable data_memory_interface_state data_memory_interface_address[0]
+ data_memory_interface_address[1] data_memory_interface_address[2] data_memory_interface_address[3]
+ data_memory_interface_address[4] data_memory_interface_address[5] data_memory_interface_address[6]
+ data_memory_interface_address[7] data_memory_interface_address[8] data_memory_interface_address[9]
+ data_memory_interface_address[10] data_memory_interface_address[11] data_memory_interface_address[12]
+ data_memory_interface_address[13] data_memory_interface_address[14] data_memory_interface_address[15]
+ data_memory_interface_address[16] data_memory_interface_address[17] data_memory_interface_address[18]
+ data_memory_interface_address[19] data_memory_interface_address[20] data_memory_interface_address[21]
+ data_memory_interface_address[22] data_memory_interface_address[23] data_memory_interface_address[24]
+ data_memory_interface_address[25] data_memory_interface_address[26] data_memory_interface_address[27]
+ data_memory_interface_address[28] data_memory_interface_address[29] data_memory_interface_address[30]
+ data_memory_interface_address[31] data_memory_interface_frame_mask[0] data_memory_interface_frame_mask[1]
+ data_memory_interface_frame_mask[2] data_memory_interface_frame_mask[3]
XFILL_9_6_0 gnd vdd FILL
XNAND2X1_580 INVX8_5/A MUX2X1_47/A gnd NAND2X1_580/Y vdd NAND2X1
XNAND2X1_591 AND2X2_56/B INVX2_55/A gnd OAI22X1_40/B vdd NAND2X1
XFILL_17_5_0 gnd vdd FILL
XFILL_41_3_0 gnd vdd FILL
XINVX1_402 INVX1_402/A gnd INVX1_402/Y vdd INVX1
XOAI21X1_360 INVX8_8/A INVX2_30/A NAND2X1_338/Y gnd OAI21X1_410/A vdd OAI21X1
XOAI21X1_371 NOR2X1_1/A AND2X2_25/Y OR2X2_44/B gnd OAI21X1_371/Y vdd OAI21X1
XOAI21X1_382 OR2X2_25/Y INVX8_5/A OAI21X1_381/Y gnd NOR2X1_223/B vdd OAI21X1
XAND2X2_5 AND2X2_5/A AND2X2_5/B gnd AND2X2_5/Y vdd AND2X2
XOAI21X1_393 BUFX4_39/Y NOR2X1_151/B OAI21X1_393/C gnd OAI21X1_393/Y vdd OAI21X1
XINVX1_413 INVX1_413/A gnd INVX1_413/Y vdd INVX1
XINVX1_424 INVX1_424/A gnd INVX1_424/Y vdd INVX1
XINVX1_435 INVX1_435/A gnd INVX1_435/Y vdd INVX1
XINVX1_468 BUFX2_39/A gnd INVX1_468/Y vdd INVX1
XINVX1_457 INVX1_457/A gnd INVX1_457/Y vdd INVX1
XINVX1_446 OR2X2_59/B gnd INVX1_446/Y vdd INVX1
XINVX1_479 BUFX2_56/A gnd INVX1_479/Y vdd INVX1
XFILL_32_3_0 gnd vdd FILL
XFILL_23_3_0 gnd vdd FILL
XFILL_6_4_0 gnd vdd FILL
XMUX2X1_17 INVX1_242/A INVX2_85/A INVX4_4/A gnd MUX2X1_17/Y vdd MUX2X1
XMUX2X1_39 MUX2X1_39/A INVX2_53/A INVX8_8/A gnd MUX2X1_43/B vdd MUX2X1
XMUX2X1_28 MUX2X1_28/A MUX2X1_28/B INVX8_4/A gnd MUX2X1_28/Y vdd MUX2X1
XFILL_14_3_0 gnd vdd FILL
XOAI21X1_190 BUFX4_13/Y BUFX4_196/Y OAI21X1_865/Y gnd NAND3X1_65/C vdd OAI21X1
XINVX1_210 INVX1_210/A gnd INVX1_210/Y vdd INVX1
XINVX1_243 INVX1_243/A gnd INVX1_243/Y vdd INVX1
XINVX1_232 NOR2X1_1/A gnd INVX1_232/Y vdd INVX1
XINVX1_221 INVX1_221/A gnd INVX1_221/Y vdd INVX1
XINVX1_254 MUX2X1_9/A gnd INVX1_254/Y vdd INVX1
XINVX1_265 OR2X2_10/Y gnd INVX1_265/Y vdd INVX1
XINVX1_276 INVX1_276/A gnd INVX1_276/Y vdd INVX1
XINVX1_287 INVX1_287/A gnd INVX1_287/Y vdd INVX1
XINVX1_298 AND2X2_19/Y gnd INVX1_298/Y vdd INVX1
XNAND2X1_21 BUFX4_18/Y NAND2X1_21/B gnd OAI21X1_21/C vdd NAND2X1
XNAND2X1_10 BUFX4_20/Y NAND2X1_10/B gnd OAI21X1_10/C vdd NAND2X1
XNAND2X1_32 BUFX4_20/Y NAND2X1_32/B gnd OAI21X1_32/C vdd NAND2X1
XNAND2X1_43 BUFX4_30/Y NAND2X1_43/B gnd OAI21X1_43/C vdd NAND2X1
XNAND2X1_76 INVX1_253/A BUFX4_163/Y gnd NAND2X1_76/Y vdd NAND2X1
XNAND2X1_65 NOR2X1_6/A NOR2X1_6/B gnd OR2X2_1/A vdd NAND2X1
XNAND2X1_54 BUFX4_30/Y NAND2X1_54/B gnd NAND2X1_54/Y vdd NAND2X1
XNAND2X1_98 NAND2X1_98/A BUFX4_156/Y gnd NAND2X1_98/Y vdd NAND2X1
XNAND2X1_87 INVX1_271/A BUFX4_158/Y gnd NAND2X1_87/Y vdd NAND2X1
XFILL_35_1 gnd vdd FILL
XAOI21X1_225 INVX1_495/A INVX1_567/Y AOI21X1_225/C gnd NAND3X1_254/C vdd AOI21X1
XAOI21X1_203 INVX1_426/Y AOI21X1_203/B INVX1_427/A gnd NOR2X1_366/B vdd AOI21X1
XAOI21X1_214 OAI21X1_773/C AND2X2_69/A INVX2_28/A gnd OAI21X1_783/A vdd AOI21X1
XAOI21X1_236 NAND2X1_962/Y NOR2X1_435/Y NOR2X1_436/Y gnd AOI21X1_236/Y vdd AOI21X1
XAOI21X1_247 AND2X2_95/Y OAI21X1_928/Y OAI21X1_930/Y gnd AOI21X1_247/Y vdd AOI21X1
XAOI21X1_258 AOI21X1_263/A AOI21X1_258/B OAI22X1_54/Y gnd OAI21X1_986/A vdd AOI21X1
XAOI21X1_269 INVX1_759/A NOR2X1_475/Y BUFX2_36/A gnd AOI21X1_271/B vdd AOI21X1
XAOI22X1_30 AOI22X1_30/A BUFX4_236/Y BUFX4_256/Y AOI22X1_30/D gnd AOI22X1_30/Y vdd
+ AOI22X1
XAOI22X1_41 NOR2X1_15/Y NOR2X1_14/Y NOR2X1_18/Y INVX1_229/A gnd AOI22X1_41/Y vdd AOI22X1
XAOI22X1_74 AOI22X1_74/A AOI21X1_98/A AOI22X1_74/C AOI22X1_85/B gnd NAND3X1_91/C vdd
+ AOI22X1
XAOI22X1_52 MUX2X1_3/A BUFX4_235/Y BUFX4_151/Y MUX2X1_3/B gnd NOR2X1_40/B vdd AOI22X1
XAOI22X1_63 AOI22X1_63/A BUFX4_233/Y AND2X2_11/A OR2X2_55/A gnd NOR2X1_55/B vdd AOI22X1
XAOI22X1_96 AOI22X1_96/A AOI22X1_96/B AOI22X1_96/C AOI22X1_96/D gnd AOI22X1_96/Y vdd
+ AOI22X1
XAOI22X1_85 BUFX4_190/Y AOI22X1_85/B NOR2X1_232/A BUFX4_154/Y gnd AOI22X1_85/Y vdd
+ AOI22X1
XNAND3X1_229 BUFX4_221/Y NAND3X1_228/Y NAND3X1_229/C gnd NAND2X1_768/B vdd NAND3X1
XNAND3X1_207 BUFX4_218/Y NAND3X1_207/B NAND3X1_207/C gnd NAND2X1_735/B vdd NAND3X1
XNAND3X1_218 INVX1_532/Y BUFX4_207/Y BUFX4_34/Y gnd NAND3X1_218/Y vdd NAND3X1
XOAI22X1_3 INVX2_3/Y BUFX2_91/A INVX2_1/A INVX1_132/Y gnd NOR3X1_16/B vdd OAI22X1
XFILL_30_6_1 gnd vdd FILL
XDFFPOSX1_328 INVX1_279/A CLKBUF1_25/Y OAI21X1_896/Y gnd vdd DFFPOSX1
XDFFPOSX1_317 INVX2_12/A CLKBUF1_56/Y OAI21X1_885/Y gnd vdd DFFPOSX1
XDFFPOSX1_306 INVX2_7/A CLKBUF1_34/Y OAI21X1_879/Y gnd vdd DFFPOSX1
XDFFPOSX1_339 XOR2X1_1/A CLKBUF1_9/Y NOR2X1_22/A gnd vdd DFFPOSX1
XNAND2X1_409 BUFX4_213/Y NAND2X1_409/B gnd INVX1_389/A vdd NAND2X1
XFILL_37_2_0 gnd vdd FILL
XFILL_38_7_1 gnd vdd FILL
XNOR2X1_420 INVX1_467/A INVX1_664/Y gnd NOR2X1_422/A vdd NOR2X1
XNOR2X1_442 NOR2X1_442/A NOR2X1_442/B gnd NOR2X1_442/Y vdd NOR2X1
XNOR2X1_431 MUX2X1_9/B INVX2_84/Y gnd NOR2X1_431/Y vdd NOR2X1
XNOR2X1_475 NOR2X1_475/A NOR2X1_475/B gnd NOR2X1_475/Y vdd NOR2X1
XNOR2X1_464 OR2X2_59/A OR2X2_59/B gnd OAI22X1_52/D vdd NOR2X1
XNOR2X1_453 OR2X2_53/B INVX1_704/Y gnd NOR2X1_453/Y vdd NOR2X1
XNOR2X1_486 INVX2_88/A NOR3X1_73/B gnd BUFX4_253/A vdd NOR2X1
XFILL_20_1_0 gnd vdd FILL
XOAI21X1_904 INVX1_700/A INVX1_671/Y NAND2X1_939/Y gnd NOR2X1_425/B vdd OAI21X1
XFILL_21_6_1 gnd vdd FILL
XOAI21X1_915 INVX1_306/A INVX2_81/Y AND2X2_82/B gnd NOR3X1_71/C vdd OAI21X1
XOAI21X1_948 NOR2X1_487/A NOR3X1_78/C INVX1_756/A gnd BUFX2_33/A vdd OAI21X1
XOAI21X1_926 NOR2X1_457/Y NOR2X1_458/Y INVX1_684/A gnd AOI21X1_246/B vdd OAI21X1
XOAI21X1_937 AOI21X1_250/Y OAI21X1_938/A OAI21X1_937/C gnd OR2X2_67/A vdd OAI21X1
XOAI21X1_959 INVX4_14/Y INVX1_721/Y OAI21X1_959/C gnd OAI21X1_959/Y vdd OAI21X1
XINVX2_12 INVX2_12/A gnd INVX2_12/Y vdd INVX2
XINVX2_34 INVX2_34/A gnd INVX2_34/Y vdd INVX2
XINVX2_45 INVX2_45/A gnd INVX2_45/Y vdd INVX2
XINVX2_23 INVX2_23/A gnd INVX2_23/Y vdd INVX2
XNAND2X1_921 NOR2X1_22/A NOR2X1_411/Y gnd NAND2X1_921/Y vdd NAND2X1
XNAND2X1_910 INVX1_636/Y BUFX4_94/Y gnd NAND3X1_321/C vdd NAND2X1
XINVX2_67 INVX2_67/A gnd INVX2_67/Y vdd INVX2
XINVX2_56 INVX2_56/A gnd INVX2_56/Y vdd INVX2
XNAND2X1_954 INVX2_85/A OR2X2_60/B gnd AOI22X1_131/B vdd NAND2X1
XNAND2X1_943 INVX1_327/A INVX1_674/Y gnd NAND2X1_943/Y vdd NAND2X1
XNAND2X1_932 INVX1_668/A INVX2_80/A gnd NAND2X1_932/Y vdd NAND2X1
XINVX2_78 INVX2_75/A gnd INVX2_78/Y vdd INVX2
XNAND2X1_998 INVX1_759/A NOR2X1_475/Y gnd BUFX2_34/A vdd NAND2X1
XNAND2X1_987 OAI21X1_912/C NAND2X1_987/B gnd NOR2X1_459/A vdd NAND2X1
XNAND2X1_976 MUX2X1_1/B INVX2_86/Y gnd AND2X2_91/B vdd NAND2X1
XNAND2X1_965 NAND2X1_963/Y AND2X2_88/Y gnd AOI21X1_239/A vdd NAND2X1
XINVX2_89 INVX2_89/A gnd INVX2_89/Y vdd INVX2
XFILL_4_7_1 gnd vdd FILL
XFILL_28_2_0 gnd vdd FILL
XFILL_29_7_1 gnd vdd FILL
XFILL_3_2_0 gnd vdd FILL
XOAI21X1_19 INVX1_19/Y BUFX4_19/Y OAI21X1_19/C gnd OAI21X1_19/Y vdd OAI21X1
XFILL_11_1_0 gnd vdd FILL
XFILL_12_6_1 gnd vdd FILL
XFILL_19_2_0 gnd vdd FILL
XDFFPOSX1_103 INVX1_216/A CLKBUF1_63/Y OAI21X1_147/C gnd vdd DFFPOSX1
XDFFPOSX1_125 DFFPOSX1_13/D CLKBUF1_51/Y INVX1_243/A gnd vdd DFFPOSX1
XDFFPOSX1_136 DFFPOSX1_24/D CLKBUF1_55/Y INVX2_14/A gnd vdd DFFPOSX1
XDFFPOSX1_114 NOR2X1_3/B CLKBUF1_62/Y NOR2X1_6/B gnd vdd DFFPOSX1
XDFFPOSX1_169 BUFX2_12/A CLKBUF1_10/Y XNOR2X1_25/Y gnd vdd DFFPOSX1
XDFFPOSX1_158 INVX2_87/A CLKBUF1_46/Y NOR2X1_69/Y gnd vdd DFFPOSX1
XDFFPOSX1_147 DFFPOSX1_35/D CLKBUF1_50/Y INVX1_285/A gnd vdd DFFPOSX1
XNAND2X1_217 INVX4_4/A AOI22X1_57/A gnd OAI21X1_295/C vdd NAND2X1
XNAND2X1_206 INVX4_4/Y INVX1_318/Y gnd OAI21X1_291/C vdd NAND2X1
XNAND2X1_228 INVX2_35/Y MUX2X1_2/Y gnd NAND2X1_228/Y vdd NAND2X1
XNAND2X1_239 INVX2_36/A INVX2_53/A gnd INVX1_329/A vdd NAND2X1
XBUFX4_190 BUFX4_188/A gnd BUFX4_190/Y vdd BUFX4
XNOR2X1_250 NOR2X1_250/A NOR2X1_247/Y gnd NOR2X1_250/Y vdd NOR2X1
XNOR2X1_261 INVX8_3/A MUX2X1_20/Y gnd INVX1_391/A vdd NOR2X1
XNOR2X1_294 OAI22X1_7/C OR2X2_34/A gnd NOR2X1_294/Y vdd NOR2X1
XNOR2X1_272 BUFX4_176/Y NOR2X1_203/B gnd AND2X2_45/A vdd NOR2X1
XNOR2X1_283 NOR3X1_56/A NOR3X1_56/C gnd NOR2X1_283/Y vdd NOR2X1
XOAI21X1_712 NOR2X1_308/B NOR2X1_143/A AOI21X1_186/Y gnd AOI21X1_203/B vdd OAI21X1
XOAI21X1_701 NAND2X1_595/B INVX8_4/A NAND2X1_572/Y gnd NOR2X1_339/B vdd OAI21X1
XOAI21X1_723 INVX2_18/A OAI21X1_722/Y OAI21X1_723/C gnd NAND3X1_165/A vdd OAI21X1
XOAI21X1_767 AND2X2_71/Y NOR2X1_371/Y AND2X2_56/B gnd OAI21X1_768/C vdd OAI21X1
XOAI21X1_745 INVX4_2/Y BUFX4_40/Y NAND2X1_334/Y gnd OAI21X1_745/Y vdd OAI21X1
XOAI21X1_734 INVX2_16/Y INVX2_17/Y OAI21X1_734/C gnd OAI21X1_734/Y vdd OAI21X1
XOAI21X1_756 NOR2X1_366/Y OAI21X1_755/Y AND2X2_69/Y gnd OAI21X1_756/Y vdd OAI21X1
XOAI21X1_778 AND2X2_74/Y AND2X2_72/Y BUFX4_127/Y gnd OAI21X1_779/C vdd OAI21X1
XOAI21X1_789 BUFX4_180/Y INVX1_442/Y OAI21X1_789/C gnd OAI21X1_789/Y vdd OAI21X1
XNAND2X1_762 NAND2X1_762/A NAND2X1_762/B gnd NAND2X1_18/B vdd NAND2X1
XNAND2X1_751 OAI21X1_79/Y BUFX4_135/Y gnd NAND2X1_753/A vdd NAND2X1
XNAND2X1_740 INVX1_523/Y BUFX4_202/Y gnd NAND3X1_211/C vdd NAND2X1
XNAND2X1_773 INVX1_545/Y BUFX4_204/Y gnd NAND3X1_233/C vdd NAND2X1
XNAND2X1_784 OAI21X1_90/Y BUFX4_132/Y gnd NAND2X1_784/Y vdd NAND2X1
XNAND2X1_795 NAND2X1_795/A NAND2X1_795/B gnd NAND2X1_29/B vdd NAND2X1
XFILL_43_0_0 gnd vdd FILL
XBUFX4_52 INVX8_3/Y gnd BUFX4_52/Y vdd BUFX4
XBUFX4_41 INVX8_8/Y gnd BUFX4_41/Y vdd BUFX4
XBUFX4_30 BUFX4_27/A gnd BUFX4_30/Y vdd BUFX4
XBUFX4_74 INVX8_1/Y gnd BUFX4_74/Y vdd BUFX4
XBUFX4_85 INVX8_9/Y gnd BUFX4_85/Y vdd BUFX4
XBUFX4_63 BUFX4_62/A gnd BUFX4_63/Y vdd BUFX4
XBUFX4_96 BUFX4_98/A gnd BUFX4_96/Y vdd BUFX4
XFILL_34_0_0 gnd vdd FILL
XFILL_35_5_1 gnd vdd FILL
XOR2X2_11 OR2X2_11/A OR2X2_11/B gnd OR2X2_11/Y vdd OR2X2
XOR2X2_33 OR2X2_33/A OR2X2_33/B gnd OR2X2_33/Y vdd OR2X2
XOR2X2_22 OR2X2_22/A OR2X2_22/B gnd OR2X2_23/B vdd OR2X2
XOR2X2_4 OR2X2_4/A OR2X2_4/B gnd OR2X2_4/Y vdd OR2X2
XOR2X2_44 OR2X2_44/A OR2X2_44/B gnd OR2X2_44/Y vdd OR2X2
XOR2X2_66 OR2X2_66/A OR2X2_66/B gnd OR2X2_67/B vdd OR2X2
XOR2X2_55 OR2X2_55/A OR2X2_55/B gnd OR2X2_55/Y vdd OR2X2
XXNOR2X1_6 XNOR2X1_6/A INVX2_6/A gnd XNOR2X1_7/B vdd XNOR2X1
XFILL_1_5_1 gnd vdd FILL
XFILL_25_0_0 gnd vdd FILL
XFILL_26_5_1 gnd vdd FILL
XFILL_0_0_0 gnd vdd FILL
XINVX8_11 INVX8_11/A gnd INVX8_11/Y vdd INVX8
XINVX1_6 gnd gnd INVX1_6/Y vdd INVX1
XOAI21X1_520 OAI21X1_520/A INVX8_3/A NAND2X1_477/Y gnd OR2X2_30/A vdd OAI21X1
XOAI21X1_531 INVX8_8/A MUX2X1_8/Y OAI21X1_351/C gnd OAI21X1_531/Y vdd OAI21X1
XOAI21X1_553 OAI22X1_9/A OAI22X1_25/C AOI22X1_71/A gnd OAI21X1_553/Y vdd OAI21X1
XOAI21X1_575 INVX1_396/Y MUX2X1_40/S NAND2X1_520/Y gnd OAI21X1_621/A vdd OAI21X1
XOAI21X1_542 INVX8_5/A MUX2X1_36/B NAND2X1_496/Y gnd NAND2X1_497/B vdd OAI21X1
XOAI21X1_564 INVX2_61/Y OAI22X1_8/A OAI21X1_564/C gnd OAI21X1_565/B vdd OAI21X1
XINVX1_617 INVX1_617/A gnd INVX1_617/Y vdd INVX1
XOAI21X1_597 INVX2_66/A INVX8_3/A AOI21X1_136/Y gnd AOI21X1_137/A vdd OAI21X1
XOAI21X1_586 MUX2X1_32/Y BUFX4_56/Y BUFX4_128/Y gnd AOI21X1_126/C vdd OAI21X1
XINVX1_606 INVX1_533/A gnd INVX1_606/Y vdd INVX1
XINVX1_628 INVX1_628/A gnd INVX1_628/Y vdd INVX1
XINVX1_639 INVX1_639/A gnd INVX1_639/Y vdd INVX1
XFILL_9_6_1 gnd vdd FILL
XFILL_8_1_0 gnd vdd FILL
XNAND2X1_570 AND2X2_52/Y NOR2X1_336/Y gnd NAND2X1_570/Y vdd NAND2X1
XNAND2X1_581 INVX4_7/A AND2X2_40/A gnd NAND2X1_581/Y vdd NAND2X1
XNAND2X1_592 INVX1_422/A NOR2X1_355/Y gnd NAND3X1_166/C vdd NAND2X1
XFILL_16_0_0 gnd vdd FILL
XFILL_17_5_1 gnd vdd FILL
XFILL_41_3_1 gnd vdd FILL
XOAI21X1_350 BUFX4_42/Y MUX2X1_7/Y OAI21X1_350/C gnd OAI21X1_350/Y vdd OAI21X1
XOAI21X1_361 NOR2X1_201/B NOR2X1_160/Y MUX2X1_47/S gnd OAI21X1_362/C vdd OAI21X1
XOAI21X1_383 INVX8_4/A OAI21X1_380/Y OAI21X1_383/C gnd NOR2X1_251/B vdd OAI21X1
XOAI21X1_372 INVX1_359/Y INVX4_4/A OAI21X1_372/C gnd OAI21X1_372/Y vdd OAI21X1
XAND2X2_6 AND2X2_6/A AND2X2_6/B gnd AND2X2_6/Y vdd AND2X2
XINVX1_403 INVX1_403/A gnd INVX1_403/Y vdd INVX1
XOAI21X1_394 INVX8_5/A OAI21X1_394/B NAND2X1_380/Y gnd OAI21X1_394/Y vdd OAI21X1
XINVX1_425 INVX1_425/A gnd INVX1_425/Y vdd INVX1
XINVX1_414 AND2X2_59/B gnd INVX1_414/Y vdd INVX1
XINVX1_469 BUFX2_40/A gnd INVX1_469/Y vdd INVX1
XINVX1_458 INVX1_458/A gnd INVX1_458/Y vdd INVX1
XINVX1_436 INVX1_436/A gnd INVX1_436/Y vdd INVX1
XINVX1_447 OR2X2_58/B gnd INVX1_447/Y vdd INVX1
XFILL_32_3_1 gnd vdd FILL
XFILL_23_3_1 gnd vdd FILL
XFILL_6_4_1 gnd vdd FILL
XMUX2X1_18 INVX1_239/A OR2X2_61/A INVX4_4/A gnd AND2X2_34/A vdd MUX2X1
XMUX2X1_29 MUX2X1_28/Y MUX2X1_29/B BUFX4_58/Y gnd MUX2X1_29/Y vdd MUX2X1
XFILL_14_3_1 gnd vdd FILL
XAOI22X1_1 INVX2_2/Y OR2X2_52/B INVX2_1/A INVX1_132/Y gnd AND2X2_3/B vdd AOI22X1
XOAI21X1_180 BUFX4_16/Y BUFX4_198/Y OAI21X1_847/Y gnd NAND3X1_45/C vdd OAI21X1
XOAI21X1_191 BUFX4_16/Y BUFX4_198/Y OAI21X1_866/Y gnd NAND3X1_67/C vdd OAI21X1
XINVX1_200 INVX1_200/A gnd INVX1_200/Y vdd INVX1
XINVX1_222 INVX1_222/A gnd INVX1_222/Y vdd INVX1
XINVX1_244 INVX1_244/A gnd INVX1_244/Y vdd INVX1
XINVX1_233 AOI21X1_7/A gnd INVX1_233/Y vdd INVX1
XINVX1_211 INVX1_211/A gnd INVX1_211/Y vdd INVX1
XINVX1_255 MUX2X1_9/B gnd INVX1_255/Y vdd INVX1
XINVX1_277 OR2X2_14/Y gnd INVX1_277/Y vdd INVX1
XINVX1_266 MUX2X1_1/A gnd INVX1_266/Y vdd INVX1
XINVX1_299 NOR2X1_64/Y gnd INVX1_299/Y vdd INVX1
XINVX1_288 INVX1_288/A gnd INVX1_288/Y vdd INVX1
XNAND2X1_22 BUFX4_24/Y NAND2X1_22/B gnd OAI21X1_22/C vdd NAND2X1
XNAND2X1_11 BUFX4_20/Y NAND2X1_11/B gnd OAI21X1_11/C vdd NAND2X1
XNAND2X1_33 NAND2X1_33/A BUFX4_28/Y gnd OAI21X1_33/C vdd NAND2X1
XNAND2X1_77 INVX2_9/A BUFX4_163/Y gnd NAND2X1_77/Y vdd NAND2X1
XNAND2X1_66 AND2X2_1/Y NOR2X1_1/Y gnd NOR2X1_2/B vdd NAND2X1
XNAND2X1_44 BUFX4_29/Y NAND2X1_44/B gnd OAI21X1_44/C vdd NAND2X1
XNAND2X1_55 BUFX4_25/Y NAND2X1_55/B gnd OAI21X1_55/C vdd NAND2X1
XNAND2X1_88 INVX1_273/A BUFX4_161/Y gnd NAND2X1_88/Y vdd NAND2X1
XNAND2X1_99 INVX1_99/Y NOR2X1_3/Y gnd BUFX4_194/A vdd NAND2X1
XFILL_35_2 gnd vdd FILL
XAOI21X1_215 INVX1_473/Y NOR2X1_382/Y BUFX2_49/A gnd AOI21X1_215/Y vdd AOI21X1
XAOI21X1_204 NOR2X1_367/Y INVX2_71/Y BUFX4_88/Y gnd AND2X2_69/B vdd AOI21X1
XAOI21X1_237 NOR2X1_438/Y AND2X2_95/A NOR2X1_437/Y gnd AOI21X1_237/Y vdd AOI21X1
XAOI21X1_248 AOI22X1_130/Y OAI21X1_910/Y AOI21X1_248/C gnd OAI21X1_932/A vdd AOI21X1
XAOI21X1_226 BUFX2_90/A INVX1_571/Y INVX1_572/Y gnd AOI21X1_226/Y vdd AOI21X1
XAOI21X1_259 AOI21X1_259/A AOI21X1_259/B INVX4_12/A gnd OAI21X1_993/B vdd AOI21X1
XAOI22X1_42 MUX2X1_14/A AND2X2_12/A AND2X2_11/A OR2X2_64/A gnd OR2X2_9/A vdd AOI22X1
XAOI22X1_31 AOI22X1_31/A BUFX4_238/Y BUFX4_259/Y AOI22X1_31/D gnd AOI22X1_31/Y vdd
+ AOI22X1
XAOI22X1_20 AOI22X1_20/A BUFX4_238/Y BUFX4_256/Y AOI22X1_20/D gnd AOI22X1_20/Y vdd
+ AOI22X1
XAOI22X1_53 AOI22X1_53/A BUFX4_231/Y BUFX4_150/Y INVX1_327/A gnd NOR2X1_41/B vdd AOI22X1
XAOI22X1_75 INVX1_349/Y AOI22X1_75/B INVX1_305/Y AOI22X1_75/D gnd AOI22X1_75/Y vdd
+ AOI22X1
XAOI22X1_64 AOI22X1_64/A BUFX4_233/Y BUFX4_148/Y OR2X2_54/A gnd NOR2X1_56/B vdd AOI22X1
XAOI22X1_97 OAI22X1_8/B BUFX4_153/Y OR2X2_24/Y AOI22X1_97/D gnd AOI22X1_97/Y vdd AOI22X1
XAOI22X1_86 AOI22X1_86/A BUFX4_154/Y OR2X2_24/Y AND2X2_35/B gnd AOI22X1_86/Y vdd AOI22X1
XNAND3X1_208 INVX1_522/Y BUFX4_206/Y BUFX4_33/Y gnd NAND3X1_208/Y vdd NAND3X1
XNAND3X1_219 BUFX4_218/Y NAND3X1_218/Y NAND3X1_219/C gnd NAND2X1_753/B vdd NAND3X1
XOAI22X1_4 INVX2_1/Y INVX1_495/A INVX2_3/A AOI22X1_6/D gnd NOR3X1_17/A vdd OAI22X1
XDFFPOSX1_329 INVX1_283/A CLKBUF1_1/Y OAI21X1_897/Y gnd vdd DFFPOSX1
XDFFPOSX1_318 INVX2_13/A CLKBUF1_42/Y OAI21X1_886/Y gnd vdd DFFPOSX1
XDFFPOSX1_307 INVX1_234/A CLKBUF1_34/Y OAI21X1_880/Y gnd vdd DFFPOSX1
XFILL_37_2_1 gnd vdd FILL
XNOR2X1_410 NOR2X1_410/A NOR2X1_410/B gnd NOR2X1_410/Y vdd NOR2X1
XNOR2X1_432 NOR2X1_432/A INVX1_691/A gnd NOR2X1_432/Y vdd NOR2X1
XNOR2X1_421 INVX1_664/A INVX1_665/Y gnd NOR2X1_422/B vdd NOR2X1
XNOR2X1_443 OR2X2_54/A OR2X2_54/B gnd OAI22X1_51/B vdd NOR2X1
XNOR2X1_465 OR2X2_68/Y NOR2X1_465/B gnd NOR2X1_465/Y vdd NOR2X1
XNOR2X1_454 NOR2X1_454/A NOR2X1_454/B gnd NOR2X1_454/Y vdd NOR2X1
XNOR2X1_476 INVX4_12/Y INVX2_87/Y gnd NOR2X1_476/Y vdd NOR2X1
XNOR2X1_487 NOR2X1_487/A NOR3X1_78/C gnd NOR2X1_487/Y vdd NOR2X1
XOAI21X1_905 INVX1_325/A INVX2_83/Y NAND2X1_943/Y gnd NOR3X1_70/A vdd OAI21X1
XOAI21X1_916 NOR2X1_445/Y NAND2X1_943/Y OAI21X1_906/C gnd AOI21X1_251/B vdd OAI21X1
XOAI21X1_927 OR2X2_65/Y AND2X2_94/Y INVX1_708/Y gnd OAI21X1_927/Y vdd OAI21X1
XFILL_20_1_1 gnd vdd FILL
XOAI21X1_938 OAI21X1_938/A NAND2X1_992/Y NOR2X1_455/Y gnd OAI21X1_938/Y vdd OAI21X1
XOAI21X1_949 NOR3X1_77/Y NOR3X1_78/Y INVX4_12/Y gnd AOI21X1_263/A vdd OAI21X1
XINVX2_35 INVX2_35/A gnd INVX2_35/Y vdd INVX2
XINVX2_13 INVX2_13/A gnd INVX2_13/Y vdd INVX2
XINVX2_24 INVX2_24/A gnd INVX2_24/Y vdd INVX2
XNAND2X1_911 NAND2X1_909/Y NAND2X1_911/B gnd NAND2X1_63/B vdd NAND2X1
XNAND2X1_900 OAI21X1_92/Y BUFX4_59/Y gnd NAND2X1_900/Y vdd NAND2X1
XNAND2X1_922 OR2X2_8/B NOR2X1_411/Y gnd OAI21X1_878/C vdd NAND2X1
XINVX2_57 INVX2_57/A gnd INVX2_57/Y vdd INVX2
XINVX2_68 INVX2_68/A gnd INVX2_68/Y vdd INVX2
XINVX2_46 INVX2_46/A gnd INVX2_46/Y vdd INVX2
XNAND2X1_955 OR2X2_61/A OR2X2_61/B gnd AOI22X1_131/C vdd NAND2X1
XNAND2X1_944 INVX1_325/A INVX2_83/Y gnd OAI21X1_906/C vdd NAND2X1
XNAND2X1_933 INVX1_668/Y INVX2_80/Y gnd NAND2X1_933/Y vdd NAND2X1
XINVX2_79 INVX2_79/A gnd INVX2_79/Y vdd INVX2
XAND2X2_100 AND2X2_100/A NAND3X1_1/B gnd AND2X2_100/Y vdd AND2X2
XNAND2X1_977 AND2X2_91/Y NAND2X1_975/Y gnd NAND2X1_977/Y vdd NAND2X1
XNAND2X1_988 AND2X2_86/A AND2X2_86/B gnd NOR2X1_459/B vdd NAND2X1
XNAND2X1_966 AND2X2_86/Y NOR2X1_430/Y gnd OAI21X1_913/A vdd NAND2X1
XNAND2X1_999 INVX2_89/Y AND2X2_98/Y gnd NOR2X1_487/A vdd NAND2X1
XFILL_3_2_1 gnd vdd FILL
XFILL_28_2_1 gnd vdd FILL
XFILL_11_1_1 gnd vdd FILL
XFILL_19_2_1 gnd vdd FILL
XDFFPOSX1_126 DFFPOSX1_14/D CLKBUF1_32/Y INVX1_245/A gnd vdd DFFPOSX1
XDFFPOSX1_137 DFFPOSX1_25/D CLKBUF1_19/Y INVX1_261/A gnd vdd DFFPOSX1
XDFFPOSX1_104 INVX1_217/A CLKBUF1_3/Y OAI21X1_149/C gnd vdd DFFPOSX1
XDFFPOSX1_115 NOR2X1_3/A CLKBUF1_62/Y NOR2X1_6/A gnd vdd DFFPOSX1
XDFFPOSX1_159 INVX4_12/A CLKBUF1_4/Y XNOR2X1_5/Y gnd vdd DFFPOSX1
XDFFPOSX1_148 DFFPOSX1_36/D CLKBUF1_19/Y INVX1_288/A gnd vdd DFFPOSX1
XNAND2X1_207 NOR2X1_99/A NOR2X1_332/B gnd AND2X2_59/A vdd NAND2X1
XNAND2X1_229 NAND2X1_228/Y INVX1_402/A gnd INVX1_403/A vdd NAND2X1
XNAND2X1_218 INVX2_32/A MUX2X1_44/A gnd INVX1_408/A vdd NAND2X1
XBUFX4_180 BUFX4_178/A gnd BUFX4_180/Y vdd BUFX4
XBUFX4_191 BUFX4_194/A gnd OR2X2_2/B vdd BUFX4
XNOR2X1_240 NOR2X1_239/Y NOR2X1_238/Y gnd INVX1_387/A vdd NOR2X1
XNOR2X1_251 INVX8_3/A NOR2X1_251/B gnd AND2X2_40/A vdd NOR2X1
XNOR2X1_273 INVX4_5/Y AND2X2_45/Y gnd NOR2X1_273/Y vdd NOR2X1
XNOR2X1_284 NOR2X1_284/A NOR2X1_284/B gnd NOR2X1_284/Y vdd NOR2X1
XNOR2X1_262 NOR2X1_262/A NOR2X1_135/B gnd AOI22X1_94/D vdd NOR2X1
XNOR2X1_295 NOR2X1_295/A NOR2X1_295/B gnd OR2X2_35/B vdd NOR2X1
XOAI21X1_702 INVX2_55/Y NOR2X1_339/B BUFX4_128/Y gnd OAI21X1_702/Y vdd OAI21X1
XOAI21X1_724 INVX4_3/Y BUFX4_38/Y NAND2X1_583/Y gnd INVX1_421/A vdd OAI21X1
XOAI21X1_713 NOR2X1_80/Y INVX2_19/Y AOI21X1_203/B gnd OAI21X1_732/A vdd OAI21X1
XOAI21X1_757 OAI21X1_736/Y AND2X2_70/B MUX2X1_49/S gnd OAI22X1_42/B vdd OAI21X1
XOAI21X1_746 INVX8_5/A OAI21X1_745/Y NAND2X1_594/Y gnd OAI21X1_747/B vdd OAI21X1
XOAI21X1_735 INVX1_422/A OAI21X1_734/Y OAI21X1_735/C gnd NAND3X1_167/A vdd OAI21X1
XOAI21X1_779 OAI21X1_779/A BUFX4_127/Y OAI21X1_779/C gnd OAI21X1_779/Y vdd OAI21X1
XOAI21X1_768 AND2X2_56/B OAI22X1_34/B OAI21X1_768/C gnd AOI21X1_210/B vdd OAI21X1
XNAND2X1_730 OAI21X1_72/Y BUFX4_132/Y gnd NAND2X1_730/Y vdd NAND2X1
XNAND2X1_741 NAND2X1_739/Y NAND2X1_741/B gnd NAND2X1_11/B vdd NAND2X1
XNAND2X1_763 OAI21X1_83/Y BUFX4_133/Y gnd NAND2X1_765/A vdd NAND2X1
XNAND2X1_752 INVX1_531/Y BUFX4_203/Y gnd NAND3X1_219/C vdd NAND2X1
XNAND2X1_774 NAND2X1_774/A NAND2X1_774/B gnd NAND2X1_22/B vdd NAND2X1
XNAND2X1_796 OAI21X1_94/Y BUFX4_131/Y gnd NAND2X1_798/A vdd NAND2X1
XNAND2X1_785 INVX1_553/Y BUFX4_205/Y gnd NAND3X1_241/C vdd NAND2X1
XFILL_43_0_1 gnd vdd FILL
XBUFX4_20 BUFX4_22/A gnd BUFX4_20/Y vdd BUFX4
XBUFX4_42 INVX8_8/Y gnd BUFX4_42/Y vdd BUFX4
XBUFX4_53 INVX8_3/Y gnd BUFX4_53/Y vdd BUFX4
XBUFX4_31 BUFX4_27/A gnd BUFX4_31/Y vdd BUFX4
XBUFX4_86 BUFX4_88/A gnd BUFX4_86/Y vdd BUFX4
XBUFX4_75 INVX8_1/Y gnd BUFX4_75/Y vdd BUFX4
XBUFX4_64 BUFX4_65/A gnd BUFX4_64/Y vdd BUFX4
XBUFX4_97 BUFX4_98/A gnd BUFX4_97/Y vdd BUFX4
XFILL_34_0_1 gnd vdd FILL
XFILL_10_1 gnd vdd FILL
XOR2X2_12 OR2X2_12/A OR2X2_12/B gnd OR2X2_12/Y vdd OR2X2
XOR2X2_23 OR2X2_23/A OR2X2_23/B gnd OR2X2_23/Y vdd OR2X2
XOR2X2_45 OR2X2_45/A OR2X2_45/B gnd OR2X2_45/Y vdd OR2X2
XOR2X2_34 OR2X2_34/A OR2X2_34/B gnd OR2X2_34/Y vdd OR2X2
XOR2X2_56 OR2X2_56/A OR2X2_56/B gnd OR2X2_56/Y vdd OR2X2
XOR2X2_67 OR2X2_67/A OR2X2_67/B gnd OR2X2_67/Y vdd OR2X2
XOR2X2_5 OR2X2_5/A OR2X2_5/B gnd OR2X2_5/Y vdd OR2X2
XXNOR2X1_7 AOI21X1_6/Y XNOR2X1_7/B gnd XNOR2X1_7/Y vdd XNOR2X1
XFILL_25_0_1 gnd vdd FILL
XFILL_0_0_1 gnd vdd FILL
XINVX8_12 INVX8_12/A gnd INVX8_12/Y vdd INVX8
XINVX1_7 gnd gnd INVX1_7/Y vdd INVX1
XOAI21X1_510 NOR2X1_149/Y OAI21X1_463/A OAI22X1_15/B gnd AOI21X1_96/B vdd OAI21X1
XOAI21X1_532 MUX2X1_40/S AOI21X1_93/Y NAND2X1_490/Y gnd OAI21X1_576/B vdd OAI21X1
XOAI21X1_521 OAI22X1_30/A OR2X2_30/Y OAI21X1_521/C gnd NOR2X1_250/A vdd OAI21X1
XOAI21X1_543 BUFX4_216/Y OAI21X1_543/B NAND2X1_497/Y gnd MUX2X1_34/A vdd OAI21X1
XOAI21X1_554 NOR2X1_253/B NOR2X1_296/A AOI21X1_114/Y gnd INVX2_61/A vdd OAI21X1
XOAI21X1_565 NOR2X1_281/A OAI21X1_565/B AOI21X1_117/Y gnd OAI21X1_565/Y vdd OAI21X1
XOAI21X1_587 OAI22X1_30/A OAI21X1_779/A AOI21X1_127/Y gnd OR2X2_35/A vdd OAI21X1
XOAI21X1_576 BUFX4_216/Y OAI21X1_576/B NAND2X1_521/Y gnd NOR2X1_329/B vdd OAI21X1
XOAI21X1_598 NOR2X1_103/Y INVX8_12/Y AOI22X1_100/Y gnd OAI21X1_598/Y vdd OAI21X1
XINVX1_607 INVX1_607/A gnd INVX1_607/Y vdd INVX1
XINVX1_618 INVX1_545/A gnd INVX1_618/Y vdd INVX1
XINVX1_629 INVX1_556/A gnd INVX1_629/Y vdd INVX1
XDFFPOSX1_490 BUFX2_57/A CLKBUF1_45/Y NAND3X1_43/Y gnd vdd DFFPOSX1
XFILL_8_1_1 gnd vdd FILL
XNAND2X1_571 INVX1_413/A INVX1_328/A gnd AND2X2_62/A vdd NAND2X1
XNAND2X1_560 BUFX4_53/Y NOR2X1_328/Y gnd AOI21X1_163/B vdd NAND2X1
XNAND2X1_593 INVX2_18/A INVX1_422/A gnd NOR2X1_356/B vdd NAND2X1
XNAND2X1_582 NOR2X1_81/Y AND2X2_64/B gnd NOR2X1_356/A vdd NAND2X1
XFILL_16_0_1 gnd vdd FILL
XFILL_10_7_0 gnd vdd FILL
XOAI21X1_340 INVX1_352/Y NOR2X1_185/B AND2X2_21/A gnd OAI21X1_341/C vdd OAI21X1
XOAI21X1_351 INVX8_8/A MUX2X1_10/Y OAI21X1_351/C gnd OR2X2_19/A vdd OAI21X1
XOAI21X1_362 OAI21X1_410/A MUX2X1_47/S OAI21X1_362/C gnd MUX2X1_26/B vdd OAI21X1
XOAI21X1_373 INVX8_8/A OAI21X1_372/Y BUFX4_187/Y gnd AND2X2_27/B vdd OAI21X1
XAND2X2_7 AND2X2_5/Y AND2X2_7/B gnd AND2X2_8/B vdd AND2X2
XINVX1_415 OR2X2_39/B gnd INVX1_415/Y vdd INVX1
XINVX1_404 INVX1_404/A gnd INVX1_404/Y vdd INVX1
XOAI21X1_384 NOR2X1_160/B BUFX4_39/Y OAI21X1_631/C gnd INVX1_362/A vdd OAI21X1
XOAI21X1_395 BUFX4_41/Y MUX2X1_10/Y NAND2X1_381/Y gnd NAND2X1_416/B vdd OAI21X1
XINVX1_426 OR2X2_15/B gnd INVX1_426/Y vdd INVX1
XINVX1_459 INVX1_459/A gnd INVX1_459/Y vdd INVX1
XINVX1_437 BUFX4_268/Y gnd INVX1_437/Y vdd INVX1
XINVX1_448 OR2X2_57/B gnd INVX1_448/Y vdd INVX1
XNAND2X1_390 INVX8_3/A NAND2X1_482/B gnd OAI21X1_406/C vdd NAND2X1
XMUX2X1_19 MUX2X1_19/A MUX2X1_19/B INVX8_5/A gnd MUX2X1_19/Y vdd MUX2X1
XFILL_42_6_0 gnd vdd FILL
XAOI22X1_2 INVX2_3/Y BUFX2_91/A INVX2_2/A AOI22X1_2/D gnd NAND3X1_2/A vdd AOI22X1
XOAI21X1_170 BUFX4_15/Y BUFX4_200/Y OAI21X1_827/Y gnd NAND3X1_25/C vdd OAI21X1
XOAI21X1_181 BUFX4_12/Y BUFX4_199/Y OAI21X1_849/Y gnd NAND3X1_47/C vdd OAI21X1
XOAI21X1_192 BUFX4_16/Y BUFX4_198/Y OAI21X1_868/Y gnd NAND3X1_69/C vdd OAI21X1
XINVX1_201 INVX1_201/A gnd INVX1_201/Y vdd INVX1
XINVX1_223 NOR2X1_8/B gnd INVX1_223/Y vdd INVX1
XINVX1_234 INVX1_234/A gnd INVX1_234/Y vdd INVX1
XINVX1_212 INVX1_212/A gnd INVX1_212/Y vdd INVX1
XINVX1_256 MUX2X1_6/B gnd INVX1_256/Y vdd INVX1
XINVX1_245 INVX1_245/A gnd INVX1_245/Y vdd INVX1
XINVX1_267 BUFX4_232/Y gnd INVX1_267/Y vdd INVX1
XINVX1_289 NOR2X1_58/Y gnd INVX1_289/Y vdd INVX1
XINVX1_278 INVX1_278/A gnd INVX1_278/Y vdd INVX1
XNAND2X1_23 BUFX4_18/Y NAND2X1_23/B gnd OAI21X1_23/C vdd NAND2X1
XNAND2X1_12 BUFX4_22/Y NAND2X1_12/B gnd OAI21X1_12/C vdd NAND2X1
XNAND2X1_34 BUFX4_28/Y NAND2X1_34/B gnd OAI21X1_34/C vdd NAND2X1
XNAND2X1_67 INVX1_230/A BUFX4_162/Y gnd NAND2X1_67/Y vdd NAND2X1
XNAND2X1_45 BUFX4_26/Y NAND2X1_45/B gnd OAI21X1_45/C vdd NAND2X1
XNAND2X1_56 BUFX4_31/Y NAND2X1_56/B gnd NAND2X1_56/Y vdd NAND2X1
XNAND2X1_89 INVX1_274/A BUFX4_157/Y gnd NAND2X1_89/Y vdd NAND2X1
XNAND2X1_78 INVX2_10/A BUFX4_159/Y gnd NAND2X1_78/Y vdd NAND2X1
XFILL_35_3 gnd vdd FILL
XFILL_33_6_0 gnd vdd FILL
XAOI21X1_216 BUFX2_53/A XNOR2X1_51/A BUFX2_54/A gnd AOI21X1_216/Y vdd AOI21X1
XAOI21X1_205 INVX8_8/A INVX2_21/A OR2X2_25/A gnd AND2X2_70/A vdd AOI21X1
XAOI21X1_238 AOI21X1_238/A NOR2X1_440/Y NOR2X1_441/Y gnd INVX1_710/A vdd AOI21X1
XAOI21X1_249 NOR2X1_459/Y INVX1_710/Y INVX1_695/A gnd AOI21X1_249/Y vdd AOI21X1
XAOI21X1_227 INVX2_78/Y BUFX2_87/A OAI22X1_47/Y gnd AOI21X1_227/Y vdd AOI21X1
XAOI22X1_10 AOI22X1_10/A BUFX4_238/Y BUFX4_256/Y AOI22X1_10/D gnd AOI22X1_10/Y vdd
+ AOI22X1
XAOI22X1_21 AOI22X1_21/A BUFX4_238/Y BUFX4_256/Y AOI22X1_21/D gnd AOI22X1_21/Y vdd
+ AOI22X1
XAOI22X1_32 AOI22X1_32/A BUFX4_238/Y BUFX4_256/Y AOI22X1_32/D gnd AOI22X1_32/Y vdd
+ AOI22X1
XAOI22X1_54 AOI22X1_54/A BUFX4_235/Y BUFX4_150/Y INVX1_325/A gnd INVX1_260/A vdd AOI22X1
XAOI22X1_43 INVX1_351/A BUFX4_231/Y BUFX4_150/Y OR2X2_63/A gnd XNOR2X1_6/A vdd AOI22X1
XAOI22X1_65 AOI22X1_65/A BUFX4_233/Y BUFX4_148/Y OR2X2_53/A gnd NOR2X1_58/B vdd AOI22X1
XAOI22X1_98 AOI22X1_98/A INVX4_9/A AOI22X1_98/C BUFX4_53/Y gnd OAI22X1_34/B vdd AOI22X1
XAOI22X1_87 AOI22X1_87/A AOI22X1_87/B NOR2X1_237/Y NOR2X1_194/Y gnd AOI22X1_87/Y vdd
+ AOI22X1
XAOI22X1_76 BUFX4_90/Y NOR2X1_196/Y NOR2X1_194/Y INVX1_370/Y gnd AOI22X1_76/Y vdd
+ AOI22X1
XFILL_24_6_0 gnd vdd FILL
XNAND3X1_209 BUFX4_220/Y NAND3X1_208/Y NAND3X1_209/C gnd NAND2X1_738/B vdd NAND3X1
XOAI22X1_5 INVX2_3/Y OR2X2_49/B INVX2_2/A AOI22X1_4/D gnd NOR3X1_17/B vdd OAI22X1
XFILL_7_7_0 gnd vdd FILL
XFILL_15_6_0 gnd vdd FILL
XDFFPOSX1_308 INVX1_243/A CLKBUF1_25/Y NOR2X1_413/Y gnd vdd DFFPOSX1
XDFFPOSX1_319 INVX2_14/A CLKBUF1_40/Y OAI21X1_887/Y gnd vdd DFFPOSX1
XNOR2X1_400 NOR2X1_400/A NOR2X1_400/B gnd AND2X2_79/A vdd NOR2X1
XNOR2X1_433 OR2X2_62/B INVX1_686/Y gnd INVX1_708/A vdd NOR2X1
XNOR2X1_422 NOR2X1_422/A NOR2X1_422/B gnd NOR2X1_422/Y vdd NOR2X1
XNOR2X1_411 OAI22X1_6/Y INVX2_79/Y gnd NOR2X1_411/Y vdd NOR2X1
XNOR2X1_455 INVX2_51/A INVX2_49/A gnd NOR2X1_455/Y vdd NOR2X1
XNOR2X1_444 OR2X2_55/A OR2X2_55/B gnd OAI22X1_51/D vdd NOR2X1
XNOR2X1_477 INVX4_12/A INVX2_87/Y gnd NOR2X1_477/Y vdd NOR2X1
XNOR2X1_466 OR2X2_69/A OR2X2_69/B gnd NOR2X1_466/Y vdd NOR2X1
XNOR2X1_488 OAI22X1_58/B NOR2X1_488/B gnd OR2X2_70/B vdd NOR2X1
XOAI21X1_906 INVX1_327/A INVX1_674/Y OAI21X1_906/C gnd NOR3X1_70/C vdd OAI21X1
XOAI21X1_928 INVX2_85/Y OR2X2_60/B NAND2X1_984/Y gnd OAI21X1_928/Y vdd OAI21X1
XOAI21X1_917 MUX2X1_1/B INVX2_86/Y NOR2X1_446/Y gnd AND2X2_91/A vdd OAI21X1
XOAI21X1_939 MUX2X1_9/B INVX2_84/Y AND2X2_87/A gnd NOR3X1_72/A vdd OAI21X1
XINVX2_36 INVX2_36/A gnd INVX2_36/Y vdd INVX2
XINVX2_25 INVX2_25/A gnd INVX2_25/Y vdd INVX2
XINVX2_14 INVX2_14/A gnd INVX2_14/Y vdd INVX2
XNAND2X1_912 OAI21X1_96/Y BUFX4_59/Y gnd NAND2X1_912/Y vdd NAND2X1
XNAND2X1_901 INVX1_630/Y BUFX4_94/Y gnd NAND3X1_315/C vdd NAND2X1
XINVX2_58 INVX2_58/A gnd INVX2_58/Y vdd INVX2
XINVX2_47 INVX2_47/A gnd INVX2_47/Y vdd INVX2
XINVX2_69 INVX2_69/A gnd INVX2_69/Y vdd INVX2
XNAND2X1_945 MUX2X1_4/B INVX1_677/Y gnd AND2X2_86/A vdd NAND2X1
XNAND2X1_934 OR2X2_54/A OR2X2_54/B gnd NAND2X1_934/Y vdd NAND2X1
XNAND2X1_923 OR2X2_8/A NOR2X1_411/Y gnd OAI21X1_879/C vdd NAND2X1
XAND2X2_101 OAI22X1_58/C AND2X2_101/B gnd AND2X2_101/Y vdd AND2X2
XNAND2X1_978 INVX1_457/A INVX1_672/Y gnd AOI21X1_241/A vdd NAND2X1
XNAND2X1_956 OR2X2_62/A OR2X2_62/B gnd NAND2X1_956/Y vdd NAND2X1
XNAND2X1_989 AND2X2_83/B AND2X2_83/A gnd NAND2X1_989/Y vdd NAND2X1
XNAND2X1_967 INVX1_449/A INVX1_679/Y gnd AOI21X1_238/A vdd NAND2X1
XFILL_30_4_0 gnd vdd FILL
XDFFPOSX1_127 DFFPOSX1_15/D CLKBUF1_12/Y INVX1_249/A gnd vdd DFFPOSX1
XDFFPOSX1_105 INVX1_218/A CLKBUF1_30/Y OAI21X1_151/C gnd vdd DFFPOSX1
XDFFPOSX1_116 INVX2_89/A CLKBUF1_62/Y OR2X2_1/B gnd vdd DFFPOSX1
XDFFPOSX1_138 DFFPOSX1_26/D CLKBUF1_42/Y INVX1_264/A gnd vdd DFFPOSX1
XDFFPOSX1_149 DFFPOSX1_37/D CLKBUF1_51/Y NOR2X1_62/A gnd vdd DFFPOSX1
XNAND2X1_208 INVX4_4/A AOI22X1_60/A gnd NAND2X1_208/Y vdd NAND2X1
XNAND2X1_219 INVX4_4/Y INVX1_322/Y gnd OAI21X1_296/C vdd NAND2X1
XFILL_38_5_0 gnd vdd FILL
XBUFX4_181 BUFX4_178/A gnd BUFX4_181/Y vdd BUFX4
XBUFX4_170 BUFX4_171/A gnd BUFX4_170/Y vdd BUFX4
XNOR2X1_241 INVX8_7/A NOR2X1_241/B gnd NOR2X1_241/Y vdd NOR2X1
XNOR2X1_230 NOR2X1_230/A NOR2X1_230/B gnd NOR2X1_230/Y vdd NOR2X1
XNOR2X1_252 INVX2_44/A MUX2X1_9/Y gnd OAI22X1_24/B vdd NOR2X1
XBUFX4_192 BUFX4_194/A gnd BUFX4_192/Y vdd BUFX4
XNOR2X1_274 INVX2_42/Y MUX2X1_35/A gnd OAI22X1_37/A vdd NOR2X1
XNOR2X1_285 INVX2_41/A MUX2X1_6/Y gnd NOR2X1_285/Y vdd NOR2X1
XNOR2X1_263 NOR2X1_255/Y NOR2X1_263/B gnd NOR2X1_263/Y vdd NOR2X1
XNOR2X1_296 NOR2X1_296/A NOR2X1_296/B gnd NOR2X1_296/Y vdd NOR2X1
XOAI21X1_703 NOR2X1_338/Y OAI21X1_702/Y INVX2_65/A gnd OAI21X1_703/Y vdd OAI21X1
XOAI21X1_714 AND2X2_64/B AND2X2_65/B BUFX4_93/Y gnd AOI21X1_187/C vdd OAI21X1
XFILL_21_4_0 gnd vdd FILL
XOAI21X1_758 BUFX4_53/Y NOR2X1_328/B NAND2X1_598/Y gnd OAI21X1_758/Y vdd OAI21X1
XOAI21X1_747 INVX8_4/A OAI21X1_747/B NAND2X1_595/Y gnd MUX2X1_54/A vdd OAI21X1
XOAI21X1_725 BUFX4_225/Y OAI21X1_725/B OAI21X1_725/C gnd OAI22X1_44/C vdd OAI21X1
XOAI21X1_736 INVX4_2/Y INVX8_8/A NAND2X1_365/Y gnd OAI21X1_736/Y vdd OAI21X1
XOAI21X1_769 BUFX4_55/Y MUX2X1_45/Y OAI21X1_769/C gnd OAI21X1_770/B vdd OAI21X1
XOAI21X1_1060 OAI21X1_993/B NOR3X1_73/B INVX1_757/A gnd NOR2X1_488/B vdd OAI21X1
XNAND2X1_720 NAND2X1_718/Y NAND2X1_720/B gnd NAND2X1_4/B vdd NAND2X1
XNAND2X1_753 NAND2X1_753/A NAND2X1_753/B gnd NAND2X1_15/B vdd NAND2X1
XNAND2X1_742 OAI21X1_76/Y BUFX4_131/Y gnd NAND2X1_742/Y vdd NAND2X1
XNAND2X1_731 INVX1_517/Y BUFX4_202/Y gnd NAND3X1_205/C vdd NAND2X1
XNAND2X1_764 INVX1_539/Y BUFX4_204/Y gnd NAND3X1_227/C vdd NAND2X1
XNAND2X1_797 INVX1_561/Y BUFX4_204/Y gnd NAND3X1_249/C vdd NAND2X1
XNAND2X1_786 NAND2X1_784/Y NAND2X1_786/B gnd NAND2X1_26/B vdd NAND2X1
XNAND2X1_775 OAI21X1_87/Y BUFX4_133/Y gnd NAND2X1_777/A vdd NAND2X1
XFILL_4_5_0 gnd vdd FILL
XFILL_29_5_0 gnd vdd FILL
XFILL_12_4_0 gnd vdd FILL
XINVX8_1 reset gnd INVX8_1/Y vdd INVX8
XBUFX4_10 BUFX4_9/A gnd BUFX4_10/Y vdd BUFX4
XBUFX4_43 INVX8_8/Y gnd BUFX4_43/Y vdd BUFX4
XBUFX4_21 BUFX4_22/A gnd BUFX4_21/Y vdd BUFX4
XBUFX4_32 BUFX4_27/A gnd BUFX4_32/Y vdd BUFX4
XBUFX4_54 INVX8_3/Y gnd BUFX4_54/Y vdd BUFX4
XBUFX4_87 BUFX4_88/A gnd BUFX4_87/Y vdd BUFX4
XBUFX4_76 INVX8_1/Y gnd BUFX4_76/Y vdd BUFX4
XBUFX4_65 BUFX4_65/A gnd BUFX4_65/Y vdd BUFX4
XBUFX4_98 BUFX4_98/A gnd BUFX4_98/Y vdd BUFX4
XFILL_10_2 gnd vdd FILL
XOR2X2_13 OR2X2_13/A OR2X2_13/B gnd OR2X2_13/Y vdd OR2X2
XOR2X2_24 OR2X2_24/A OR2X2_24/B gnd OR2X2_24/Y vdd OR2X2
XOR2X2_35 OR2X2_35/A OR2X2_35/B gnd OR2X2_35/Y vdd OR2X2
XOR2X2_46 OR2X2_46/A OR2X2_46/B gnd OR2X2_46/Y vdd OR2X2
XOR2X2_57 OR2X2_57/A OR2X2_57/B gnd OR2X2_57/Y vdd OR2X2
XOR2X2_6 OR2X2_6/A OR2X2_6/B gnd OR2X2_6/Y vdd OR2X2
XOR2X2_68 OR2X2_68/A OR2X2_68/B gnd OR2X2_68/Y vdd OR2X2
XXNOR2X1_8 XNOR2X1_6/A INVX2_6/Y gnd XNOR2X1_8/Y vdd XNOR2X1
XINVX8_13 INVX8_13/A gnd INVX8_13/Y vdd INVX8
XOAI21X1_522 INVX1_365/Y BUFX4_52/Y NAND2X1_482/Y gnd OAI21X1_523/A vdd OAI21X1
XOAI21X1_500 OAI22X1_11/A INVX8_12/Y AOI22X1_86/Y gnd AOI21X1_89/C vdd OAI21X1
XOAI21X1_511 OAI22X1_11/A AOI22X1_74/C AOI22X1_74/A gnd AOI21X1_96/C vdd OAI21X1
XINVX1_8 gnd gnd INVX1_8/Y vdd INVX1
XOAI21X1_544 OR2X2_30/B OAI22X1_30/A INVX4_6/A gnd AOI21X1_110/B vdd OAI21X1
XOAI21X1_566 OAI21X1_472/Y BUFX4_52/Y BUFX4_128/Y gnd AOI21X1_118/C vdd OAI21X1
XOAI21X1_533 OAI21X1_576/B INVX8_4/A NAND2X1_489/Y gnd NOR2X1_315/A vdd OAI21X1
XOAI21X1_555 AOI22X1_97/D INVX2_61/A NOR2X1_276/Y gnd OAI21X1_555/Y vdd OAI21X1
XOAI21X1_599 INVX2_65/Y OAI21X1_599/B AOI21X1_140/Y gnd NOR2X1_300/B vdd OAI21X1
XOAI21X1_588 OAI22X1_8/D OAI21X1_564/C OAI21X1_588/C gnd OAI21X1_588/Y vdd OAI21X1
XOAI21X1_577 INVX8_3/A NOR2X1_329/B OAI21X1_577/C gnd NOR2X1_373/B vdd OAI21X1
XINVX1_608 INVX1_535/A gnd INVX1_608/Y vdd INVX1
XINVX1_619 INVX1_619/A gnd INVX1_619/Y vdd INVX1
XDFFPOSX1_480 BUFX2_47/A CLKBUF1_7/Y NAND3X1_23/Y gnd vdd DFFPOSX1
XDFFPOSX1_491 BUFX2_58/A CLKBUF1_45/Y NAND3X1_45/Y gnd vdd DFFPOSX1
XNAND2X1_550 INVX8_5/A MUX2X1_42/Y gnd NAND2X1_550/Y vdd NAND2X1
XNAND2X1_572 INVX8_4/A NAND2X1_572/B gnd NAND2X1_572/Y vdd NAND2X1
XNAND2X1_561 INVX4_9/A NAND2X1_561/B gnd NAND2X1_561/Y vdd NAND2X1
XNAND2X1_594 INVX8_5/A INVX1_421/Y gnd NAND2X1_594/Y vdd NAND2X1
XNAND2X1_583 BUFX4_38/Y INVX2_17/A gnd NAND2X1_583/Y vdd NAND2X1
XFILL_9_1 gnd vdd FILL
XFILL_35_3_0 gnd vdd FILL
XFILL_1_3_0 gnd vdd FILL
XFILL_26_3_0 gnd vdd FILL
XOAI21X1_330 NOR2X1_281/A NAND2X1_500/A OAI21X1_330/C gnd AOI21X1_42/B vdd OAI21X1
XFILL_10_7_1 gnd vdd FILL
XOAI21X1_341 NAND3X1_94/Y OAI22X1_10/Y OAI21X1_341/C gnd OAI21X1_341/Y vdd OAI21X1
XOAI21X1_363 MUX2X1_2/Y INVX8_8/A OAI21X1_648/C gnd OAI21X1_411/B vdd OAI21X1
XOAI21X1_352 BUFX4_227/Y OAI21X1_350/Y OR2X2_19/Y gnd OAI21X1_353/B vdd OAI21X1
XOAI21X1_374 OR2X2_24/Y BUFX4_90/Y OAI21X1_375/C gnd AND2X2_27/A vdd OAI21X1
XOAI21X1_385 MUX2X1_2/Y BUFX4_39/Y OAI21X1_385/C gnd MUX2X1_23/B vdd OAI21X1
XOAI21X1_396 BUFX4_41/Y MUX2X1_16/Y OAI21X1_469/C gnd INVX1_366/A vdd OAI21X1
XINVX1_405 INVX1_405/A gnd INVX1_405/Y vdd INVX1
XINVX1_416 NOR2X1_80/Y gnd INVX1_416/Y vdd INVX1
XAND2X2_8 AND2X2_8/A AND2X2_8/B gnd AND2X2_8/Y vdd AND2X2
XINVX1_427 INVX1_427/A gnd INVX1_427/Y vdd INVX1
XINVX1_438 OR2X2_64/B gnd INVX1_438/Y vdd INVX1
XINVX1_449 INVX1_449/A gnd INVX1_449/Y vdd INVX1
XFILL_9_4_0 gnd vdd FILL
XNAND2X1_380 INVX8_5/A OAI21X1_393/Y gnd NAND2X1_380/Y vdd NAND2X1
XNAND2X1_391 AOI21X1_59/Y NAND2X1_377/Y gnd NAND2X1_391/Y vdd NAND2X1
XFILL_17_3_0 gnd vdd FILL
XFILL_42_6_1 gnd vdd FILL
XFILL_41_1_0 gnd vdd FILL
XAOI22X1_3 INVX2_1/Y BUFX2_87/A INVX2_3/A AOI22X1_3/D gnd NAND3X1_2/B vdd AOI22X1
XOAI21X1_160 BUFX4_186/Y INVX1_130/Y OAI21X1_159/Y gnd INVX1_639/A vdd OAI21X1
XOAI21X1_171 BUFX4_14/Y BUFX4_197/Y OAI21X1_829/Y gnd NAND3X1_27/C vdd OAI21X1
XOAI21X1_182 BUFX4_12/Y BUFX4_199/Y OAI21X1_182/C gnd NAND3X1_49/C vdd OAI21X1
XINVX1_224 NOR2X1_9/B gnd INVX1_224/Y vdd INVX1
XINVX1_235 OR2X2_61/A gnd INVX1_235/Y vdd INVX1
XOAI21X1_193 BUFX4_141/Y INVX1_188/Y AOI22X1_8/Y gnd OAI21X1_193/Y vdd OAI21X1
XINVX1_213 INVX1_213/A gnd INVX1_213/Y vdd INVX1
XINVX1_202 INVX1_202/A gnd INVX1_202/Y vdd INVX1
XINVX1_257 MUX2X1_6/A gnd INVX1_257/Y vdd INVX1
XINVX1_246 INVX1_690/A gnd INVX1_246/Y vdd INVX1
XINVX1_268 INVX1_268/A gnd INVX1_268/Y vdd INVX1
XINVX1_279 INVX1_279/A gnd INVX1_279/Y vdd INVX1
XNAND2X1_24 BUFX4_21/Y NAND2X1_24/B gnd OAI21X1_24/C vdd NAND2X1
XNAND2X1_13 BUFX4_17/Y NAND2X1_13/B gnd OAI21X1_13/C vdd NAND2X1
XNAND2X1_35 BUFX4_30/Y NAND2X1_35/B gnd NAND2X1_35/Y vdd NAND2X1
XNAND2X1_68 INVX2_5/A BUFX4_156/Y gnd OAI21X1_66/C vdd NAND2X1
XNAND2X1_46 BUFX4_25/Y NAND2X1_46/B gnd NAND2X1_46/Y vdd NAND2X1
XNAND2X1_57 BUFX4_27/Y NAND2X1_57/B gnd NAND2X1_57/Y vdd NAND2X1
XNAND2X1_79 INVX2_11/A BUFX4_163/Y gnd NAND2X1_79/Y vdd NAND2X1
XFILL_32_1_0 gnd vdd FILL
XFILL_33_6_1 gnd vdd FILL
XAOI21X1_206 INVX2_65/A MUX2X1_55/Y OAI21X1_761/Y gnd AOI21X1_206/Y vdd AOI21X1
XAOI21X1_217 INVX1_480/Y NOR3X1_65/Y BUFX2_57/A gnd AOI21X1_217/Y vdd AOI21X1
XAOI21X1_239 AOI21X1_239/A INVX1_691/Y OAI21X1_913/Y gnd AOI21X1_240/A vdd AOI21X1
XAOI21X1_228 BUFX2_90/A INVX1_575/Y INVX1_577/Y gnd NAND2X1_820/A vdd AOI21X1
XAOI22X1_33 AOI22X1_33/A BUFX4_238/Y BUFX4_256/Y AOI22X1_33/D gnd AOI22X1_33/Y vdd
+ AOI22X1
XAOI22X1_22 AOI22X1_22/A BUFX4_237/Y BUFX4_259/Y AOI22X1_22/D gnd AOI22X1_22/Y vdd
+ AOI22X1
XAOI22X1_11 AOI22X1_11/A BUFX4_237/Y BUFX4_257/Y AOI22X1_11/D gnd AOI22X1_11/Y vdd
+ AOI22X1
XAOI22X1_44 INVX1_350/A BUFX4_231/Y BUFX4_150/Y OR2X2_62/A gnd XNOR2X1_9/A vdd AOI22X1
XAOI22X1_55 INVX1_239/A BUFX4_232/Y BUFX4_146/Y OR2X2_61/A gnd XNOR2X1_37/A vdd AOI22X1
XAOI22X1_66 AOI22X1_66/A AND2X2_12/A AND2X2_11/A INVX1_668/A gnd INVX1_291/A vdd AOI22X1
XAOI22X1_88 AOI22X1_88/A AOI21X1_88/A AOI22X1_88/C AOI22X1_88/D gnd AOI22X1_88/Y vdd
+ AOI22X1
XAOI22X1_99 AOI22X1_99/A AOI22X1_99/B AOI22X1_99/C AOI22X1_99/D gnd AOI22X1_99/Y vdd
+ AOI22X1
XAOI22X1_77 BUFX4_187/Y AOI21X1_69/A AOI21X1_69/C BUFX4_155/Y gnd AOI22X1_77/Y vdd
+ AOI22X1
XNOR3X1_1 NOR3X1_4/A NOR3X1_1/B NOR3X1_4/C gnd NOR3X1_1/Y vdd NOR3X1
XFILL_24_6_1 gnd vdd FILL
XFILL_23_1_0 gnd vdd FILL
XOAI22X1_6 OR2X2_5/Y OAI22X1_6/B OR2X2_6/Y OR2X2_7/Y gnd OAI22X1_6/Y vdd OAI22X1
XFILL_7_7_1 gnd vdd FILL
XFILL_6_2_0 gnd vdd FILL
XFILL_15_6_1 gnd vdd FILL
XFILL_14_1_0 gnd vdd FILL
XDFFPOSX1_309 INVX1_245/A CLKBUF1_25/Y NOR2X1_414/Y gnd vdd DFFPOSX1
XNOR2X1_401 NOR2X1_401/A OAI22X1_46/Y gnd NOR2X1_401/Y vdd NOR2X1
XNOR2X1_434 OR2X2_63/B OR2X2_65/A gnd NOR2X1_434/Y vdd NOR2X1
XNOR2X1_423 INVX1_306/A INVX2_81/Y gnd NOR2X1_423/Y vdd NOR2X1
XNOR2X1_412 INVX2_79/A INVX1_643/Y gnd NOR2X1_412/Y vdd NOR2X1
XNOR2X1_456 INVX2_49/A OR2X2_66/B gnd AND2X2_93/A vdd NOR2X1
XNOR2X1_445 INVX1_325/A INVX2_83/Y gnd NOR2X1_445/Y vdd NOR2X1
XFILL_33_1 gnd vdd FILL
XNOR2X1_467 NOR2X1_3/B NOR3X1_76/A gnd NOR2X1_467/Y vdd NOR2X1
XNOR2X1_478 INVX8_15/Y INVX8_17/Y gnd BUFX4_107/A vdd NOR2X1
XOAI21X1_907 AOI22X1_133/Y INVX1_684/Y OAI21X1_907/C gnd OAI21X1_907/Y vdd OAI21X1
XOAI21X1_929 INVX1_689/A INVX1_709/Y NOR2X1_438/Y gnd OAI21X1_929/Y vdd OAI21X1
XOAI21X1_918 NAND3X1_337/Y INVX1_711/A INVX1_712/A gnd OAI21X1_918/Y vdd OAI21X1
XNAND2X1_913 INVX1_638/Y BUFX4_98/Y gnd NAND3X1_323/C vdd NAND2X1
XINVX2_15 INVX2_15/A gnd INVX2_15/Y vdd INVX2
XINVX2_26 INVX2_26/A gnd INVX2_26/Y vdd INVX2
XNAND2X1_902 NAND2X1_900/Y NAND2X1_902/B gnd NAND2X1_60/B vdd NAND2X1
XINVX2_59 INVX2_59/A gnd INVX2_59/Y vdd INVX2
XINVX2_37 INVX2_37/A gnd INVX2_37/Y vdd INVX2
XINVX2_48 INVX2_48/A gnd INVX2_48/Y vdd INVX2
XNAND2X1_946 INVX1_450/A INVX1_678/Y gnd AND2X2_86/B vdd NAND2X1
XNAND2X1_935 OR2X2_55/A OR2X2_55/B gnd AOI22X1_127/C vdd NAND2X1
XNAND2X1_924 NOR2X1_23/A NOR2X1_411/Y gnd OAI21X1_880/C vdd NAND2X1
XNAND2X1_957 OR2X2_63/A OR2X2_63/B gnd AOI22X1_132/C vdd NAND2X1
XNAND2X1_968 MUX2X1_3/B INVX1_676/Y gnd OAI21X1_912/C vdd NAND2X1
XNAND2X1_979 OR2X2_54/A INVX1_702/Y gnd NAND2X1_979/Y vdd NAND2X1
XFILL_30_4_1 gnd vdd FILL
XDFFPOSX1_128 DFFPOSX1_16/D CLKBUF1_18/Y INVX2_8/A gnd vdd DFFPOSX1
XDFFPOSX1_117 AND2X2_99/B CLKBUF1_22/Y INVX2_51/A gnd vdd DFFPOSX1
XDFFPOSX1_106 INVX1_219/A CLKBUF1_61/Y OAI21X1_153/C gnd vdd DFFPOSX1
XDFFPOSX1_139 DFFPOSX1_27/D CLKBUF1_42/Y INVX1_268/A gnd vdd DFFPOSX1
XNAND2X1_209 INVX1_317/A MUX2X1_46/B gnd AND2X2_59/B vdd NAND2X1
XFILL_37_0_0 gnd vdd FILL
XFILL_38_5_1 gnd vdd FILL
XBUFX4_160 NOR2X1_2/Y gnd BUFX4_160/Y vdd BUFX4
XBUFX4_182 OR2X2_2/Y gnd BUFX4_182/Y vdd BUFX4
XBUFX4_171 BUFX4_171/A gnd BUFX4_171/Y vdd BUFX4
XNOR2X1_220 NOR2X1_220/A BUFX4_275/Y gnd AOI21X1_80/B vdd NOR2X1
XNOR2X1_242 INVX2_45/A MUX2X1_10/Y gnd OAI22X1_24/D vdd NOR2X1
XNOR2X1_231 NOR2X1_227/Y NOR2X1_231/B gnd NOR2X1_231/Y vdd NOR2X1
XBUFX4_193 BUFX4_194/A gnd BUFX4_193/Y vdd BUFX4
XNOR2X1_253 NOR2X1_253/A NOR2X1_253/B gnd NOR2X1_254/B vdd NOR2X1
XNOR2X1_275 OR2X2_32/B INVX2_61/Y gnd NOR2X1_275/Y vdd NOR2X1
XNOR2X1_264 OR2X2_31/B OR2X2_23/A gnd AND2X2_43/A vdd NOR2X1
XNOR2X1_297 INVX2_42/A MUX2X1_7/Y gnd OAI22X1_37/B vdd NOR2X1
XNOR2X1_286 BUFX4_86/Y AND2X2_46/Y gnd NOR2X1_286/Y vdd NOR2X1
XOAI21X1_704 NOR2X1_340/Y NOR2X1_339/Y BUFX4_128/Y gnd OAI21X1_704/Y vdd OAI21X1
XOAI21X1_715 INVX1_420/Y INVX8_5/A NAND2X1_580/Y gnd MUX2X1_49/A vdd OAI21X1
XFILL_21_4_1 gnd vdd FILL
XOAI21X1_748 NOR2X1_359/Y NOR2X1_360/Y NOR3X1_56/Y gnd OAI21X1_748/Y vdd OAI21X1
XOAI21X1_726 OAI22X1_44/C INVX8_4/A NAND2X1_585/Y gnd AND2X2_66/A vdd OAI21X1
XOAI21X1_737 OAI21X1_736/Y INVX8_5/A OAI21X1_737/C gnd NAND2X1_590/B vdd OAI21X1
XOAI21X1_759 INVX8_7/A OAI21X1_758/Y NOR3X1_56/Y gnd OAI21X1_759/Y vdd OAI21X1
XOAI21X1_1050 BUFX4_64/Y BUFX4_68/Y AOI22X1_166/Y gnd OAI21X1_1050/Y vdd OAI21X1
XOAI21X1_1061 AND2X2_101/Y NOR2X1_488/B NOR2X1_487/Y gnd OR2X2_70/A vdd OAI21X1
XNAND2X1_721 OAI21X1_69/Y BUFX4_135/Y gnd NAND2X1_723/A vdd NAND2X1
XNAND2X1_710 AOI21X1_224/Y NAND2X1_710/B gnd NOR2X1_402/B vdd NAND2X1
XNAND2X1_732 NAND2X1_730/Y NAND2X1_732/B gnd NAND2X1_8/B vdd NAND2X1
XNAND2X1_754 OAI21X1_80/Y BUFX4_135/Y gnd NAND2X1_754/Y vdd NAND2X1
XNAND2X1_743 INVX1_525/Y BUFX4_202/Y gnd NAND2X1_743/Y vdd NAND2X1
XNAND2X1_787 OAI21X1_91/Y BUFX4_135/Y gnd NAND2X1_787/Y vdd NAND2X1
XNAND2X1_765 NAND2X1_765/A NAND2X1_765/B gnd NAND2X1_19/B vdd NAND2X1
XNAND2X1_776 INVX1_547/Y BUFX4_201/Y gnd NAND3X1_235/C vdd NAND2X1
XFILL_4_5_1 gnd vdd FILL
XFILL_28_0_0 gnd vdd FILL
XFILL_29_5_1 gnd vdd FILL
XNAND2X1_798 NAND2X1_798/A NAND2X1_798/B gnd NAND2X1_30/B vdd NAND2X1
XFILL_3_0_0 gnd vdd FILL
XINVX8_2 INVX8_2/A gnd INVX8_2/Y vdd INVX8
XFILL_12_4_1 gnd vdd FILL
XBUFX4_11 BUFX4_9/A gnd BUFX4_11/Y vdd BUFX4
XBUFX4_44 INVX8_8/Y gnd BUFX4_44/Y vdd BUFX4
XBUFX4_22 BUFX4_22/A gnd BUFX4_22/Y vdd BUFX4
XBUFX4_33 BUFX4_37/A gnd BUFX4_33/Y vdd BUFX4
XBUFX4_77 INVX8_6/Y gnd BUFX4_77/Y vdd BUFX4
XBUFX4_55 INVX8_3/Y gnd BUFX4_55/Y vdd BUFX4
XBUFX4_66 BUFX4_65/A gnd BUFX4_66/Y vdd BUFX4
XBUFX4_88 BUFX4_88/A gnd BUFX4_88/Y vdd BUFX4
XFILL_19_0_0 gnd vdd FILL
XBUFX4_99 BUFX4_99/A gnd BUFX4_99/Y vdd BUFX4
XNAND3X1_360 NAND3X1_360/A NAND3X1_360/B OAI21X1_968/C gnd NAND3X1_360/Y vdd NAND3X1
XOR2X2_14 OR2X2_14/A OR2X2_14/B gnd OR2X2_14/Y vdd OR2X2
XOR2X2_47 OR2X2_47/A OR2X2_47/B gnd OR2X2_47/Y vdd OR2X2
XOR2X2_58 MUX2X1_7/B OR2X2_58/B gnd OR2X2_58/Y vdd OR2X2
XOR2X2_36 OR2X2_36/A OR2X2_36/B gnd OR2X2_36/Y vdd OR2X2
XOR2X2_25 OR2X2_25/A OR2X2_25/B gnd OR2X2_25/Y vdd OR2X2
XOR2X2_7 OR2X2_5/B OR2X2_7/B gnd OR2X2_7/Y vdd OR2X2
XOR2X2_69 OR2X2_69/A OR2X2_69/B gnd OR2X2_69/Y vdd OR2X2
XXNOR2X1_9 XNOR2X1_9/A INVX2_7/Y gnd XNOR2X1_9/Y vdd XNOR2X1
XINVX8_14 INVX8_14/A gnd INVX8_14/Y vdd INVX8
XOAI21X1_501 OAI22X1_17/B AOI22X1_88/D AOI22X1_88/A gnd AOI21X1_91/A vdd OAI21X1
XOAI21X1_512 AOI21X1_74/Y NAND2X1_474/Y AOI21X1_96/Y gnd OAI21X1_513/C vdd OAI21X1
XOAI21X1_523 OAI21X1_523/A INVX8_7/A OAI21X1_523/C gnd AOI22X1_91/B vdd OAI21X1
XINVX1_9 gnd gnd INVX1_9/Y vdd INVX1
XOAI21X1_545 NOR2X1_271/Y NOR2X1_270/Y BUFX4_128/Y gnd OAI21X1_545/Y vdd OAI21X1
XOAI21X1_556 INVX8_5/A INVX1_396/A NAND2X1_503/Y gnd INVX1_398/A vdd OAI21X1
XOAI21X1_534 BUFX4_57/Y INVX1_389/Y OAI21X1_534/C gnd NOR2X1_256/B vdd OAI21X1
XOAI21X1_567 AND2X2_45/Y INVX4_5/Y OAI21X1_567/C gnd OAI21X1_568/A vdd OAI21X1
XOAI21X1_589 OAI22X1_7/A AOI22X1_70/C OAI22X1_36/B gnd OAI21X1_589/Y vdd OAI21X1
XOAI21X1_578 OAI22X1_30/C NAND2X1_523/Y OAI21X1_578/C gnd NOR2X1_290/B vdd OAI21X1
XINVX1_609 INVX1_609/A gnd INVX1_609/Y vdd INVX1
XDFFPOSX1_481 XOR2X1_8/B CLKBUF1_33/Y NAND3X1_25/Y gnd vdd DFFPOSX1
XDFFPOSX1_492 BUFX2_59/A CLKBUF1_45/Y NAND3X1_47/Y gnd vdd DFFPOSX1
XDFFPOSX1_470 NAND3X1_66/A CLKBUF1_36/Y BUFX2_69/A gnd vdd DFFPOSX1
XNAND2X1_540 BUFX4_126/Y NAND2X1_540/B gnd INVX1_400/A vdd NAND2X1
XNAND2X1_551 INVX8_4/A MUX2X1_40/Y gnd NAND2X1_551/Y vdd NAND2X1
XNAND2X1_562 INVX1_412/A AOI22X1_69/C gnd INVX2_70/A vdd NAND2X1
XNAND2X1_595 INVX8_4/A NAND2X1_595/B gnd NAND2X1_595/Y vdd NAND2X1
XNAND2X1_573 BUFX4_38/Y INVX2_50/A gnd OAI21X1_699/C vdd NAND2X1
XNAND2X1_584 BUFX4_225/Y INVX1_421/Y gnd OAI21X1_725/C vdd NAND2X1
XFILL_35_3_1 gnd vdd FILL
XNAND3X1_190 INVX1_503/Y BUFX4_206/Y BUFX4_33/Y gnd NAND3X1_190/Y vdd NAND3X1
XFILL_1_3_1 gnd vdd FILL
XFILL_26_3_1 gnd vdd FILL
XOAI21X1_320 INVX1_341/Y INVX4_4/A NAND2X1_277/Y gnd MUX2X1_31/B vdd OAI21X1
XOAI21X1_331 OAI22X1_38/B AOI22X1_99/C AOI22X1_99/B gnd AOI21X1_42/C vdd OAI21X1
XOAI21X1_342 BUFX4_44/Y MUX2X1_24/B OAI21X1_342/C gnd OAI21X1_343/A vdd OAI21X1
XOAI21X1_353 INVX8_4/A OAI21X1_353/B OAI21X1_353/C gnd AOI21X1_52/B vdd OAI21X1
XOAI21X1_364 INVX2_53/Y INVX8_8/A OAI21X1_364/C gnd INVX1_354/A vdd OAI21X1
XOAI21X1_386 INVX1_362/Y BUFX4_228/Y NAND2X1_370/Y gnd OAI21X1_390/B vdd OAI21X1
XOAI21X1_397 INVX1_366/Y INVX8_5/A OAI21X1_397/C gnd MUX2X1_27/B vdd OAI21X1
XINVX1_417 INVX1_417/A gnd INVX1_417/Y vdd INVX1
XINVX1_406 INVX1_406/A gnd INVX1_406/Y vdd INVX1
XOAI21X1_375 NOR2X1_176/Y NOR2X1_178/A OAI21X1_375/C gnd OAI21X1_376/C vdd OAI21X1
XAND2X2_9 AND2X2_1/A AND2X2_1/B gnd AND2X2_9/Y vdd AND2X2
XINVX1_439 OR2X2_62/B gnd INVX1_439/Y vdd INVX1
XINVX1_428 INVX1_428/A gnd INVX1_428/Y vdd INVX1
XFILL_9_4_1 gnd vdd FILL
XNAND2X1_370 BUFX4_223/Y MUX2X1_23/B gnd NAND2X1_370/Y vdd NAND2X1
XNAND2X1_381 BUFX4_41/Y MUX2X1_31/B gnd NAND2X1_381/Y vdd NAND2X1
XNAND2X1_392 BUFX4_82/Y NOR2X1_188/Y gnd INVX1_370/A vdd NAND2X1
XFILL_17_3_1 gnd vdd FILL
XFILL_41_1_1 gnd vdd FILL
XAOI22X1_4 INVX2_1/Y INVX1_495/A INVX2_2/A AOI22X1_4/D gnd AND2X2_4/B vdd AOI22X1
XOAI21X1_172 BUFX4_14/Y BUFX4_197/Y OAI21X1_832/Y gnd NAND3X1_29/C vdd OAI21X1
XOAI21X1_183 BUFX4_16/Y BUFX4_198/Y OAI21X1_854/Y gnd NAND3X1_51/C vdd OAI21X1
XOAI21X1_161 BUFX4_13/Y BUFX4_196/Y OAI21X1_161/C gnd AOI21X1_1/B vdd OAI21X1
XOAI21X1_150 BUFX4_185/Y INVX1_125/Y OAI21X1_150/C gnd INVX1_556/A vdd OAI21X1
XOAI21X1_194 OR2X2_4/A INVX1_192/Y AOI22X1_9/Y gnd OAI21X1_194/Y vdd OAI21X1
XINVX1_203 INVX1_203/A gnd INVX1_203/Y vdd INVX1
XINVX1_214 INVX1_214/A gnd INVX1_214/Y vdd INVX1
XINVX1_225 INVX1_225/A gnd NOR2X1_20/B vdd INVX1
XINVX1_247 INVX1_247/A gnd INVX1_247/Y vdd INVX1
XINVX1_258 INVX1_258/A gnd INVX1_258/Y vdd INVX1
XINVX1_236 NOR2X1_6/A gnd INVX1_236/Y vdd INVX1
XINVX1_269 INVX1_269/A gnd INVX1_269/Y vdd INVX1
XNAND2X1_25 BUFX4_21/Y NAND2X1_25/B gnd OAI21X1_25/C vdd NAND2X1
XNAND2X1_14 BUFX4_17/Y NAND2X1_14/B gnd OAI21X1_14/C vdd NAND2X1
XNAND2X1_47 BUFX4_28/Y NAND2X1_47/B gnd OAI21X1_47/C vdd NAND2X1
XNAND2X1_58 BUFX4_29/Y NAND2X1_58/B gnd NAND2X1_58/Y vdd NAND2X1
XNAND2X1_36 BUFX4_31/Y NAND2X1_36/B gnd NAND2X1_36/Y vdd NAND2X1
XNAND2X1_69 INVX2_6/A BUFX4_160/Y gnd NAND2X1_69/Y vdd NAND2X1
XAOI21X1_207 NOR2X1_85/B INVX2_71/A NOR2X1_87/Y gnd OAI21X1_763/C vdd AOI21X1
XFILL_32_1_1 gnd vdd FILL
XAOI21X1_229 BUFX2_87/A INVX1_640/Y OAI21X1_874/Y gnd NAND3X1_324/C vdd AOI21X1
XAOI21X1_218 AND2X2_78/A NOR3X1_65/Y BUFX2_59/A gnd AOI21X1_218/Y vdd AOI21X1
XAOI22X1_23 AOI22X1_23/A BUFX4_236/Y BUFX4_258/Y AOI22X1_23/D gnd AOI22X1_23/Y vdd
+ AOI22X1
XAOI22X1_12 AOI22X1_12/A BUFX4_237/Y BUFX4_259/Y AOI22X1_12/D gnd AOI22X1_12/Y vdd
+ AOI22X1
XAOI22X1_56 MUX2X1_2/A BUFX4_231/Y BUFX4_147/Y MUX2X1_2/B gnd OR2X2_10/A vdd AOI22X1
XAOI22X1_45 INVX1_242/A BUFX4_232/Y BUFX4_147/Y INVX2_85/A gnd AOI22X1_45/Y vdd AOI22X1
XAOI22X1_34 AOI22X1_34/A BUFX4_237/Y BUFX4_257/Y AOI22X1_34/D gnd AOI22X1_34/Y vdd
+ AOI22X1
XAOI22X1_89 AOI22X1_89/A AOI22X1_89/B AOI22X1_89/C AOI22X1_89/D gnd AOI21X1_96/A vdd
+ AOI22X1
XAOI22X1_78 INVX8_11/Y AOI22X1_78/B AOI21X1_64/A OR2X2_24/Y gnd AOI22X1_78/Y vdd AOI22X1
XAOI22X1_67 AOI22X1_67/A BUFX4_233/Y BUFX4_148/Y INVX1_667/A gnd NOR2X1_65/B vdd AOI22X1
XNOR3X1_2 NOR3X1_9/A NOR3X1_2/B NOR3X1_9/C gnd NOR3X1_2/Y vdd NOR3X1
XFILL_23_1_1 gnd vdd FILL
XOAI22X1_7 OAI22X1_7/A OAI22X1_7/B OAI22X1_7/C OAI22X1_7/D gnd OAI22X1_7/Y vdd OAI22X1
XFILL_6_2_1 gnd vdd FILL
XFILL_14_1_1 gnd vdd FILL
XNOR2X1_413 INVX1_648/Y BUFX4_260/Y gnd NOR2X1_413/Y vdd NOR2X1
XNOR2X1_424 NOR2X1_424/A NOR2X1_424/B gnd NOR2X1_424/Y vdd NOR2X1
XNOR2X1_402 NOR2X1_402/A NOR2X1_402/B gnd BUFX4_37/A vdd NOR2X1
XNOR2X1_435 OR2X2_61/B INVX1_688/Y gnd NOR2X1_435/Y vdd NOR2X1
XNOR2X1_457 OR2X2_64/A INVX1_683/Y gnd NOR2X1_457/Y vdd NOR2X1
XNOR2X1_446 INVX1_454/A INVX1_698/Y gnd NOR2X1_446/Y vdd NOR2X1
XFILL_33_2 gnd vdd FILL
XNOR2X1_468 AND2X2_99/B INVX8_15/A gnd INVX2_90/A vdd NOR2X1
XFILL_26_1 gnd vdd FILL
XNOR2X1_479 INVX1_733/Y BUFX4_118/Y gnd NOR2X1_479/Y vdd NOR2X1
XOAI21X1_908 NAND2X1_961/Y AOI21X1_236/Y AOI21X1_237/Y gnd OAI21X1_908/Y vdd OAI21X1
XOAI21X1_919 NOR2X1_423/Y AND2X2_82/B AND2X2_82/A gnd OAI21X1_919/Y vdd OAI21X1
XINVX2_16 INVX2_16/A gnd INVX2_16/Y vdd INVX2
XINVX2_27 INVX2_27/A gnd INVX2_27/Y vdd INVX2
XNAND2X1_903 OAI21X1_93/Y BUFX4_62/Y gnd NAND2X1_903/Y vdd NAND2X1
XINVX2_38 INVX2_38/A gnd INVX2_38/Y vdd INVX2
XINVX2_49 INVX2_49/A gnd INVX2_49/Y vdd INVX2
XNAND2X1_936 INVX1_306/A INVX2_81/Y gnd AND2X2_82/A vdd NAND2X1
XNAND2X1_925 INVX1_643/A NOR2X1_22/B gnd NAND2X1_925/Y vdd NAND2X1
XNAND2X1_914 NAND2X1_912/Y NAND2X1_914/B gnd NAND2X1_64/B vdd NAND2X1
XNAND2X1_958 OR2X2_64/A INVX1_683/Y gnd INVX1_684/A vdd NAND2X1
XNAND2X1_947 MUX2X1_6/B INVX1_449/A gnd NAND2X1_947/Y vdd NAND2X1
XNAND2X1_969 INVX1_664/A INVX1_665/Y gnd NAND2X1_970/A vdd NAND2X1
XDFFPOSX1_118 INVX8_15/A CLKBUF1_38/Y INVX2_49/A gnd vdd DFFPOSX1
XDFFPOSX1_107 INVX1_220/A CLKBUF1_61/Y OAI21X1_155/C gnd vdd DFFPOSX1
XDFFPOSX1_129 DFFPOSX1_17/D CLKBUF1_2/Y INVX1_253/A gnd vdd DFFPOSX1
XCLKBUF1_1 BUFX4_6/Y gnd CLKBUF1_1/Y vdd CLKBUF1
XBUFX4_150 BUFX4_148/A gnd BUFX4_150/Y vdd BUFX4
XBUFX4_161 NOR2X1_2/Y gnd BUFX4_161/Y vdd BUFX4
XFILL_37_0_1 gnd vdd FILL
XBUFX4_172 BUFX4_171/A gnd BUFX4_172/Y vdd BUFX4
XNOR2X1_221 INVX8_7/A AND2X2_34/A gnd OAI22X1_17/D vdd NOR2X1
XNOR2X1_232 NOR2X1_232/A AOI21X1_87/Y gnd NOR2X1_232/Y vdd NOR2X1
XNOR2X1_243 INVX1_342/A MUX2X1_15/Y gnd OAI22X1_22/B vdd NOR2X1
XNOR2X1_210 AOI21X1_64/A NOR2X1_210/B gnd NOR2X1_210/Y vdd NOR2X1
XBUFX4_183 OR2X2_2/Y gnd BUFX4_183/Y vdd BUFX4
XBUFX4_194 BUFX4_194/A gnd BUFX4_194/Y vdd BUFX4
XNOR2X1_254 NOR2X1_254/A NOR2X1_254/B gnd NOR2X1_254/Y vdd NOR2X1
XNOR2X1_276 BUFX4_274/Y NOR2X1_275/Y gnd NOR2X1_276/Y vdd NOR2X1
XNOR2X1_265 INVX8_9/A NOR2X1_256/B gnd NOR2X1_265/Y vdd NOR2X1
XNOR2X1_287 INVX2_41/Y MUX2X1_37/A gnd OAI22X1_31/C vdd NOR2X1
XNOR2X1_298 INVX8_6/A OR2X2_23/Y gnd INVX2_65/A vdd NOR2X1
XOAI21X1_705 INVX1_387/A BUFX4_128/Y OAI21X1_704/Y gnd AND2X2_63/A vdd OAI21X1
XOAI21X1_727 AND2X2_66/Y AND2X2_67/Y BUFX4_129/Y gnd OAI21X1_728/C vdd OAI21X1
XOAI21X1_738 MUX2X1_47/Y MUX2X1_49/S OAI21X1_738/C gnd MUX2X1_50/B vdd OAI21X1
XOAI21X1_716 MUX2X1_49/Y INVX8_3/A NAND2X1_579/Y gnd NOR2X1_344/B vdd OAI21X1
XOAI21X1_749 INVX8_12/Y NOR2X1_85/A OAI21X1_749/C gnd NOR2X1_361/B vdd OAI21X1
XOAI21X1_1040 BUFX4_66/Y BUFX4_71/Y AOI22X1_156/Y gnd OAI21X1_1040/Y vdd OAI21X1
XOAI21X1_1051 BUFX4_66/Y BUFX4_71/Y AOI22X1_167/Y gnd OAI21X1_1051/Y vdd OAI21X1
XOAI21X1_1062 AOI21X1_263/A INVX2_87/Y AND2X2_101/B gnd OAI21X1_1062/Y vdd OAI21X1
XNAND2X1_711 NAND2X1_711/A NAND2X1_711/B gnd NAND2X1_1/A vdd NAND2X1
XNAND2X1_700 INVX2_73/A INVX1_497/Y gnd NAND3X1_187/A vdd NAND2X1
XNAND2X1_733 OAI21X1_73/Y BUFX4_135/Y gnd NAND2X1_733/Y vdd NAND2X1
XNAND2X1_744 NAND2X1_742/Y NAND2X1_744/B gnd NAND2X1_12/B vdd NAND2X1
XNAND2X1_755 INVX1_533/Y BUFX4_201/Y gnd NAND3X1_221/C vdd NAND2X1
XNAND2X1_722 INVX1_511/Y BUFX4_201/Y gnd NAND3X1_199/C vdd NAND2X1
XNAND2X1_788 INVX1_555/Y BUFX4_203/Y gnd NAND3X1_243/C vdd NAND2X1
XNAND2X1_766 OAI21X1_84/Y BUFX4_133/Y gnd NAND2X1_768/A vdd NAND2X1
XNAND2X1_777 NAND2X1_777/A NAND2X1_777/B gnd NAND2X1_23/B vdd NAND2X1
XNAND2X1_799 OAI21X1_95/Y BUFX4_132/Y gnd NAND2X1_799/Y vdd NAND2X1
XFILL_3_0_1 gnd vdd FILL
XFILL_28_0_1 gnd vdd FILL
XINVX8_3 INVX8_3/A gnd INVX8_3/Y vdd INVX8
XFILL_40_7_0 gnd vdd FILL
XBUFX4_12 BUFX4_13/A gnd BUFX4_12/Y vdd BUFX4
XBUFX4_23 BUFX4_22/A gnd BUFX4_23/Y vdd BUFX4
XBUFX4_34 BUFX4_37/A gnd BUFX4_34/Y vdd BUFX4
XBUFX4_78 INVX8_6/Y gnd BUFX4_78/Y vdd BUFX4
XBUFX4_56 INVX8_3/Y gnd BUFX4_56/Y vdd BUFX4
XBUFX4_45 BUFX4_46/A gnd BUFX4_45/Y vdd BUFX4
XBUFX4_67 BUFX4_65/A gnd BUFX4_67/Y vdd BUFX4
XBUFX4_89 BUFX4_88/A gnd INVX8_10/A vdd BUFX4
XFILL_19_0_1 gnd vdd FILL
XFILL_31_7_0 gnd vdd FILL
XNAND3X1_350 NOR3X1_75/Y BUFX4_11/Y NOR3X1_76/Y gnd AOI21X1_259/B vdd NAND3X1
XNAND3X1_361 NAND3X1_361/A NAND3X1_361/B NAND3X1_361/C gnd NAND3X1_361/Y vdd NAND3X1
XOR2X2_15 OR2X2_15/A OR2X2_15/B gnd OR2X2_15/Y vdd OR2X2
XOR2X2_37 OR2X2_37/A OR2X2_37/B gnd OR2X2_37/Y vdd OR2X2
XOR2X2_26 OR2X2_26/A INVX8_3/A gnd OR2X2_27/B vdd OR2X2
XOR2X2_48 OR2X2_48/A OR2X2_48/B gnd OR2X2_48/Y vdd OR2X2
XOR2X2_59 OR2X2_59/A OR2X2_59/B gnd OR2X2_59/Y vdd OR2X2
XOR2X2_8 OR2X2_8/A OR2X2_8/B gnd OR2X2_8/Y vdd OR2X2
XINVX8_15 INVX8_15/A gnd INVX8_15/Y vdd INVX8
XFILL_22_7_0 gnd vdd FILL
XOAI21X1_513 OAI22X1_24/C OAI22X1_24/D OAI21X1_513/C gnd AOI22X1_90/A vdd OAI21X1
XOAI21X1_502 AND2X2_37/Y AOI22X1_89/D AOI22X1_89/A gnd AOI21X1_91/C vdd OAI21X1
XOAI21X1_546 OR2X2_41/A INVX8_3/A INVX8_7/A gnd OAI21X1_546/Y vdd OAI21X1
XOAI21X1_557 INVX8_4/A INVX1_398/A NAND2X1_502/Y gnd NOR2X1_323/B vdd OAI21X1
XOAI21X1_524 INVX1_388/Y OAI21X1_523/A OAI21X1_524/C gnd AOI22X1_91/C vdd OAI21X1
XOAI21X1_535 AND2X2_42/Y OR2X2_24/B INVX2_59/A gnd OAI21X1_535/Y vdd OAI21X1
XOAI21X1_568 OAI21X1_568/A AOI21X1_118/Y AOI21X1_119/Y gnd NOR2X1_284/A vdd OAI21X1
XOAI21X1_579 MUX2X1_28/Y BUFX4_58/Y BUFX4_129/Y gnd AOI21X1_124/C vdd OAI21X1
XDFFPOSX1_482 BUFX2_49/A CLKBUF1_7/Y NAND3X1_27/Y gnd vdd DFFPOSX1
XDFFPOSX1_460 NAND3X1_46/A CLKBUF1_45/Y BUFX2_59/A gnd vdd DFFPOSX1
XDFFPOSX1_471 NAND3X1_68/A CLKBUF1_27/Y BUFX2_70/A gnd vdd DFFPOSX1
XNAND2X1_530 INVX2_36/Y INVX2_53/Y gnd NAND2X1_530/Y vdd NAND2X1
XDFFPOSX1_493 BUFX2_60/A CLKBUF1_35/Y NAND3X1_49/Y gnd vdd DFFPOSX1
XNAND2X1_541 BUFX4_216/Y MUX2X1_45/B gnd OAI21X1_621/C vdd NAND2X1
XNAND2X1_563 INVX8_7/A NOR2X1_229/Y gnd AOI21X1_170/A vdd NAND2X1
XNAND2X1_552 MUX2X1_54/B BUFX4_81/Y gnd INVX1_425/A vdd NAND2X1
XNAND2X1_585 INVX8_4/A MUX2X1_45/A gnd NAND2X1_585/Y vdd NAND2X1
XNAND2X1_574 BUFX4_225/Y OAI21X1_725/B gnd OAI21X1_700/C vdd NAND2X1
XNAND2X1_596 NOR2X1_85/B BUFX4_152/Y gnd OAI21X1_749/C vdd NAND2X1
XFILL_13_7_0 gnd vdd FILL
XNAND3X1_180 BUFX2_44/A INVX2_72/A BUFX2_46/A gnd NOR2X1_382/B vdd NAND3X1
XNAND3X1_191 BUFX4_220/Y NAND3X1_190/Y NAND3X1_191/C gnd NAND2X1_711/B vdd NAND3X1
XOAI21X1_332 AOI21X1_43/Y NOR2X1_143/A AOI21X1_39/Y gnd AOI21X1_46/B vdd OAI21X1
XOAI21X1_321 INVX1_343/Y INVX4_4/A OAI21X1_321/C gnd MUX2X1_30/B vdd OAI21X1
XOAI21X1_310 INVX1_333/Y INVX4_4/A OAI21X1_310/C gnd MUX2X1_37/A vdd OAI21X1
XOAI21X1_354 INVX8_3/A OAI21X1_354/B AOI21X1_52/Y gnd AOI21X1_57/A vdd OAI21X1
XOAI21X1_365 BUFX4_223/Y OAI21X1_411/B NAND2X1_341/Y gnd NAND2X1_342/B vdd OAI21X1
XOAI21X1_343 OAI21X1_343/A BUFX4_223/Y BUFX4_215/Y gnd OAI21X1_346/B vdd OAI21X1
XINVX1_407 INVX1_407/A gnd INVX1_407/Y vdd INVX1
XOAI21X1_398 INVX8_4/A OAI21X1_394/Y OAI21X1_398/C gnd OAI21X1_398/Y vdd OAI21X1
XOAI21X1_376 OAI22X1_30/A NOR2X1_299/B OAI21X1_376/C gnd AOI21X1_56/C vdd OAI21X1
XOAI21X1_387 INVX2_50/Y BUFX4_38/Y NAND2X1_371/Y gnd INVX1_363/A vdd OAI21X1
XINVX1_418 INVX1_418/A gnd INVX1_418/Y vdd INVX1
XINVX1_429 INVX1_429/A gnd INVX1_429/Y vdd INVX1
XDFFPOSX1_290 NOR2X1_6/B CLKBUF1_34/Y NAND3X1_7/Y gnd vdd DFFPOSX1
XXOR2X1_10 OR2X2_49/B INVX2_3/A gnd XOR2X1_10/Y vdd XOR2X1
XNAND2X1_360 BUFX4_80/Y INVX1_360/Y gnd OAI22X1_30/A vdd NAND2X1
XNAND2X1_371 BUFX4_38/Y MUX2X1_46/B gnd NAND2X1_371/Y vdd NAND2X1
XNAND2X1_382 INVX8_5/A NAND2X1_416/B gnd OAI21X1_397/C vdd NAND2X1
XNAND2X1_393 MUX2X1_47/S MUX2X1_14/Y gnd AOI21X1_69/A vdd NAND2X1
XFILL_36_6_0 gnd vdd FILL
XFILL_2_6_0 gnd vdd FILL
XFILL_27_6_0 gnd vdd FILL
XFILL_10_5_0 gnd vdd FILL
XOAI21X1_140 BUFX4_185/Y INVX1_120/Y OAI21X1_139/Y gnd INVX1_619/A vdd OAI21X1
XAOI22X1_5 INVX2_3/Y OR2X2_49/B INVX2_1/A INVX1_136/Y gnd AOI22X1_5/Y vdd AOI22X1
XOAI21X1_173 BUFX4_14/Y BUFX4_197/Y OAI21X1_173/C gnd NAND3X1_31/C vdd OAI21X1
XOAI21X1_162 BUFX4_13/Y BUFX4_196/Y OAI21X1_816/Y gnd AOI21X1_2/B vdd OAI21X1
XOAI21X1_151 BUFX4_269/Y BUFX4_192/Y OAI21X1_151/C gnd OAI21X1_152/C vdd OAI21X1
XOAI21X1_184 BUFX4_16/Y BUFX4_198/Y OAI21X1_856/Y gnd NAND3X1_53/C vdd OAI21X1
XINVX1_226 NOR2X1_14/A gnd INVX1_226/Y vdd INVX1
XOAI21X1_195 BUFX4_144/Y INVX1_193/Y AOI22X1_10/Y gnd OAI21X1_195/Y vdd OAI21X1
XINVX1_215 INVX1_215/A gnd INVX1_215/Y vdd INVX1
XINVX1_204 INVX1_204/A gnd INVX1_204/Y vdd INVX1
XINVX1_259 NOR2X1_41/Y gnd INVX1_259/Y vdd INVX1
XINVX1_248 INVX1_248/A gnd INVX1_248/Y vdd INVX1
XINVX1_237 OR2X2_1/B gnd NOR3X1_47/C vdd INVX1
XNAND2X1_15 BUFX4_19/Y NAND2X1_15/B gnd OAI21X1_15/C vdd NAND2X1
XNAND2X1_26 BUFX4_17/Y NAND2X1_26/B gnd OAI21X1_26/C vdd NAND2X1
XNAND2X1_37 BUFX4_28/Y NAND2X1_37/B gnd OAI21X1_37/C vdd NAND2X1
XNAND2X1_48 BUFX4_25/Y NAND2X1_48/B gnd NAND2X1_48/Y vdd NAND2X1
XNAND2X1_59 BUFX4_25/Y NAND2X1_59/B gnd OAI21X1_59/C vdd NAND2X1
XNAND2X1_190 INVX1_296/Y NOR2X1_65/B gnd AND2X2_19/B vdd NAND2X1
XFILL_18_6_0 gnd vdd FILL
XAOI21X1_219 BUFX2_61/A NOR2X1_392/B BUFX2_62/A gnd AOI21X1_219/Y vdd AOI21X1
XAOI21X1_208 OAI21X1_763/C AOI21X1_208/B INVX2_28/Y gnd NOR2X1_370/B vdd AOI21X1
XAOI22X1_13 AOI22X1_13/A AOI22X1_9/B OR2X2_3/A AOI22X1_13/D gnd AOI22X1_13/Y vdd AOI22X1
XAOI22X1_24 AOI22X1_24/A OR2X2_3/B BUFX4_257/Y AOI22X1_24/D gnd AOI22X1_24/Y vdd AOI22X1
XAOI22X1_46 INVX1_251/A BUFX4_231/Y BUFX4_147/Y INVX1_689/A gnd XNOR2X1_16/A vdd AOI22X1
XAOI22X1_57 AOI22X1_57/A BUFX4_232/Y BUFX4_146/Y OR2X2_56/A gnd OR2X2_12/A vdd AOI22X1
XAOI22X1_35 AOI22X1_35/A BUFX4_237/Y BUFX4_259/Y AOI22X1_35/D gnd AOI22X1_35/Y vdd
+ AOI22X1
XAOI22X1_79 AOI22X1_79/A AOI21X1_64/Y BUFX4_154/Y AOI22X1_79/D gnd AOI22X1_79/Y vdd
+ AOI22X1
XAOI22X1_68 AOI22X1_68/A AND2X2_12/A AND2X2_11/A INVX1_664/A gnd XNOR2X1_48/A vdd
+ AOI22X1
XNOR3X1_3 NOR3X1_3/A NOR3X1_3/B NOR3X1_4/C gnd NOR3X1_3/Y vdd NOR3X1
XOAI22X1_8 OAI22X1_8/A OAI22X1_8/B OAI22X1_8/C OAI22X1_8/D gnd OAI22X1_8/Y vdd OAI22X1
XFILL_42_4_0 gnd vdd FILL
XAOI21X1_90 INVX4_6/Y INVX1_385/A AOI21X1_90/C gnd AOI21X1_90/Y vdd AOI21X1
XNOR2X1_403 XOR2X1_12/Y XOR2X1_13/Y gnd NOR2X1_403/Y vdd NOR2X1
XNOR2X1_425 NOR2X1_425/A NOR2X1_425/B gnd AND2X2_83/A vdd NOR2X1
XNOR2X1_414 INVX1_649/Y BUFX4_260/Y gnd NOR2X1_414/Y vdd NOR2X1
XNOR2X1_436 OR2X2_60/B INVX2_85/Y gnd NOR2X1_436/Y vdd NOR2X1
XNOR2X1_458 INVX1_685/A INVX1_707/Y gnd NOR2X1_458/Y vdd NOR2X1
XNOR2X1_447 INVX1_459/A INVX2_82/Y gnd INVX1_699/A vdd NOR2X1
XFILL_33_3 gnd vdd FILL
XFILL_26_2 gnd vdd FILL
XFILL_33_4_0 gnd vdd FILL
XNOR2X1_469 NOR2X1_3/A INVX2_89/A gnd AND2X2_100/A vdd NOR2X1
XOAI21X1_909 AOI21X1_235/Y OAI21X1_908/Y NOR2X1_432/Y gnd OAI21X1_909/Y vdd OAI21X1
XINVX2_17 INVX2_17/A gnd INVX2_17/Y vdd INVX2
XINVX1_590 INVX1_517/A gnd INVX1_590/Y vdd INVX1
XNAND2X1_904 INVX1_632/Y BUFX4_96/Y gnd NAND2X1_904/Y vdd NAND2X1
XNAND2X1_915 DFFPOSX1_41/Q INVX2_76/Y gnd NAND2X1_915/Y vdd NAND2X1
XINVX2_39 INVX2_39/A gnd INVX2_39/Y vdd INVX2
XINVX2_28 INVX2_28/A gnd INVX2_28/Y vdd INVX2
XNAND2X1_937 INVX1_669/A INVX1_670/Y gnd AND2X2_82/B vdd NAND2X1
XNAND2X1_926 NOR2X1_411/Y OAI21X1_881/Y gnd NAND2X1_926/Y vdd NAND2X1
XNAND2X1_959 OR2X2_64/A OR2X2_64/B gnd NAND2X1_959/Y vdd NAND2X1
XNAND2X1_948 INVX1_679/Y INVX1_680/Y gnd NAND2X1_948/Y vdd NAND2X1
XFILL_24_4_0 gnd vdd FILL
XFILL_7_5_0 gnd vdd FILL
XFILL_15_4_0 gnd vdd FILL
XMUX2X1_1 MUX2X1_1/A MUX2X1_1/B INVX4_4/A gnd MUX2X1_1/Y vdd MUX2X1
XDFFPOSX1_108 INVX1_221/A CLKBUF1_15/Y OAI21X1_157/C gnd vdd DFFPOSX1
XDFFPOSX1_119 INVX2_88/A CLKBUF1_8/Y AND2X2_93/B gnd vdd DFFPOSX1
XCLKBUF1_2 BUFX4_6/Y gnd CLKBUF1_2/Y vdd CLKBUF1
XBUFX4_151 BUFX4_148/A gnd BUFX4_151/Y vdd BUFX4
XBUFX4_173 BUFX4_175/A gnd OR2X2_30/B vdd BUFX4
XNOR2X1_200 NOR2X1_200/A NOR2X1_200/B gnd NOR2X1_200/Y vdd NOR2X1
XBUFX4_140 OAI22X1_1/Y gnd AND2X2_2/A vdd BUFX4
XBUFX4_162 NOR2X1_2/Y gnd BUFX4_162/Y vdd BUFX4
XNOR2X1_211 INVX8_4/A MUX2X1_12/Y gnd AOI21X1_78/B vdd NOR2X1
XNOR2X1_222 INVX8_3/A NOR2X1_222/B gnd AND2X2_55/A vdd NOR2X1
XNOR2X1_233 AND2X2_35/B AND2X2_35/A gnd NOR2X1_233/Y vdd NOR2X1
XBUFX4_195 BUFX4_194/A gnd BUFX4_195/Y vdd BUFX4
XBUFX4_184 OR2X2_2/Y gnd BUFX4_184/Y vdd BUFX4
XNOR2X1_255 NOR2X1_255/A AND2X2_41/Y gnd NOR2X1_255/Y vdd NOR2X1
XNOR2X1_244 INVX2_46/Y MUX2X1_30/B gnd NOR2X1_244/Y vdd NOR2X1
XNOR2X1_266 INVX8_3/A AND2X2_29/Y gnd NOR2X1_267/A vdd NOR2X1
XNOR2X1_299 BUFX4_126/Y NOR2X1_299/B gnd NOR2X1_299/Y vdd NOR2X1
XNOR2X1_288 OR2X2_30/B NOR2X1_329/B gnd AOI22X1_98/C vdd NOR2X1
XNOR2X1_277 INVX8_7/A OR2X2_33/A gnd NOR2X1_277/Y vdd NOR2X1
XOAI21X1_706 OR2X2_24/A OR2X2_24/B NOR2X1_81/Y gnd OAI21X1_706/Y vdd OAI21X1
XOAI21X1_728 BUFX4_129/Y NOR2X1_256/B OAI21X1_728/C gnd AND2X2_68/B vdd OAI21X1
XOAI21X1_717 NOR2X1_344/Y NOR2X1_345/Y NOR3X1_56/Y gnd NAND3X1_163/A vdd OAI21X1
XOAI21X1_739 NOR2X1_76/Y INVX8_12/Y OAI21X1_739/C gnd NOR2X1_352/B vdd OAI21X1
XOAI21X1_1030 BUFX4_65/Y BUFX4_69/Y AOI22X1_149/Y gnd OAI21X1_1030/Y vdd OAI21X1
XOAI21X1_1052 BUFX4_254/Y OAI21X1_956/Y AOI22X1_168/Y gnd OAI21X1_1052/Y vdd OAI21X1
XOAI21X1_1041 BUFX4_66/Y BUFX4_71/Y AOI22X1_157/Y gnd OAI21X1_1041/Y vdd OAI21X1
XOAI21X1_1063 INVX2_93/Y INVX1_758/Y OAI21X1_1062/Y gnd OAI21X1_1064/A vdd OAI21X1
XNAND2X1_712 OAI21X1_66/Y BUFX4_131/Y gnd NAND2X1_712/Y vdd NAND2X1
XNAND2X1_701 XOR2X1_2/A INVX2_74/Y gnd NAND3X1_187/B vdd NAND2X1
XNAND2X1_745 OAI21X1_77/Y BUFX4_132/Y gnd NAND2X1_747/A vdd NAND2X1
XNAND2X1_723 NAND2X1_723/A NAND2X1_723/B gnd NAND2X1_5/B vdd NAND2X1
XNAND2X1_734 INVX1_519/Y BUFX4_205/Y gnd NAND3X1_207/C vdd NAND2X1
XNAND2X1_767 INVX1_541/Y BUFX4_203/Y gnd NAND3X1_229/C vdd NAND2X1
XNAND2X1_778 OAI21X1_88/Y BUFX4_134/Y gnd NAND2X1_780/A vdd NAND2X1
XNAND2X1_756 NAND2X1_754/Y NAND2X1_756/B gnd NAND2X1_16/B vdd NAND2X1
XNAND2X1_789 NAND2X1_787/Y NAND2X1_789/B gnd NAND2X1_27/B vdd NAND2X1
XFILL_40_7_1 gnd vdd FILL
XINVX8_4 INVX8_4/A gnd INVX8_4/Y vdd INVX8
XDFFPOSX1_90 INVX1_203/A CLKBUF1_50/Y OAI21X1_121/C gnd vdd DFFPOSX1
XBUFX4_13 BUFX4_13/A gnd BUFX4_13/Y vdd BUFX4
XBUFX4_24 BUFX4_22/A gnd BUFX4_24/Y vdd BUFX4
XBUFX4_35 BUFX4_37/A gnd BUFX4_35/Y vdd BUFX4
XBUFX4_57 INVX8_3/Y gnd BUFX4_57/Y vdd BUFX4
XBUFX4_46 BUFX4_46/A gnd NOR3X1_8/C vdd BUFX4
XBUFX4_68 BUFX4_69/A gnd BUFX4_68/Y vdd BUFX4
XBUFX4_79 INVX8_6/Y gnd BUFX4_79/Y vdd BUFX4
XNAND3X1_340 AND2X2_83/A AND2X2_83/B NOR3X1_70/Y gnd NOR2X1_462/B vdd NAND3X1
XFILL_31_7_1 gnd vdd FILL
XNAND3X1_351 INVX8_15/A NAND3X1_1/B INVX2_89/Y gnd NOR2X1_474/B vdd NAND3X1
XNAND3X1_362 NAND3X1_362/A NAND3X1_362/B OAI21X1_971/C gnd NAND3X1_362/Y vdd NAND3X1
XFILL_30_2_0 gnd vdd FILL
XOR2X2_49 OR2X2_49/A OR2X2_49/B gnd OR2X2_49/Y vdd OR2X2
XOR2X2_27 INVX4_6/A OR2X2_27/B gnd OR2X2_27/Y vdd OR2X2
XOR2X2_38 OR2X2_38/A OR2X2_38/B gnd OR2X2_38/Y vdd OR2X2
XOR2X2_16 OR2X2_16/A NOR2X1_1/A gnd OR2X2_16/Y vdd OR2X2
XOR2X2_9 OR2X2_9/A INVX2_5/Y gnd OR2X2_9/Y vdd OR2X2
XFILL_38_3_0 gnd vdd FILL
XINVX8_16 INVX8_16/A gnd INVX8_16/Y vdd INVX8
XFILL_22_7_1 gnd vdd FILL
XOAI21X1_514 OAI22X1_21/Y AOI21X1_69/Y AOI21X1_97/Y gnd AOI21X1_99/B vdd OAI21X1
XOAI21X1_503 AOI21X1_77/Y NAND3X1_91/Y AOI21X1_91/Y gnd AOI21X1_92/B vdd OAI21X1
XFILL_21_2_0 gnd vdd FILL
XOAI21X1_547 NAND2X1_498/Y NOR2X1_273/Y AOI21X1_109/Y gnd OAI21X1_547/Y vdd OAI21X1
XOAI21X1_525 NOR2X1_253/B INVX4_8/Y AND2X2_36/A gnd XNOR2X1_49/A vdd OAI21X1
XOAI21X1_536 NOR2X1_260/Y NOR2X1_259/Y BUFX4_124/Y gnd OAI21X1_536/Y vdd OAI21X1
XOAI21X1_569 INVX1_395/Y BUFX4_214/Y OAI21X1_569/C gnd NAND2X1_561/B vdd OAI21X1
XOAI21X1_558 INVX8_3/A OAI21X1_558/B OAI21X1_558/C gnd NOR2X1_278/B vdd OAI21X1
XDFFPOSX1_483 BUFX2_50/A CLKBUF1_7/Y NAND3X1_29/Y gnd vdd DFFPOSX1
XDFFPOSX1_450 NAND3X1_26/A CLKBUF1_7/Y BUFX2_49/A gnd vdd DFFPOSX1
XDFFPOSX1_461 NAND3X1_48/A CLKBUF1_52/Y BUFX2_60/A gnd vdd DFFPOSX1
XDFFPOSX1_472 BUFX2_39/A CLKBUF1_5/Y AOI21X1_1/Y gnd vdd DFFPOSX1
XNAND2X1_520 MUX2X1_40/S MUX2X1_37/Y gnd NAND2X1_520/Y vdd NAND2X1
XDFFPOSX1_494 BUFX2_61/A CLKBUF1_27/Y NAND3X1_51/Y gnd vdd DFFPOSX1
XNAND2X1_531 INVX1_329/A NAND2X1_530/Y gnd INVX1_399/A vdd NAND2X1
XNAND2X1_542 BUFX4_81/Y AND2X2_67/A gnd NOR2X1_314/B vdd NAND2X1
XNAND2X1_553 INVX8_7/A NOR2X1_217/Y gnd AOI21X1_160/B vdd NAND2X1
XNAND2X1_564 INVX8_5/A NAND2X1_564/B gnd NAND2X1_564/Y vdd NAND2X1
XNAND2X1_575 INVX2_62/Y AND2X2_39/Y gnd NAND2X1_575/Y vdd NAND2X1
XNAND2X1_586 INVX4_7/A INVX1_391/A gnd NAND2X1_586/Y vdd NAND2X1
XNAND2X1_597 INVX1_311/Y NOR2X1_362/B gnd AND2X2_69/A vdd NAND2X1
XFILL_4_3_0 gnd vdd FILL
XFILL_29_3_0 gnd vdd FILL
XFILL_13_7_1 gnd vdd FILL
XFILL_12_2_0 gnd vdd FILL
XNAND3X1_192 INVX1_506/Y BUFX4_210/Y BUFX4_37/Y gnd NAND3X1_192/Y vdd NAND3X1
XNAND3X1_181 OR2X2_45/A AND2X2_76/Y AND2X2_77/Y gnd NOR3X1_65/C vdd NAND3X1
XNAND3X1_170 INVX8_11/Y OAI21X1_753/Y NAND3X1_170/C gnd NAND3X1_171/A vdd NAND3X1
XOAI21X1_300 INVX1_327/Y INVX4_4/A OAI21X1_300/C gnd INVX2_53/A vdd OAI21X1
XOAI21X1_311 INVX1_334/Y INVX4_4/A NAND2X1_252/Y gnd MUX2X1_35/A vdd OAI21X1
XOAI21X1_322 INVX1_344/Y INVX4_4/A OAI21X1_322/C gnd MUX2X1_30/A vdd OAI21X1
XOAI21X1_344 BUFX4_39/Y MUX2X1_17/Y OAI21X1_452/C gnd OAI21X1_344/Y vdd OAI21X1
XOAI21X1_355 INVX2_24/Y BUFX4_40/Y NAND2X1_334/Y gnd MUX2X1_19/B vdd OAI21X1
XOAI21X1_333 NOR2X1_137/Y NOR2X1_138/Y INVX1_428/A gnd OAI21X1_333/Y vdd OAI21X1
XOAI21X1_399 NOR2X1_191/Y NOR2X1_192/Y INVX8_5/A gnd OAI21X1_399/Y vdd OAI21X1
XOAI21X1_366 BUFX4_213/Y MUX2X1_26/B NAND2X1_342/Y gnd OAI21X1_366/Y vdd OAI21X1
XINVX1_408 INVX1_408/A gnd INVX1_408/Y vdd INVX1
XOAI21X1_388 INVX2_30/Y BUFX4_44/Y NAND2X1_372/Y gnd NAND2X1_373/B vdd OAI21X1
XOAI21X1_377 AOI21X1_46/Y OAI21X1_341/Y AOI21X1_57/Y gnd INVX1_65/A vdd OAI21X1
XINVX1_419 INVX1_419/A gnd AND2X2_65/B vdd INVX1
XDFFPOSX1_280 AOI22X1_63/A CLKBUF1_36/Y NAND3X1_58/A gnd vdd DFFPOSX1
XDFFPOSX1_291 NOR2X1_6/A CLKBUF1_34/Y NOR3X1_14/Y gnd vdd DFFPOSX1
XXOR2X1_11 OR2X2_50/B INVX2_2/A gnd XOR2X1_11/Y vdd XOR2X1
XNAND2X1_361 BUFX4_127/Y NOR3X1_56/Y gnd INVX4_6/A vdd NAND2X1
XNAND2X1_372 BUFX4_44/Y MUX2X1_44/B gnd NAND2X1_372/Y vdd NAND2X1
XNAND2X1_350 AND2X2_25/Y INVX1_358/Y gnd NAND3X1_102/C vdd NAND2X1
XNAND2X1_383 BUFX4_41/Y MUX2X1_30/A gnd OAI21X1_469/C vdd NAND2X1
XNAND2X1_394 AOI22X1_87/A OAI21X1_391/Y gnd NAND2X1_394/Y vdd NAND2X1
XFILL_7_1 gnd vdd FILL
XFILL_36_6_1 gnd vdd FILL
XFILL_35_1_0 gnd vdd FILL
XNAND3X1_1 INVX1_715/A NAND3X1_1/B NOR2X1_4/Y gnd NAND3X1_1/Y vdd NAND3X1
XFILL_2_6_1 gnd vdd FILL
XFILL_27_6_1 gnd vdd FILL
XFILL_1_1_0 gnd vdd FILL
XFILL_26_1_0 gnd vdd FILL
XFILL_10_5_1 gnd vdd FILL
XOAI21X1_130 BUFX4_185/Y INVX1_115/Y OAI21X1_130/C gnd INVX1_609/A vdd OAI21X1
XOAI21X1_163 BUFX4_12/Y BUFX4_199/Y OAI21X1_163/C gnd NAND3X1_11/C vdd OAI21X1
XOAI21X1_174 BUFX4_15/Y BUFX4_200/Y OAI21X1_835/Y gnd NAND3X1_33/C vdd OAI21X1
XOAI21X1_141 BUFX4_273/Y BUFX4_193/Y OAI21X1_141/C gnd OAI21X1_141/Y vdd OAI21X1
XOAI21X1_152 BUFX4_184/Y INVX1_126/Y OAI21X1_152/C gnd INVX1_558/A vdd OAI21X1
XAOI22X1_6 INVX2_2/Y OR2X2_50/B INVX2_3/A AOI22X1_6/D gnd AOI22X1_6/Y vdd AOI22X1
XOAI21X1_185 BUFX4_16/Y BUFX4_198/Y OAI21X1_857/Y gnd NAND3X1_55/C vdd OAI21X1
XINVX1_216 INVX1_216/A gnd INVX1_216/Y vdd INVX1
XINVX1_205 INVX1_205/A gnd INVX1_205/Y vdd INVX1
XOAI21X1_196 BUFX4_142/Y INVX1_194/Y AOI22X1_11/Y gnd OAI21X1_196/Y vdd OAI21X1
XINVX1_249 INVX1_249/A gnd INVX1_249/Y vdd INVX1
XINVX1_238 INVX1_66/A gnd NOR3X1_48/A vdd INVX1
XINVX1_227 NOR2X1_18/A gnd INVX1_227/Y vdd INVX1
XFILL_9_2_0 gnd vdd FILL
XNAND2X1_16 BUFX4_19/Y NAND2X1_16/B gnd OAI21X1_16/C vdd NAND2X1
XNAND2X1_180 NAND2X1_180/A INVX2_15/Y gnd XOR2X1_6/B vdd NAND2X1
XNAND2X1_27 BUFX4_19/Y NAND2X1_27/B gnd OAI21X1_27/C vdd NAND2X1
XNAND2X1_38 BUFX4_29/Y NAND2X1_38/B gnd OAI21X1_38/C vdd NAND2X1
XNAND2X1_49 BUFX4_25/Y NAND2X1_49/B gnd OAI21X1_49/C vdd NAND2X1
XNAND2X1_191 INVX1_295/Y AOI21X1_35/B gnd NOR2X1_66/B vdd NAND2X1
XFILL_18_6_1 gnd vdd FILL
XFILL_17_1_0 gnd vdd FILL
XAOI21X1_209 AOI21X1_89/A OAI22X1_33/B AOI21X1_209/C gnd AOI21X1_209/Y vdd AOI21X1
XAOI22X1_14 AOI22X1_14/A BUFX4_237/Y BUFX4_259/Y AOI22X1_14/D gnd AOI22X1_14/Y vdd
+ AOI22X1
XAOI22X1_47 MUX2X1_10/A BUFX4_235/Y BUFX4_151/Y INVX1_681/A gnd AOI22X1_47/Y vdd AOI22X1
XAOI22X1_25 AOI22X1_25/A OR2X2_3/B BUFX4_257/Y AOI22X1_25/D gnd AOI22X1_25/Y vdd AOI22X1
XAOI22X1_36 AOI22X1_36/A AOI22X1_9/B OR2X2_3/A AOI22X1_36/D gnd AOI22X1_36/Y vdd AOI22X1
XAOI22X1_58 AOI22X1_58/A AND2X2_12/A BUFX4_146/Y INVX1_672/A gnd OR2X2_13/A vdd AOI22X1
XAOI22X1_69 AND2X2_59/A AND2X2_59/B AOI22X1_69/C INVX1_412/A gnd INVX1_328/A vdd AOI22X1
XNOR3X1_4 NOR3X1_4/A NOR3X1_4/B NOR3X1_4/C gnd NOR3X1_4/Y vdd NOR3X1
XINVX1_750 data_memory_interface_data[22] gnd INVX1_750/Y vdd INVX1
XBUFX2_90 BUFX2_90/A gnd BUFX2_90/Y vdd BUFX2
XOAI22X1_9 OAI22X1_9/A OAI22X1_9/B OAI22X1_9/C OAI22X1_9/D gnd OAI22X1_9/Y vdd OAI22X1
XFILL_42_4_1 gnd vdd FILL
XAOI21X1_80 AOI21X1_80/A AOI21X1_80/B AOI21X1_80/C gnd AOI21X1_80/Y vdd AOI21X1
XAOI21X1_91 AOI21X1_91/A NAND3X1_91/C AOI21X1_91/C gnd AOI21X1_91/Y vdd AOI21X1
XNOR2X1_404 NOR2X1_404/A NOR2X1_404/B gnd NOR2X1_404/Y vdd NOR2X1
XNOR2X1_415 INVX1_650/Y BUFX4_260/Y gnd NOR2X1_415/Y vdd NOR2X1
XNOR2X1_448 OR2X2_56/B INVX1_701/Y gnd NOR2X1_448/Y vdd NOR2X1
XNOR2X1_437 INVX1_443/A INVX1_689/Y gnd NOR2X1_437/Y vdd NOR2X1
XNOR2X1_426 MUX2X1_1/B INVX2_86/A gnd NOR2X1_426/Y vdd NOR2X1
XNOR2X1_459 NOR2X1_459/A NOR2X1_459/B gnd NOR2X1_459/Y vdd NOR2X1
XFILL_26_3 gnd vdd FILL
XFILL_33_4_1 gnd vdd FILL
XINVX2_18 INVX2_18/A gnd INVX2_18/Y vdd INVX2
XINVX1_580 INVX1_507/A gnd INVX1_580/Y vdd INVX1
XNAND2X1_916 DFFPOSX1_43/Q INVX2_77/Y gnd OAI21X1_875/C vdd NAND2X1
XINVX2_29 INVX2_29/A gnd INVX2_29/Y vdd INVX2
XNAND2X1_927 NAND2X1_927/A NAND2X1_927/B gnd NOR2X1_419/B vdd NAND2X1
XNAND2X1_905 NAND2X1_903/Y NAND2X1_905/B gnd NAND2X1_61/B vdd NAND2X1
XINVX1_591 INVX1_591/A gnd INVX1_591/Y vdd INVX1
XNAND2X1_938 INVX1_700/A INVX1_671/Y gnd NAND3X1_337/A vdd NAND2X1
XNAND2X1_949 OR2X2_57/A OR2X2_57/B gnd AOI22X1_129/A vdd NAND2X1
XFILL_24_4_1 gnd vdd FILL
XFILL_7_5_1 gnd vdd FILL
XFILL_6_0_0 gnd vdd FILL
XXOR2X1_1 XOR2X1_1/A INVX2_76/A gnd XOR2X1_1/Y vdd XOR2X1
XFILL_15_4_1 gnd vdd FILL
XMUX2X1_2 MUX2X1_2/A MUX2X1_2/B INVX4_4/A gnd MUX2X1_2/Y vdd MUX2X1
XDFFPOSX1_109 INVX1_222/A CLKBUF1_31/Y OAI21X1_159/C gnd vdd DFFPOSX1
XCLKBUF1_3 BUFX4_4/Y gnd CLKBUF1_3/Y vdd CLKBUF1
XBUFX4_130 INVX8_7/Y gnd AND2X2_56/B vdd BUFX4
XBUFX4_152 BUFX4_152/A gnd BUFX4_152/Y vdd BUFX4
XBUFX4_163 NOR2X1_2/Y gnd BUFX4_163/Y vdd BUFX4
XBUFX4_141 OR2X2_3/Y gnd BUFX4_141/Y vdd BUFX4
XNOR2X1_234 INVX8_3/A MUX2X1_38/B gnd INVX1_385/A vdd NOR2X1
XNOR2X1_212 MUX2X1_47/S MUX2X1_21/A gnd NOR2X1_212/Y vdd NOR2X1
XBUFX4_174 BUFX4_175/A gnd INVX8_9/A vdd BUFX4
XNOR2X1_201 NOR2X1_160/Y NOR2X1_201/B gnd NOR2X1_201/Y vdd NOR2X1
XBUFX4_196 INVX8_2/Y gnd BUFX4_196/Y vdd BUFX4
XNOR2X1_223 INVX8_4/A NOR2X1_223/B gnd NOR2X1_223/Y vdd NOR2X1
XBUFX4_185 OR2X2_2/Y gnd BUFX4_185/Y vdd BUFX4
XNOR2X1_245 INVX2_46/A MUX2X1_16/Y gnd OAI22X1_22/D vdd NOR2X1
XNOR2X1_267 NOR2X1_267/A NOR2X1_267/B gnd AOI22X1_95/B vdd NOR2X1
XNOR2X1_256 INVX8_7/A NOR2X1_256/B gnd NOR2X1_256/Y vdd NOR2X1
XFILL_31_1 gnd vdd FILL
XNOR2X1_278 INVX8_7/A NOR2X1_278/B gnd NOR2X1_278/Y vdd NOR2X1
XNOR2X1_289 INVX8_3/A MUX2X1_29/B gnd OAI22X1_33/B vdd NOR2X1
XOAI21X1_718 OR2X2_30/A OR2X2_33/B INVX8_7/A gnd NAND3X1_161/C vdd OAI21X1
XOAI21X1_707 OAI22X1_20/A INVX2_19/A OAI21X1_706/Y gnd OAI21X1_707/Y vdd OAI21X1
XOAI21X1_729 INVX2_18/Y OAI22X1_43/B NAND2X1_587/Y gnd NOR2X1_347/B vdd OAI21X1
XOAI21X1_1020 INVX1_742/Y INVX2_93/A OAI21X1_1019/Y gnd AOI22X1_146/C vdd OAI21X1
XOAI21X1_1031 INVX1_754/Y INVX2_93/Y NAND2X1_1020/Y gnd AOI22X1_150/C vdd OAI21X1
XOAI21X1_1053 BUFX4_252/Y OAI21X1_963/C AOI22X1_169/Y gnd OAI21X1_1053/Y vdd OAI21X1
XOAI21X1_1042 BUFX4_64/Y BUFX4_68/Y AOI22X1_158/Y gnd OAI21X1_1042/Y vdd OAI21X1
XOAI21X1_1064 OAI21X1_1064/A INVX1_757/Y NOR2X1_487/Y gnd OAI21X1_1064/Y vdd OAI21X1
XNAND2X1_702 OAI21X1_65/Y BUFX4_132/Y gnd NAND2X1_711/A vdd NAND2X1
XNAND2X1_713 INVX1_505/Y BUFX4_204/Y gnd NAND3X1_193/C vdd NAND2X1
XNAND2X1_724 OAI21X1_70/Y BUFX4_133/Y gnd NAND2X1_724/Y vdd NAND2X1
XNAND2X1_735 NAND2X1_733/Y NAND2X1_735/B gnd NAND2X1_9/B vdd NAND2X1
XNAND2X1_746 INVX1_527/Y BUFX4_202/Y gnd NAND3X1_215/C vdd NAND2X1
XNAND2X1_757 OAI21X1_81/Y BUFX4_134/Y gnd NAND2X1_759/A vdd NAND2X1
XNAND2X1_768 NAND2X1_768/A NAND2X1_768/B gnd NAND2X1_20/B vdd NAND2X1
XNAND2X1_779 INVX1_549/Y BUFX4_201/Y gnd NAND3X1_237/C vdd NAND2X1
XINVX8_5 INVX8_5/A gnd INVX8_5/Y vdd INVX8
XDFFPOSX1_80 INVX1_193/A CLKBUF1_11/Y OAI21X1_101/C gnd vdd DFFPOSX1
XDFFPOSX1_91 INVX1_204/A CLKBUF1_11/Y OAI21X1_123/C gnd vdd DFFPOSX1
XBUFX4_14 BUFX4_13/A gnd BUFX4_14/Y vdd BUFX4
XBUFX4_25 BUFX4_27/A gnd BUFX4_25/Y vdd BUFX4
XBUFX4_58 INVX8_3/Y gnd BUFX4_58/Y vdd BUFX4
XBUFX4_47 BUFX4_46/A gnd NOR3X1_9/C vdd BUFX4
XBUFX4_69 BUFX4_69/A gnd BUFX4_69/Y vdd BUFX4
XBUFX4_36 BUFX4_37/A gnd BUFX4_36/Y vdd BUFX4
XNAND3X1_341 NOR2X1_459/Y NAND3X1_341/B NOR3X1_72/Y gnd NOR2X1_465/B vdd NAND3X1
XNAND3X1_330 AND2X2_81/Y NOR2X1_422/Y AOI22X1_126/Y gnd NOR2X1_424/B vdd NAND3X1
XNAND3X1_352 NOR2X1_3/A NOR3X1_76/Y NOR2X1_474/Y gnd NAND3X1_352/Y vdd NAND3X1
XFILL_30_2_1 gnd vdd FILL
XOR2X2_39 OR2X2_39/A OR2X2_39/B gnd OR2X2_39/Y vdd OR2X2
XOR2X2_28 OR2X2_28/A INVX2_47/A gnd OR2X2_28/Y vdd OR2X2
XOR2X2_17 OR2X2_17/A OR2X2_17/B gnd OR2X2_17/Y vdd OR2X2
XFILL_38_3_1 gnd vdd FILL
XINVX8_17 INVX8_17/A gnd INVX8_17/Y vdd INVX8
XOAI21X1_504 INVX4_8/Y AOI21X1_92/B AOI21X1_92/Y gnd NAND3X1_122/A vdd OAI21X1
XFILL_21_2_1 gnd vdd FILL
XOAI21X1_526 INVX2_58/A OAI21X1_526/B BUFX4_92/Y gnd OAI21X1_526/Y vdd OAI21X1
XOAI21X1_515 NOR2X1_246/B AOI21X1_86/Y AOI21X1_98/Y gnd AOI21X1_99/C vdd OAI21X1
XOAI21X1_548 NOR2X1_152/A AOI21X1_88/Y AOI21X1_111/Y gnd OAI21X1_548/Y vdd OAI21X1
XOAI21X1_537 OAI21X1_537/A OR2X2_40/B NAND2X1_494/Y gnd AOI22X1_95/C vdd OAI21X1
XOAI21X1_559 NOR2X1_278/Y NOR2X1_279/Y INVX4_5/Y gnd NAND3X1_134/A vdd OAI21X1
XDFFPOSX1_440 NAND3X1_8/A CLKBUF1_5/Y BUFX2_39/A gnd vdd DFFPOSX1
XDFFPOSX1_451 NAND3X1_28/A CLKBUF1_7/Y BUFX2_50/A gnd vdd DFFPOSX1
XDFFPOSX1_462 NAND3X1_50/A CLKBUF1_27/Y BUFX2_61/A gnd vdd DFFPOSX1
XDFFPOSX1_473 BUFX2_40/A CLKBUF1_5/Y AOI21X1_2/Y gnd vdd DFFPOSX1
XNAND2X1_521 BUFX4_217/Y OAI21X1_621/A gnd NAND2X1_521/Y vdd NAND2X1
XDFFPOSX1_484 BUFX2_51/A CLKBUF1_41/Y NAND3X1_31/Y gnd vdd DFFPOSX1
XNAND2X1_510 INVX2_40/A MUX2X1_35/B gnd OAI21X1_564/C vdd NAND2X1
XDFFPOSX1_495 BUFX2_62/A CLKBUF1_27/Y NAND3X1_53/Y gnd vdd DFFPOSX1
XNAND2X1_532 BUFX4_217/Y MUX2X1_40/Y gnd OAI21X1_596/C vdd NAND2X1
XNAND2X1_543 INVX8_7/A NOR2X1_209/Y gnd NAND2X1_543/Y vdd NAND2X1
XNAND2X1_554 INVX1_408/Y BUFX4_155/Y gnd NAND2X1_554/Y vdd NAND2X1
XNAND2X1_576 INVX4_7/A AND2X2_38/Y gnd NAND3X1_158/A vdd NAND2X1
XNAND2X1_565 INVX1_412/Y BUFX4_155/Y gnd NAND2X1_565/Y vdd NAND2X1
XNAND2X1_587 NOR2X1_72/Y BUFX4_152/Y gnd NAND2X1_587/Y vdd NAND2X1
XFILL_4_3_1 gnd vdd FILL
XNAND2X1_598 BUFX4_55/Y OAI22X1_42/Y gnd NAND2X1_598/Y vdd NAND2X1
XFILL_29_3_1 gnd vdd FILL
XFILL_12_2_1 gnd vdd FILL
XNAND3X1_193 BUFX4_222/Y NAND3X1_192/Y NAND3X1_193/C gnd NAND2X1_714/B vdd NAND3X1
XNAND3X1_182 BUFX2_51/A NOR2X1_386/Y NOR2X1_382/Y gnd NOR2X1_387/B vdd NAND3X1
XNAND3X1_160 INVX4_10/Y AND2X2_51/Y NOR2X1_341/Y gnd NOR2X1_342/B vdd NAND3X1
XNAND3X1_171 NAND3X1_171/A OAI21X1_756/Y AOI21X1_206/Y gnd INVX1_95/A vdd NAND3X1
XOAI21X1_323 INVX1_345/Y INVX4_4/A NAND2X1_287/Y gnd NOR2X1_151/B vdd OAI21X1
XOAI21X1_301 INVX1_325/Y INVX4_4/A NAND2X1_233/Y gnd MUX2X1_42/A vdd OAI21X1
XOAI21X1_312 INVX1_335/Y INVX4_4/A NAND2X1_255/Y gnd NOR2X1_123/B vdd OAI21X1
XOAI21X1_345 INVX8_5/A OAI21X1_344/Y NAND2X1_326/Y gnd INVX1_375/A vdd OAI21X1
XOAI21X1_356 INVX2_25/Y BUFX4_40/Y NAND2X1_335/Y gnd MUX2X1_19/A vdd OAI21X1
XOAI21X1_334 INVX2_16/Y INVX2_17/A OAI21X1_334/C gnd AOI22X1_75/B vdd OAI21X1
XOAI21X1_367 INVX8_3/A OAI21X1_366/Y OAI21X1_367/C gnd AOI21X1_54/B vdd OAI21X1
XOAI21X1_389 INVX1_363/Y BUFX4_225/Y NAND2X1_373/Y gnd INVX1_364/A vdd OAI21X1
XOAI21X1_378 INVX4_2/Y INVX8_8/A OAI21X1_378/C gnd INVX1_361/A vdd OAI21X1
XINVX1_409 INVX1_409/A gnd INVX1_409/Y vdd INVX1
XXOR2X1_12 OR2X2_49/B XOR2X1_12/B gnd XOR2X1_12/Y vdd XOR2X1
XDFFPOSX1_270 AOI22X1_53/A CLKBUF1_45/Y NAND3X1_38/A gnd vdd DFFPOSX1
XDFFPOSX1_281 AOI22X1_64/A CLKBUF1_47/Y NAND3X1_60/A gnd vdd DFFPOSX1
XDFFPOSX1_292 OR2X2_1/B CLKBUF1_40/Y NOR3X1_15/Y gnd vdd DFFPOSX1
XNAND2X1_362 BUFX4_217/Y NOR2X1_187/Y gnd NOR2X1_188/B vdd NAND2X1
XNAND2X1_340 INVX8_8/A MUX2X1_42/A gnd OAI21X1_364/C vdd NAND2X1
XNAND2X1_351 INVX2_51/A AND2X2_24/Y gnd OR2X2_23/A vdd NAND2X1
XNAND2X1_384 INVX8_4/A MUX2X1_27/B gnd OAI21X1_398/C vdd NAND2X1
XNAND2X1_373 BUFX4_225/Y NAND2X1_373/B gnd NAND2X1_373/Y vdd NAND2X1
XNAND2X1_395 INVX8_5/A MUX2X1_19/B gnd OAI21X1_408/C vdd NAND2X1
XNOR3X1_80 NOR3X1_80/A INVX8_16/Y NOR3X1_80/C gnd NOR3X1_80/Y vdd NOR3X1
XOAI21X1_890 INVX1_661/Y OAI21X1_887/B INVX4_11/Y gnd OAI21X1_890/Y vdd OAI21X1
XFILL_7_2 gnd vdd FILL
XFILL_35_1_1 gnd vdd FILL
XNAND3X1_2 NAND3X1_2/A NAND3X1_2/B XNOR2X1_2/Y gnd OAI22X1_1/A vdd NAND3X1
XFILL_1_1_1 gnd vdd FILL
XFILL_26_1_1 gnd vdd FILL
XOAI21X1_131 BUFX4_270/Y OR2X2_2/B DFFPOSX1_95/D gnd OAI21X1_132/C vdd OAI21X1
XOAI21X1_120 BUFX4_186/Y INVX1_110/Y OAI21X1_120/C gnd INVX1_599/A vdd OAI21X1
XOAI21X1_164 BUFX4_12/Y BUFX4_199/Y OAI21X1_164/C gnd NAND3X1_13/C vdd OAI21X1
XOAI21X1_142 BUFX4_183/Y INVX1_121/Y OAI21X1_141/Y gnd INVX1_621/A vdd OAI21X1
XAOI22X1_7 AOI22X1_7/A AND2X2_3/Y AND2X2_4/Y NOR3X1_17/Y gnd BUFX4_13/A vdd AOI22X1
XOAI21X1_153 OR2X2_2/A BUFX4_194/Y OAI21X1_153/C gnd OAI21X1_154/C vdd OAI21X1
XOAI21X1_175 BUFX4_15/Y BUFX4_200/Y OAI21X1_836/Y gnd NAND3X1_35/C vdd OAI21X1
XOAI21X1_186 BUFX4_13/Y BUFX4_196/Y OAI21X1_858/Y gnd NAND3X1_57/C vdd OAI21X1
XINVX1_206 INVX1_206/A gnd INVX1_206/Y vdd INVX1
XOAI21X1_197 BUFX4_145/Y INVX1_195/Y AOI22X1_12/Y gnd OAI21X1_197/Y vdd OAI21X1
XINVX1_217 INVX1_217/A gnd INVX1_217/Y vdd INVX1
XINVX1_239 INVX1_239/A gnd INVX1_239/Y vdd INVX1
XINVX1_228 INVX1_228/A gnd INVX1_228/Y vdd INVX1
XFILL_9_2_1 gnd vdd FILL
XNAND2X1_170 NAND2X1_170/A OR2X2_13/Y gnd NOR2X1_45/B vdd NAND2X1
XNAND2X1_17 BUFX4_24/Y NAND2X1_17/B gnd OAI21X1_17/C vdd NAND2X1
XNAND2X1_28 BUFX4_22/Y NAND2X1_28/B gnd OAI21X1_28/C vdd NAND2X1
XNAND2X1_39 BUFX4_27/Y NAND2X1_39/B gnd OAI21X1_39/C vdd NAND2X1
XNAND2X1_192 NAND3X1_87/Y OAI21X1_280/Y gnd NAND2X1_192/Y vdd NAND2X1
XNAND2X1_181 INVX1_279/Y NOR2X1_53/B gnd NAND2X1_182/A vdd NAND2X1
XFILL_17_1_1 gnd vdd FILL
XAOI22X1_15 AOI22X1_15/A BUFX4_238/Y BUFX4_256/Y AOI22X1_15/D gnd AOI22X1_15/Y vdd
+ AOI22X1
XAOI22X1_48 MUX2X1_8/A BUFX4_235/Y BUFX4_151/Y OR2X2_59/A gnd NOR2X1_31/B vdd AOI22X1
XAOI22X1_26 AOI22X1_26/A OR2X2_3/B BUFX4_257/Y AOI22X1_26/D gnd AOI22X1_26/Y vdd AOI22X1
XAOI22X1_37 AOI22X1_37/A AOI22X1_9/B OR2X2_3/A AOI22X1_37/D gnd AOI22X1_37/Y vdd AOI22X1
XAOI22X1_59 AOI22X1_59/A AND2X2_12/A AND2X2_11/A INVX1_700/A gnd OR2X2_14/A vdd AOI22X1
XNOR3X1_5 NOR3X1_9/A NOR3X1_5/B NOR3X1_9/C gnd NOR3X1_5/Y vdd NOR3X1
XINVX1_751 data_memory_interface_data[13] gnd INVX1_751/Y vdd INVX1
XINVX1_740 data_memory_interface_data[2] gnd INVX1_740/Y vdd INVX1
XBUFX2_80 BUFX2_80/A gnd BUFX2_80/Y vdd BUFX2
XBUFX2_91 BUFX2_91/A gnd BUFX2_91/Y vdd BUFX2
XAOI21X1_70 INVX1_373/Y INVX8_11/Y OR2X2_24/Y gnd AOI21X1_70/Y vdd AOI21X1
XAOI21X1_92 INVX4_8/Y AOI21X1_92/B BUFX4_86/Y gnd AOI21X1_92/Y vdd AOI21X1
XAOI21X1_81 INVX2_47/Y AOI21X1_81/B BUFX4_275/Y gnd AOI21X1_81/Y vdd AOI21X1
XNOR2X1_416 INVX1_651/Y BUFX4_261/Y gnd NOR2X1_416/Y vdd NOR2X1
XNOR2X1_405 XOR2X1_14/Y XOR2X1_15/Y gnd AND2X2_80/B vdd NOR2X1
XNOR2X1_449 INVX1_457/A INVX1_672/Y gnd NOR2X1_449/Y vdd NOR2X1
XNOR2X1_438 INVX1_442/A INVX1_690/Y gnd NOR2X1_438/Y vdd NOR2X1
XNOR2X1_427 MUX2X1_2/B INVX1_454/A gnd INVX1_697/A vdd NOR2X1
XINVX1_581 INVX1_581/A gnd INVX1_581/Y vdd INVX1
XINVX1_570 XOR2X1_1/A gnd INVX1_570/Y vdd INVX1
XINVX2_19 INVX2_19/A gnd INVX2_19/Y vdd INVX2
XNAND2X1_928 INVX1_467/A INVX1_664/Y gnd AOI21X1_245/A vdd NAND2X1
XNAND2X1_917 INVX2_79/A INVX1_642/Y gnd OAI22X1_49/A vdd NAND2X1
XNAND2X1_906 OAI21X1_94/Y BUFX4_59/Y gnd NAND2X1_906/Y vdd NAND2X1
XINVX1_592 INVX1_592/A gnd INVX1_592/Y vdd INVX1
XNAND2X1_939 INVX1_459/A INVX2_82/Y gnd NAND2X1_939/Y vdd NAND2X1
XFILL_6_0_1 gnd vdd FILL
XXOR2X1_2 XOR2X1_2/A INVX2_74/A gnd XOR2X1_2/Y vdd XOR2X1
XFILL_43_7_0 gnd vdd FILL
XMUX2X1_3 MUX2X1_3/A MUX2X1_3/B INVX4_4/A gnd MUX2X1_3/Y vdd MUX2X1
XCLKBUF1_4 BUFX4_6/Y gnd CLKBUF1_4/Y vdd CLKBUF1
XBUFX4_120 BUFX4_122/A gnd BUFX4_120/Y vdd BUFX4
XBUFX4_153 BUFX4_152/A gnd BUFX4_153/Y vdd BUFX4
XBUFX4_131 AND2X2_79/Y gnd BUFX4_131/Y vdd BUFX4
XBUFX4_142 OR2X2_3/Y gnd BUFX4_142/Y vdd BUFX4
XBUFX4_164 BUFX4_164/A gnd BUFX4_164/Y vdd BUFX4
XBUFX4_197 INVX8_2/Y gnd BUFX4_197/Y vdd BUFX4
XNOR2X1_224 INVX8_6/A MUX2X1_17/Y gnd AOI21X1_88/C vdd NOR2X1
XNOR2X1_213 INVX8_5/A MUX2X1_14/Y gnd AOI21X1_63/C vdd NOR2X1
XNOR2X1_202 BUFX4_129/Y NOR2X1_203/B gnd INVX2_54/A vdd NOR2X1
XBUFX4_175 BUFX4_175/A gnd OR2X2_33/B vdd BUFX4
XBUFX4_186 OR2X2_2/Y gnd BUFX4_186/Y vdd BUFX4
XNOR2X1_246 NOR2X1_246/A NOR2X1_246/B gnd NOR2X1_246/Y vdd NOR2X1
XNOR2X1_235 INVX8_5/A NOR2X1_235/B gnd INVX1_381/A vdd NOR2X1
XNOR2X1_257 INVX1_356/A INVX1_390/Y gnd NOR2X1_257/Y vdd NOR2X1
XFILL_31_2 gnd vdd FILL
XFILL_34_7_0 gnd vdd FILL
XNOR2X1_268 INVX2_43/A MUX2X1_8/Y gnd NOR2X1_269/A vdd NOR2X1
XNOR2X1_279 BUFX4_127/Y OR2X2_42/B gnd NOR2X1_279/Y vdd NOR2X1
XFILL_24_1 gnd vdd FILL
XOAI21X1_708 NOR2X1_342/B INVX1_405/A OAI21X1_708/C gnd OAI21X1_708/Y vdd OAI21X1
XOAI21X1_719 OAI21X1_719/A INVX4_9/Y OAI21X1_719/C gnd OAI21X1_719/Y vdd OAI21X1
XOAI21X1_1021 BUFX4_65/Y BUFX4_69/Y AOI22X1_146/Y gnd OAI21X1_1021/Y vdd OAI21X1
XOAI21X1_1010 INVX2_91/Y OAI21X1_981/B NAND2X1_1018/Y gnd AOI22X1_144/C vdd OAI21X1
XOAI21X1_1054 BUFX4_252/Y OAI21X1_965/C AOI22X1_170/Y gnd OAI21X1_1054/Y vdd OAI21X1
XOAI21X1_1043 BUFX4_64/Y BUFX4_68/Y AOI22X1_159/Y gnd OAI21X1_1043/Y vdd OAI21X1
XOAI21X1_1032 BUFX4_64/Y BUFX4_68/Y AOI22X1_150/Y gnd OAI21X1_1032/Y vdd OAI21X1
XOAI21X1_1065 INVX4_13/Y INVX8_16/Y AND2X2_101/B gnd OAI21X1_1066/C vdd OAI21X1
XNAND2X1_703 AND2X2_79/B AND2X2_79/A gnd BUFX4_222/A vdd NAND2X1
XNAND2X1_736 OAI21X1_74/Y BUFX4_131/Y gnd NAND2X1_738/A vdd NAND2X1
XNAND2X1_714 NAND2X1_712/Y NAND2X1_714/B gnd NAND2X1_2/B vdd NAND2X1
XNAND2X1_725 INVX1_513/Y BUFX4_203/Y gnd NAND3X1_201/C vdd NAND2X1
XNAND2X1_747 NAND2X1_747/A NAND2X1_747/B gnd NAND2X1_13/B vdd NAND2X1
XNAND2X1_769 OAI21X1_85/Y BUFX4_133/Y gnd NAND2X1_769/Y vdd NAND2X1
XNAND2X1_758 INVX1_535/Y BUFX4_203/Y gnd NAND3X1_223/C vdd NAND2X1
XFILL_0_7_0 gnd vdd FILL
XFILL_25_7_0 gnd vdd FILL
XINVX8_6 INVX8_6/A gnd INVX8_6/Y vdd INVX8
XDFFPOSX1_70 AOI22X1_32/A CLKBUF1_11/Y INVX1_123/A gnd vdd DFFPOSX1
XDFFPOSX1_81 INVX1_194/A CLKBUF1_3/Y DFFPOSX1_81/D gnd vdd DFFPOSX1
XDFFPOSX1_92 INVX1_205/A CLKBUF1_11/Y DFFPOSX1_92/D gnd vdd DFFPOSX1
XBUFX4_15 BUFX4_13/A gnd BUFX4_15/Y vdd BUFX4
XBUFX4_26 BUFX4_27/A gnd BUFX4_26/Y vdd BUFX4
XBUFX4_59 BUFX4_62/A gnd BUFX4_59/Y vdd BUFX4
XBUFX4_48 BUFX4_46/A gnd BUFX4_48/Y vdd BUFX4
XBUFX4_37 BUFX4_37/A gnd BUFX4_37/Y vdd BUFX4
XFILL_16_7_0 gnd vdd FILL
XNAND3X1_342 AND2X2_93/A NOR2X1_465/Y NOR2X1_462/Y gnd NAND2X1_993/A vdd NAND3X1
XNAND3X1_331 AOI22X1_127/Y NAND3X1_331/B AND2X2_82/Y gnd NOR2X1_424/A vdd NAND3X1
XNAND3X1_320 INVX1_637/Y BUFX4_100/Y BUFX4_165/Y gnd NAND3X1_321/B vdd NAND3X1
XNAND3X1_353 AND2X2_100/Y BUFX4_11/Y NOR3X1_76/Y gnd AOI21X1_259/A vdd NAND3X1
XOR2X2_18 INVX4_4/A OR2X2_62/A gnd OR2X2_18/Y vdd OR2X2
XOR2X2_29 OR2X2_29/A OR2X2_29/B gnd OR2X2_29/Y vdd OR2X2
XOAI21X1_505 BUFX4_227/Y INVX1_386/Y OAI21X1_505/C gnd NAND2X1_472/B vdd OAI21X1
XOAI21X1_527 NOR2X1_249/Y AND2X2_36/A AOI22X1_72/A gnd NOR2X1_254/A vdd OAI21X1
XOAI21X1_516 NOR2X1_238/Y NOR2X1_239/Y BUFX4_81/Y gnd OR2X2_29/A vdd OAI21X1
XOAI21X1_538 AND2X2_44/Y BUFX4_58/Y BUFX4_124/Y gnd NOR2X1_267/B vdd OAI21X1
XOAI21X1_549 NOR2X1_124/Y OAI21X1_526/B NAND2X1_297/Y gnd AOI21X1_113/B vdd OAI21X1
XDFFPOSX1_430 OR2X2_52/B CLKBUF1_39/Y NOR3X1_37/Y gnd vdd DFFPOSX1
XDFFPOSX1_474 BUFX2_41/A CLKBUF1_45/Y NAND3X1_11/Y gnd vdd DFFPOSX1
XDFFPOSX1_452 NAND3X1_30/A CLKBUF1_41/Y BUFX2_51/A gnd vdd DFFPOSX1
XDFFPOSX1_463 NAND3X1_52/A CLKBUF1_27/Y BUFX2_62/A gnd vdd DFFPOSX1
XDFFPOSX1_441 NAND3X1_9/A CLKBUF1_5/Y BUFX2_40/A gnd vdd DFFPOSX1
XNAND2X1_500 NAND2X1_500/A NAND2X1_500/B gnd AOI22X1_97/D vdd NAND2X1
XDFFPOSX1_485 BUFX2_52/A CLKBUF1_41/Y NAND3X1_33/Y gnd vdd DFFPOSX1
XDFFPOSX1_496 BUFX2_63/A CLKBUF1_36/Y NAND3X1_55/Y gnd vdd DFFPOSX1
XNAND2X1_511 BUFX4_55/Y NOR2X1_223/Y gnd NOR2X1_369/A vdd NAND2X1
XNAND2X1_533 INVX8_7/A NOR2X1_182/Y gnd NAND2X1_533/Y vdd NAND2X1
XNAND2X1_544 INVX1_402/Y BUFX4_154/Y gnd NAND2X1_544/Y vdd NAND2X1
XNAND2X1_522 INVX8_3/A AOI22X1_98/A gnd OAI21X1_577/C vdd NAND2X1
XNAND2X1_577 AND2X2_52/B AND2X2_52/A gnd NOR2X1_342/A vdd NAND2X1
XNAND2X1_555 INVX2_32/Y MUX2X1_44/A gnd INVX1_409/A vdd NAND2X1
XNAND2X1_566 MUX2X1_20/S MUX2X1_47/Y gnd OAI21X1_685/C vdd NAND2X1
XNAND2X1_588 INVX2_18/A OAI21X1_722/Y gnd OAI21X1_734/C vdd NAND2X1
XNAND2X1_599 NOR2X1_87/Y BUFX4_152/Y gnd OAI21X1_760/C vdd NAND2X1
XFILL_40_5_0 gnd vdd FILL
XAOI21X1_190 NAND2X1_578/Y AOI21X1_190/B NAND3X1_163/Y gnd AOI21X1_190/Y vdd AOI21X1
XNAND3X1_150 OAI21X1_655/Y NAND2X1_554/Y NAND3X1_150/C gnd NAND3X1_150/Y vdd NAND3X1
XFILL_31_5_0 gnd vdd FILL
XNAND3X1_183 NOR2X1_386/Y NOR2X1_389/Y NOR2X1_382/Y gnd NOR3X1_66/C vdd NAND3X1
XNAND3X1_161 INVX2_65/A OAI21X1_719/Y NAND3X1_161/C gnd NAND3X1_161/Y vdd NAND3X1
XNAND3X1_172 BUFX4_93/Y NAND2X1_602/Y OR2X2_43/Y gnd NAND3X1_172/Y vdd NAND3X1
XNAND3X1_194 INVX1_508/Y BUFX4_207/Y BUFX4_35/Y gnd NAND3X1_194/Y vdd NAND3X1
XFILL_39_6_0 gnd vdd FILL
XFILL_22_5_0 gnd vdd FILL
XOAI21X1_313 INVX1_336/Y INVX4_4/A NAND2X1_258/Y gnd NOR2X1_249/B vdd OAI21X1
XOAI21X1_302 NOR2X1_97/Y NOR2X1_98/Y INVX1_326/Y gnd OAI21X1_302/Y vdd OAI21X1
XOAI21X1_346 AOI21X1_50/Y OAI21X1_346/B NAND2X1_327/Y gnd OAI21X1_354/B vdd OAI21X1
XOAI21X1_324 AND2X2_35/B AOI22X1_89/C AOI22X1_89/B gnd AOI21X1_41/C vdd OAI21X1
XOAI21X1_335 AND2X2_64/B NAND2X1_319/Y NAND2X1_318/Y gnd AOI22X1_75/D vdd OAI21X1
XOAI21X1_368 BUFX4_82/Y INVX8_7/A BUFX4_78/Y gnd OR2X2_36/B vdd OAI21X1
XOAI21X1_357 NOR2X1_158/Y NOR2X1_159/Y BUFX4_225/Y gnd OAI21X1_357/Y vdd OAI21X1
XOAI21X1_379 INVX4_3/Y INVX8_8/A NAND2X1_365/Y gnd OAI21X1_379/Y vdd OAI21X1
XDFFPOSX1_260 INVX1_247/A CLKBUF1_54/Y NAND3X1_18/A gnd vdd DFFPOSX1
XDFFPOSX1_271 AOI22X1_54/A CLKBUF1_10/Y NAND3X1_40/A gnd vdd DFFPOSX1
XDFFPOSX1_282 AOI22X1_65/A CLKBUF1_17/Y NAND3X1_62/A gnd vdd DFFPOSX1
XXOR2X1_13 OR2X2_50/B XOR2X1_13/B gnd XOR2X1_13/Y vdd XOR2X1
XDFFPOSX1_293 INVX2_51/A CLKBUF1_25/Y NOR3X1_9/Y gnd vdd DFFPOSX1
XNAND2X1_341 BUFX4_227/Y INVX1_354/Y gnd NAND2X1_341/Y vdd NAND2X1
XNAND2X1_330 BUFX4_42/Y MUX2X1_35/B gnd OAI21X1_348/C vdd NAND2X1
XNAND2X1_363 NOR2X1_188/Y INVX4_6/Y gnd NAND2X1_363/Y vdd NAND2X1
XNAND2X1_352 NOR2X1_179/Y AND2X2_42/A gnd BUFX4_88/A vdd NAND2X1
XNAND2X1_374 INVX8_4/A INVX1_364/Y gnd NAND2X1_374/Y vdd NAND2X1
XFILL_5_6_0 gnd vdd FILL
XNAND2X1_385 BUFX4_42/Y NOR2X1_249/B gnd NAND2X1_385/Y vdd NAND2X1
XNAND2X1_396 INVX8_4/A MUX2X1_28/B gnd OAI21X1_412/C vdd NAND2X1
XNOR3X1_70 NOR3X1_70/A NOR3X1_70/B NOR3X1_70/C gnd NOR3X1_70/Y vdd NOR3X1
XNOR3X1_81 NOR3X1_79/Y data_memory_interface_data[31] NOR3X1_80/Y gnd NOR3X1_81/Y
+ vdd NOR3X1
XFILL_13_5_0 gnd vdd FILL
XOAI21X1_891 INVX8_14/Y AOI21X1_231/Y OAI21X1_891/C gnd OAI21X1_891/Y vdd OAI21X1
XOAI21X1_880 OAI21X1_877/A INVX1_647/Y OAI21X1_880/C gnd OAI21X1_880/Y vdd OAI21X1
XFILL_7_3 gnd vdd FILL
XNAND3X1_3 AOI22X1_5/Y AOI22X1_6/Y NAND3X1_3/C gnd OAI22X1_1/D vdd NAND3X1
XOAI21X1_121 BUFX4_272/Y BUFX4_195/Y OAI21X1_121/C gnd OAI21X1_121/Y vdd OAI21X1
XOAI21X1_110 BUFX4_184/Y INVX1_105/Y OAI21X1_109/Y gnd INVX1_589/A vdd OAI21X1
XOAI21X1_165 BUFX4_15/Y BUFX4_200/Y OAI21X1_819/Y gnd NAND3X1_15/C vdd OAI21X1
XAOI22X1_8 AOI22X1_8/A BUFX4_236/Y BUFX4_258/Y AOI22X1_8/D gnd AOI22X1_8/Y vdd AOI22X1
XOAI21X1_143 BUFX4_273/Y BUFX4_193/Y OAI21X1_143/C gnd OAI21X1_144/C vdd OAI21X1
XOAI21X1_132 BUFX4_185/Y INVX1_116/Y OAI21X1_132/C gnd INVX1_611/A vdd OAI21X1
XOAI21X1_154 BUFX4_186/Y INVX1_127/Y OAI21X1_154/C gnd INVX1_560/A vdd OAI21X1
XOAI21X1_198 OR2X2_4/A INVX1_196/Y AOI22X1_13/Y gnd OAI21X1_198/Y vdd OAI21X1
XOAI21X1_176 BUFX4_15/Y BUFX4_200/Y OAI21X1_838/Y gnd NAND3X1_37/C vdd OAI21X1
XOAI21X1_187 BUFX4_13/Y BUFX4_196/Y OAI21X1_859/Y gnd NAND3X1_59/C vdd OAI21X1
XINVX1_207 INVX1_207/A gnd INVX1_207/Y vdd INVX1
XINVX1_229 INVX1_229/A gnd OAI22X1_6/B vdd INVX1
XINVX1_218 INVX1_218/A gnd INVX1_218/Y vdd INVX1
XNAND2X1_160 OR2X2_10/B OR2X2_10/A gnd AOI21X1_27/A vdd NAND2X1
XNAND2X1_171 OR2X2_14/B OR2X2_14/A gnd NAND2X1_172/A vdd NAND2X1
XNAND2X1_18 BUFX4_18/Y NAND2X1_18/B gnd OAI21X1_18/C vdd NAND2X1
XNAND2X1_29 BUFX4_22/Y NAND2X1_29/B gnd OAI21X1_29/C vdd NAND2X1
XNAND2X1_193 AOI21X1_5/A AOI21X1_5/B gnd NOR2X1_68/B vdd NAND2X1
XNAND2X1_182 NAND2X1_182/A INVX1_280/Y gnd NOR2X1_54/B vdd NAND2X1
XAOI22X1_16 AOI22X1_16/A BUFX4_236/Y BUFX4_258/Y AOI22X1_16/D gnd AOI22X1_16/Y vdd
+ AOI22X1
XAOI22X1_38 AOI22X1_38/A BUFX4_236/Y BUFX4_258/Y AOI22X1_38/D gnd AOI22X1_38/Y vdd
+ AOI22X1
XAOI22X1_27 AOI22X1_27/A BUFX4_237/Y BUFX4_259/Y AOI22X1_27/D gnd AOI22X1_27/Y vdd
+ AOI22X1
XAOI22X1_49 MUX2X1_7/A BUFX4_235/Y BUFX4_151/Y MUX2X1_7/B gnd NOR2X1_32/B vdd AOI22X1
XNOR3X1_6 NOR3X1_9/A NOR3X1_6/B NOR3X1_9/C gnd NOR3X1_6/Y vdd NOR3X1
XINVX1_730 INVX1_730/A gnd INVX1_730/Y vdd INVX1
XINVX1_752 data_memory_interface_data[6] gnd INVX1_752/Y vdd INVX1
XINVX1_741 data_memory_interface_data[19] gnd INVX1_741/Y vdd INVX1
XFILL_36_4_0 gnd vdd FILL
XBUFX2_81 BUFX2_81/A gnd BUFX2_81/Y vdd BUFX2
XBUFX2_70 BUFX2_70/A gnd instruction_memory_interface_address[31] vdd BUFX2
XBUFX2_92 BUFX2_92/A gnd BUFX2_92/Y vdd BUFX2
XFILL_2_4_0 gnd vdd FILL
XFILL_27_4_0 gnd vdd FILL
XFILL_10_3_0 gnd vdd FILL
XAOI21X1_71 AOI21X1_71/A AOI21X1_70/Y AOI22X1_80/A gnd AOI21X1_71/Y vdd AOI21X1
XAOI21X1_60 INVX1_369/A AOI21X1_56/A INVX8_11/A gnd AOI21X1_60/Y vdd AOI21X1
XAOI21X1_82 AOI21X1_86/A BUFX4_189/Y AOI21X1_82/C gnd AOI21X1_82/Y vdd AOI21X1
XAOI21X1_93 BUFX4_41/Y NOR2X1_125/B AOI21X1_93/C gnd AOI21X1_93/Y vdd AOI21X1
XFILL_18_4_0 gnd vdd FILL
XNOR2X1_406 NOR2X1_406/A NOR2X1_406/B gnd AND2X2_80/A vdd NOR2X1
XNOR2X1_428 INVX1_451/A INVX1_675/Y gnd NOR2X1_428/Y vdd NOR2X1
XNOR2X1_417 INVX1_652/Y BUFX4_260/Y gnd NOR2X1_417/Y vdd NOR2X1
XNOR2X1_439 OR2X2_59/B INVX1_693/Y gnd NOR2X1_439/Y vdd NOR2X1
XINVX1_571 XOR2X1_2/A gnd INVX1_571/Y vdd INVX1
XINVX1_560 INVX1_560/A gnd INVX1_560/Y vdd INVX1
XNAND2X1_907 INVX1_634/Y BUFX4_98/Y gnd NAND3X1_319/C vdd NAND2X1
XNAND2X1_918 OAI22X1_6/Y INVX2_79/Y gnd OAI21X1_887/B vdd NAND2X1
XINVX1_593 INVX1_593/A gnd INVX1_593/Y vdd INVX1
XINVX1_582 INVX1_509/A gnd INVX1_582/Y vdd INVX1
XNAND2X1_929 INVX1_667/A INVX1_666/Y gnd AND2X2_81/A vdd NAND2X1
XXOR2X1_3 XOR2X1_3/A XOR2X1_3/B gnd XOR2X1_3/Y vdd XOR2X1
XFILL_43_7_1 gnd vdd FILL
XFILL_42_2_0 gnd vdd FILL
XMUX2X1_4 MUX2X1_4/A MUX2X1_4/B INVX4_4/A gnd MUX2X1_4/Y vdd MUX2X1
XCLKBUF1_5 BUFX4_5/Y gnd CLKBUF1_5/Y vdd CLKBUF1
XBUFX4_110 NOR2X1_7/Y gnd BUFX4_110/Y vdd BUFX4
XAOI22X1_170 BUFX4_254/Y INVX1_732/A AOI22X1_170/C BUFX4_106/Y gnd AOI22X1_170/Y vdd
+ AOI22X1
XBUFX4_121 BUFX4_122/A gnd BUFX4_121/Y vdd BUFX4
XBUFX4_154 BUFX4_152/A gnd BUFX4_154/Y vdd BUFX4
XBUFX4_132 AND2X2_79/Y gnd BUFX4_132/Y vdd BUFX4
XBUFX4_143 OR2X2_3/Y gnd OR2X2_4/A vdd BUFX4
XNOR2X1_214 NOR2X1_214/A BUFX4_87/Y gnd AOI21X1_72/C vdd NOR2X1
XNOR2X1_225 INVX8_3/A NOR2X1_225/B gnd NOR2X1_225/Y vdd NOR2X1
XBUFX4_176 BUFX4_175/A gnd BUFX4_176/Y vdd BUFX4
XNOR2X1_203 INVX8_7/A NOR2X1_203/B gnd INVX1_371/A vdd NOR2X1
XBUFX4_187 BUFX4_188/A gnd BUFX4_187/Y vdd BUFX4
XBUFX4_165 BUFX4_164/A gnd BUFX4_165/Y vdd BUFX4
XNOR2X1_247 OR2X2_30/A INVX4_6/A gnd NOR2X1_247/Y vdd NOR2X1
XBUFX4_198 INVX8_2/Y gnd BUFX4_198/Y vdd BUFX4
XNOR2X1_258 OR2X2_22/B OR2X2_31/B gnd AND2X2_42/B vdd NOR2X1
XNOR2X1_236 INVX8_4/A INVX1_381/Y gnd NOR2X1_236/Y vdd NOR2X1
XFILL_34_7_1 gnd vdd FILL
XNOR2X1_269 NOR2X1_269/A AND2X2_41/Y gnd NOR2X1_269/Y vdd NOR2X1
XFILL_24_2 gnd vdd FILL
XFILL_33_2_0 gnd vdd FILL
XOAI21X1_709 OAI21X1_743/A NOR2X1_80/Y INVX2_19/A gnd AND2X2_64/A vdd OAI21X1
XOAI21X1_1000 INVX1_747/Y OAI21X1_992/B OAI21X1_999/Y gnd AOI21X1_263/B vdd OAI21X1
XOAI21X1_1022 NOR2X1_481/Y INVX4_12/A data_memory_interface_data[27] gnd OAI21X1_1022/Y
+ vdd OAI21X1
XOAI21X1_1011 AOI21X1_265/Y OAI21X1_994/B AOI22X1_144/Y gnd OAI21X1_1011/Y vdd OAI21X1
XOAI21X1_1055 BUFX4_252/Y OAI21X1_967/C AOI22X1_171/Y gnd OAI21X1_1055/Y vdd OAI21X1
XOAI21X1_1044 BUFX4_67/Y BUFX4_70/Y AOI22X1_160/Y gnd OAI21X1_1044/Y vdd OAI21X1
XOAI21X1_1033 NOR2X1_481/Y INVX4_12/A data_memory_interface_data[31] gnd OAI21X1_1034/C
+ vdd OAI21X1
XOAI21X1_1066 INVX8_17/A BUFX4_253/Y OAI21X1_1066/C gnd OAI21X1_1066/Y vdd OAI21X1
XNAND2X1_704 OR2X2_49/A OR2X2_49/B gnd NAND2X1_704/Y vdd NAND2X1
XINVX1_390 INVX1_390/A gnd INVX1_390/Y vdd INVX1
XNAND2X1_715 OAI21X1_67/Y BUFX4_134/Y gnd NAND2X1_717/A vdd NAND2X1
XNAND2X1_726 NAND2X1_724/Y NAND2X1_726/B gnd NAND2X1_6/B vdd NAND2X1
XNAND2X1_737 INVX1_521/Y BUFX4_202/Y gnd NAND3X1_209/C vdd NAND2X1
XNAND2X1_759 NAND2X1_759/A NAND2X1_759/B gnd NAND2X1_17/B vdd NAND2X1
XNAND2X1_748 OAI21X1_78/Y BUFX4_132/Y gnd NAND2X1_750/A vdd NAND2X1
XFILL_0_7_1 gnd vdd FILL
XFILL_25_7_1 gnd vdd FILL
XFILL_24_2_0 gnd vdd FILL
XINVX8_7 INVX8_7/A gnd INVX8_7/Y vdd INVX8
XDFFPOSX1_71 AOI22X1_33/A CLKBUF1_24/Y INVX1_124/A gnd vdd DFFPOSX1
XDFFPOSX1_60 AOI22X1_22/A CLKBUF1_30/Y INVX1_113/A gnd vdd DFFPOSX1
XDFFPOSX1_93 INVX1_206/A CLKBUF1_15/Y OAI21X1_127/C gnd vdd DFFPOSX1
XDFFPOSX1_82 INVX1_195/A CLKBUF1_11/Y OAI21X1_105/C gnd vdd DFFPOSX1
XFILL_7_3_0 gnd vdd FILL
XBUFX4_16 BUFX4_13/A gnd BUFX4_16/Y vdd BUFX4
XBUFX4_38 INVX8_8/Y gnd BUFX4_38/Y vdd BUFX4
XBUFX4_49 BUFX4_46/A gnd BUFX4_49/Y vdd BUFX4
XBUFX4_27 BUFX4_27/A gnd BUFX4_27/Y vdd BUFX4
XFILL_16_7_1 gnd vdd FILL
XFILL_15_2_0 gnd vdd FILL
XNAND3X1_332 AND2X2_83/Y NOR3X1_70/Y NOR2X1_424/Y gnd OAI21X1_938/A vdd NAND3X1
XNAND3X1_310 INVX1_627/Y BUFX4_102/Y BUFX4_168/Y gnd NAND3X1_311/B vdd NAND3X1
XNAND3X1_321 BUFX4_121/Y NAND3X1_321/B NAND3X1_321/C gnd NAND2X1_911/B vdd NAND3X1
XNAND3X1_354 INVX1_717/Y NOR3X1_76/Y NOR2X1_474/Y gnd NAND3X1_354/Y vdd NAND3X1
XNAND3X1_343 OR2X2_67/Y AOI22X1_136/Y NAND3X1_343/C gnd NAND3X1_343/Y vdd NAND3X1
XOR2X2_19 OR2X2_19/A INVX8_5/A gnd OR2X2_19/Y vdd OR2X2
XOAI21X1_506 BUFX4_213/Y OAI21X1_506/B NAND2X1_472/Y gnd NOR2X1_238/B vdd OAI21X1
XOAI21X1_528 INVX2_59/Y NOR2X1_254/Y AOI21X1_103/Y gnd OAI21X1_528/Y vdd OAI21X1
XOAI21X1_539 NOR2X1_254/B NOR2X1_254/A INVX2_59/A gnd INVX1_392/A vdd OAI21X1
XOAI21X1_517 BUFX4_42/Y MUX2X1_10/Y NAND2X1_385/Y gnd NAND2X1_496/B vdd OAI21X1
XDFFPOSX1_420 BUFX2_84/A CLKBUF1_47/Y NOR3X1_27/Y gnd vdd DFFPOSX1
XDFFPOSX1_431 BUFX2_90/A CLKBUF1_59/Y NOR3X1_38/Y gnd vdd DFFPOSX1
XDFFPOSX1_442 NAND3X1_10/A CLKBUF1_52/Y BUFX2_41/A gnd vdd DFFPOSX1
XDFFPOSX1_453 NAND3X1_32/A CLKBUF1_41/Y BUFX2_52/A gnd vdd DFFPOSX1
XDFFPOSX1_464 NAND3X1_54/A CLKBUF1_27/Y BUFX2_63/A gnd vdd DFFPOSX1
XDFFPOSX1_475 BUFX2_42/A CLKBUF1_10/Y NAND3X1_13/Y gnd vdd DFFPOSX1
XDFFPOSX1_486 BUFX2_53/A CLKBUF1_41/Y NAND3X1_35/Y gnd vdd DFFPOSX1
XNAND2X1_501 INVX8_3/A OR2X2_26/A gnd NAND2X1_501/Y vdd NAND2X1
XNAND2X1_512 INVX8_7/A NOR2X1_369/A gnd OAI21X1_567/C vdd NAND2X1
XDFFPOSX1_497 BUFX2_64/A CLKBUF1_36/Y NAND3X1_57/Y gnd vdd DFFPOSX1
XNAND2X1_545 INVX1_403/A NOR2X1_316/Y gnd NAND3X1_144/C vdd NAND2X1
XNAND2X1_534 NOR2X1_302/Y NOR2X1_304/Y gnd OAI21X1_603/B vdd NAND2X1
XNAND2X1_523 BUFX4_127/Y NOR2X1_373/B gnd NAND2X1_523/Y vdd NAND2X1
XNAND2X1_556 INVX8_4/A NAND2X1_556/B gnd NAND2X1_556/Y vdd NAND2X1
XNAND2X1_567 INVX8_7/A NOR2X1_237/Y gnd NAND2X1_567/Y vdd NAND2X1
XNAND2X1_578 NOR2X1_82/Y AOI21X1_203/B gnd NAND2X1_578/Y vdd NAND2X1
XNAND2X1_589 INVX8_5/A MUX2X1_48/Y gnd OAI21X1_737/C vdd NAND2X1
XFILL_40_5_1 gnd vdd FILL
XAOI21X1_180 NOR2X1_337/Y AOI21X1_180/B AOI21X1_180/C gnd OAI21X1_698/B vdd AOI21X1
XAOI21X1_191 INVX2_19/Y AND2X2_64/B NOR2X1_78/Y gnd OAI21X1_722/C vdd AOI21X1
XNAND3X1_140 AOI22X1_97/D NOR2X1_281/A AOI22X1_99/Y gnd NOR2X1_296/B vdd NAND3X1
XFILL_31_5_1 gnd vdd FILL
XNAND3X1_184 AND2X2_78/Y INVX1_487/A NOR3X1_65/Y gnd NOR3X1_68/C vdd NAND3X1
XNAND3X1_151 NAND3X1_151/A OAI21X1_647/Y NOR3X1_59/Y gnd INVX1_86/A vdd NAND3X1
XNAND3X1_162 NAND2X1_581/Y NAND3X1_162/B NAND3X1_162/C gnd AOI21X1_189/C vdd NAND3X1
XNAND3X1_173 NAND3X1_173/A NAND3X1_172/Y AOI21X1_210/Y gnd INVX1_96/A vdd NAND3X1
XFILL_30_0_0 gnd vdd FILL
XNAND3X1_195 BUFX4_219/Y NAND3X1_194/Y NAND3X1_195/C gnd NAND2X1_717/B vdd NAND3X1
XFILL_39_6_1 gnd vdd FILL
XFILL_38_1_0 gnd vdd FILL
XFILL_22_5_1 gnd vdd FILL
XOAI21X1_303 OAI21X1_302/Y OR2X2_39/B AOI21X1_37/Y gnd AOI21X1_39/A vdd OAI21X1
XOAI21X1_314 INVX1_337/Y INVX4_4/A NAND2X1_261/Y gnd NOR2X1_125/B vdd OAI21X1
XFILL_21_0_0 gnd vdd FILL
XOAI21X1_325 INVX2_47/Y AOI22X1_88/C AOI21X1_88/A gnd AOI21X1_41/B vdd OAI21X1
XOAI21X1_347 BUFX4_43/Y MUX2X1_3/Y NAND2X1_328/Y gnd NAND2X1_400/B vdd OAI21X1
XOAI21X1_336 AOI22X1_75/Y INVX1_311/A OAI21X1_333/Y gnd AOI21X1_45/B vdd OAI21X1
XOAI21X1_369 AOI21X1_54/B BUFX4_124/Y INVX4_5/Y gnd OAI21X1_370/C vdd OAI21X1
XOAI21X1_358 AOI21X1_53/Y BUFX4_225/Y OAI21X1_357/Y gnd MUX2X1_26/A vdd OAI21X1
XBUFX4_1 CLK gnd BUFX4_1/Y vdd BUFX4
XDFFPOSX1_272 MUX2X1_2/A CLKBUF1_52/Y NAND3X1_42/A gnd vdd DFFPOSX1
XDFFPOSX1_261 INVX1_251/A CLKBUF1_26/Y NAND3X1_20/A gnd vdd DFFPOSX1
XDFFPOSX1_250 OAI21X1_153/C CLKBUF1_60/Y INVX1_94/A gnd vdd DFFPOSX1
XNAND2X1_320 INVX4_4/A INVX1_350/Y gnd AOI21X1_47/B vdd NAND2X1
XDFFPOSX1_283 AOI22X1_66/A CLKBUF1_36/Y NAND3X1_64/A gnd vdd DFFPOSX1
XDFFPOSX1_294 INVX2_49/A CLKBUF1_12/Y NOR3X1_10/Y gnd vdd DFFPOSX1
XXOR2X1_14 BUFX2_91/A INVX2_3/A gnd XOR2X1_14/Y vdd XOR2X1
XNAND2X1_342 BUFX4_217/Y NAND2X1_342/B gnd NAND2X1_342/Y vdd NAND2X1
XNAND2X1_331 INVX8_4/A NAND2X1_427/B gnd OAI21X1_353/C vdd NAND2X1
XNAND2X1_353 INVX1_347/Y AND2X2_23/Y gnd NOR2X1_180/A vdd NAND2X1
XNAND2X1_375 BUFX4_52/Y INVX1_365/Y gnd NAND2X1_375/Y vdd NAND2X1
XFILL_5_6_1 gnd vdd FILL
XNAND2X1_386 BUFX4_43/Y MUX2X1_39/A gnd OAI21X1_583/C vdd NAND2X1
XNAND2X1_364 INVX8_8/A INVX2_21/A gnd OAI21X1_378/C vdd NAND2X1
XFILL_4_1_0 gnd vdd FILL
XNAND2X1_397 INVX8_5/A NOR2X1_201/Y gnd OAI21X1_411/C vdd NAND2X1
XFILL_29_1_0 gnd vdd FILL
XNOR3X1_60 NOR3X1_60/A NOR3X1_60/B NOR3X1_60/C gnd NOR3X1_60/Y vdd NOR3X1
XNOR3X1_71 NOR3X1_71/A NOR3X1_71/B NOR3X1_71/C gnd NOR3X1_71/Y vdd NOR3X1
XFILL_13_5_1 gnd vdd FILL
XFILL_12_0_0 gnd vdd FILL
XINVX4_1 INVX4_1/A gnd INVX4_1/Y vdd INVX4
XOAI21X1_870 INVX1_495/A INVX1_567/Y NAND2X1_805/Y gnd AOI21X1_225/C vdd OAI21X1
XOAI21X1_892 INVX8_14/Y AOI21X1_231/Y OAI21X1_892/C gnd OAI21X1_892/Y vdd OAI21X1
XOAI21X1_881 INVX8_14/Y INVX1_643/A NAND2X1_925/Y gnd OAI21X1_881/Y vdd OAI21X1
XNAND3X1_4 INVX1_138/Y INVX1_572/A NOR2X1_6/Y gnd NOR2X1_7/B vdd NAND3X1
XOAI21X1_100 BUFX4_186/Y INVX1_100/Y OAI21X1_99/Y gnd INVX1_579/A vdd OAI21X1
XOAI21X1_122 BUFX4_183/Y INVX1_111/Y OAI21X1_121/Y gnd INVX1_601/A vdd OAI21X1
XOAI21X1_111 BUFX4_269/Y BUFX4_192/Y OAI21X1_111/C gnd OAI21X1_111/Y vdd OAI21X1
XAOI22X1_9 AOI22X1_9/A AOI22X1_9/B OR2X2_3/A AOI22X1_9/D gnd AOI22X1_9/Y vdd AOI22X1
XOAI21X1_144 BUFX4_182/Y INVX1_122/Y OAI21X1_144/C gnd INVX1_623/A vdd OAI21X1
XOAI21X1_133 BUFX4_270/Y OR2X2_2/B OAI21X1_133/C gnd OAI21X1_133/Y vdd OAI21X1
XOAI21X1_155 OR2X2_2/A BUFX4_194/Y OAI21X1_155/C gnd OAI21X1_155/Y vdd OAI21X1
XOAI21X1_177 BUFX4_12/Y BUFX4_197/Y OAI21X1_840/Y gnd NAND3X1_39/C vdd OAI21X1
XOAI21X1_166 BUFX4_15/Y BUFX4_200/Y OAI21X1_821/Y gnd NAND3X1_17/C vdd OAI21X1
XOAI21X1_188 BUFX4_13/Y BUFX4_196/Y OAI21X1_861/Y gnd NAND3X1_61/C vdd OAI21X1
XINVX1_208 INVX1_208/A gnd INVX1_208/Y vdd INVX1
XOAI21X1_199 BUFX4_145/Y INVX1_197/Y AOI22X1_14/Y gnd OAI21X1_199/Y vdd OAI21X1
XINVX1_219 INVX1_219/A gnd INVX1_219/Y vdd INVX1
XNAND2X1_150 NOR2X1_38/Y NOR2X1_39/Y gnd AOI21X1_26/C vdd NAND2X1
XNAND2X1_161 AOI21X1_27/A OR2X2_10/Y gnd OR2X2_11/B vdd NAND2X1
XNAND2X1_19 BUFX4_19/Y NAND2X1_19/B gnd OAI21X1_19/C vdd NAND2X1
XNAND2X1_172 NAND2X1_172/A OR2X2_14/Y gnd XOR2X1_5/B vdd NAND2X1
XNAND2X1_194 INVX1_66/A AND2X2_20/Y gnd NOR2X1_71/A vdd NAND2X1
XNAND2X1_183 INVX1_283/Y NOR2X1_55/B gnd AOI21X1_30/A vdd NAND2X1
XAOI22X1_39 AOI22X1_39/A AOI22X1_9/B OR2X2_3/A AOI22X1_39/D gnd AOI22X1_39/Y vdd AOI22X1
XAOI22X1_17 AOI22X1_17/A BUFX4_236/Y BUFX4_258/Y AOI22X1_17/D gnd AOI22X1_17/Y vdd
+ AOI22X1
XAOI22X1_28 AOI22X1_28/A OR2X2_3/B BUFX4_257/Y AOI22X1_28/D gnd AOI22X1_28/Y vdd AOI22X1
XNOR3X1_7 NOR3X1_9/A NOR3X1_7/B NOR3X1_9/C gnd NOR3X1_7/Y vdd NOR3X1
XINVX1_720 INVX1_720/A gnd INVX1_720/Y vdd INVX1
XINVX1_742 data_memory_interface_data[10] gnd INVX1_742/Y vdd INVX1
XINVX1_731 INVX1_731/A gnd INVX1_731/Y vdd INVX1
XINVX1_753 INVX1_753/A gnd INVX1_753/Y vdd INVX1
XFILL_5_1 gnd vdd FILL
XXNOR2X1_50 INVX1_470/A INVX2_72/Y gnd XNOR2X1_50/Y vdd XNOR2X1
XFILL_36_4_1 gnd vdd FILL
XBUFX2_71 BUFX4_75/Y gnd instruction_memory_interface_enable vdd BUFX2
XBUFX2_60 BUFX2_60/A gnd instruction_memory_interface_address[21] vdd BUFX2
XBUFX2_93 BUFX2_93/A gnd BUFX2_93/Y vdd BUFX2
XBUFX2_82 BUFX2_82/A gnd BUFX2_82/Y vdd BUFX2
XFILL_2_4_1 gnd vdd FILL
XFILL_27_4_1 gnd vdd FILL
XFILL_10_3_1 gnd vdd FILL
XAOI21X1_50 AOI21X1_50/A INVX2_52/Y INVX8_5/A gnd AOI21X1_50/Y vdd AOI21X1
XAOI21X1_61 BUFX4_83/Y NOR2X1_205/B INVX8_3/A gnd NOR2X1_204/A vdd AOI21X1
XAOI21X1_72 INVX1_373/A INVX8_11/Y AOI21X1_72/C gnd AOI21X1_72/Y vdd AOI21X1
XAOI21X1_83 AND2X2_55/A INVX4_6/Y AOI21X1_83/C gnd AOI21X1_83/Y vdd AOI21X1
XAOI21X1_94 AND2X2_36/B BUFX4_189/Y AOI21X1_94/C gnd AOI21X1_94/Y vdd AOI21X1
XOAI21X1_1 INVX1_1/Y BUFX4_23/Y OAI21X1_1/C gnd OAI21X1_1/Y vdd OAI21X1
XFILL_9_0_0 gnd vdd FILL
XFILL_18_4_1 gnd vdd FILL
XNOR2X1_407 NOR2X1_407/A OAI22X1_48/Y gnd NOR2X1_407/Y vdd NOR2X1
XNOR2X1_429 MUX2X1_3/B INVX1_676/Y gnd NOR2X1_429/Y vdd NOR2X1
XNOR2X1_418 INVX1_653/Y BUFX4_260/Y gnd NOR2X1_418/Y vdd NOR2X1
XINVX1_561 INVX1_561/A gnd INVX1_561/Y vdd INVX1
XINVX1_550 INVX1_623/A gnd INVX1_550/Y vdd INVX1
XINVX1_572 INVX1_572/A gnd INVX1_572/Y vdd INVX1
XNAND2X1_919 OAI22X1_49/A OAI21X1_887/B gnd OAI22X1_49/C vdd NAND2X1
XNAND2X1_908 NAND2X1_906/Y NAND2X1_908/B gnd NAND2X1_62/B vdd NAND2X1
XINVX1_583 INVX1_583/A gnd INVX1_583/Y vdd INVX1
XINVX1_594 INVX1_521/A gnd INVX1_594/Y vdd INVX1
XXOR2X1_4 XOR2X1_4/A OR2X2_11/A gnd XOR2X1_4/Y vdd XOR2X1
XFILL_42_2_1 gnd vdd FILL
XMUX2X1_5 MUX2X1_5/A OR2X2_57/A INVX4_4/A gnd MUX2X1_5/Y vdd MUX2X1
XCLKBUF1_6 BUFX4_5/Y gnd CLKBUF1_6/Y vdd CLKBUF1
XBUFX4_111 NOR2X1_7/Y gnd BUFX4_111/Y vdd BUFX4
XAOI22X1_171 BUFX4_252/Y INVX1_733/A AOI22X1_171/C BUFX4_106/Y gnd AOI22X1_171/Y vdd
+ AOI22X1
XBUFX4_100 BUFX4_99/A gnd BUFX4_100/Y vdd BUFX4
XAOI22X1_160 data_memory_interface_data[24] BUFX4_109/Y BUFX4_171/Y BUFX4_251/Y gnd
+ AOI22X1_160/Y vdd AOI22X1
XBUFX4_155 BUFX4_152/A gnd BUFX4_155/Y vdd BUFX4
XBUFX4_144 OR2X2_3/Y gnd BUFX4_144/Y vdd BUFX4
XBUFX4_133 AND2X2_79/Y gnd BUFX4_133/Y vdd BUFX4
XBUFX4_122 BUFX4_122/A gnd BUFX4_122/Y vdd BUFX4
XNOR2X1_215 BUFX4_176/Y INVX1_374/A gnd AOI22X1_80/D vdd NOR2X1
XNOR2X1_204 NOR2X1_204/A INVX1_371/Y gnd NOR2X1_204/Y vdd NOR2X1
XBUFX4_188 BUFX4_188/A gnd INVX8_12/A vdd BUFX4
XBUFX4_177 BUFX4_178/A gnd BUFX4_177/Y vdd BUFX4
XBUFX4_166 BUFX4_164/A gnd BUFX4_166/Y vdd BUFX4
XNOR2X1_248 INVX2_44/Y MUX2X1_9/Y gnd NOR2X1_248/Y vdd NOR2X1
XBUFX4_199 INVX8_2/Y gnd BUFX4_199/Y vdd BUFX4
XNOR2X1_237 BUFX4_176/Y INVX1_385/Y gnd NOR2X1_237/Y vdd NOR2X1
XNOR2X1_226 INVX8_9/A INVX1_371/Y gnd INVX1_388/A vdd NOR2X1
XNOR2X1_259 INVX8_3/A AND2X2_29/A gnd NOR2X1_259/Y vdd NOR2X1
XFILL_33_2_1 gnd vdd FILL
XOAI21X1_1001 INVX1_747/Y OAI21X1_993/B NAND2X1_1016/Y gnd AOI22X1_142/C vdd OAI21X1
XOAI21X1_1012 AND2X2_99/B INVX2_88/A INVX8_15/A gnd INVX1_753/A vdd OAI21X1
XOAI21X1_1045 BUFX4_67/Y BUFX4_70/Y AOI22X1_161/Y gnd OAI21X1_1045/Y vdd OAI21X1
XOAI21X1_1034 INVX1_755/Y INVX2_93/A OAI21X1_1034/C gnd BUFX4_171/A vdd OAI21X1
XOAI21X1_1023 INVX1_745/Y INVX2_93/A OAI21X1_1022/Y gnd AOI22X1_147/C vdd OAI21X1
XOAI21X1_1056 NOR2X1_481/Y INVX4_12/A BUFX4_11/Y gnd AOI21X1_270/C vdd OAI21X1
XOAI21X1_1067 AOI21X1_271/Y OAI21X1_1066/Y NOR2X1_487/Y gnd OAI21X1_1067/Y vdd OAI21X1
XINVX1_380 INVX1_242/A gnd INVX1_380/Y vdd INVX1
XNAND2X1_705 OR2X2_50/A OR2X2_50/B gnd NAND2X1_705/Y vdd NAND2X1
XINVX1_391 INVX1_391/A gnd INVX1_391/Y vdd INVX1
XNAND2X1_727 OAI21X1_71/Y BUFX4_135/Y gnd NAND2X1_727/Y vdd NAND2X1
XNAND2X1_716 INVX1_507/Y BUFX4_201/Y gnd NAND3X1_195/C vdd NAND2X1
XNAND2X1_738 NAND2X1_738/A NAND2X1_738/B gnd NAND2X1_10/B vdd NAND2X1
XNAND2X1_749 INVX1_529/Y BUFX4_205/Y gnd NAND3X1_217/C vdd NAND2X1
XFILL_24_2_1 gnd vdd FILL
XINVX8_8 INVX8_8/A gnd INVX8_8/Y vdd INVX8
XDFFPOSX1_61 AOI22X1_23/A CLKBUF1_15/Y INVX1_114/A gnd vdd DFFPOSX1
XDFFPOSX1_50 AOI22X1_12/A CLKBUF1_30/Y INVX1_103/A gnd vdd DFFPOSX1
XDFFPOSX1_72 AOI22X1_34/A CLKBUF1_3/Y INVX1_125/A gnd vdd DFFPOSX1
XDFFPOSX1_83 INVX1_196/A CLKBUF1_31/Y DFFPOSX1_83/D gnd vdd DFFPOSX1
XDFFPOSX1_94 INVX1_207/A CLKBUF1_3/Y OAI21X1_129/C gnd vdd DFFPOSX1
XFILL_7_3_1 gnd vdd FILL
XBUFX4_17 BUFX4_22/A gnd BUFX4_17/Y vdd BUFX4
XBUFX4_39 INVX8_8/Y gnd BUFX4_39/Y vdd BUFX4
XBUFX4_28 BUFX4_27/A gnd BUFX4_28/Y vdd BUFX4
XFILL_15_2_1 gnd vdd FILL
XNAND3X1_322 INVX1_639/Y BUFX4_103/Y BUFX4_164/Y gnd NAND3X1_322/Y vdd NAND3X1
XNAND3X1_300 INVX1_617/Y BUFX4_103/Y BUFX4_164/Y gnd NAND3X1_300/Y vdd NAND3X1
XNAND3X1_333 AND2X2_86/Y NOR2X1_430/Y NAND3X1_341/B gnd INVX1_691/A vdd NAND3X1
XNAND3X1_311 BUFX4_120/Y NAND3X1_311/B NAND3X1_311/C gnd NAND2X1_896/B vdd NAND3X1
XNAND3X1_355 NAND3X1_349/A OAI22X1_58/B INVX2_93/A gnd BUFX2_36/A vdd NAND3X1
XNAND3X1_344 INVX2_88/Y INVX2_89/Y AND2X2_98/Y gnd NOR3X1_79/A vdd NAND3X1
XOAI21X1_507 OAI21X1_366/Y BUFX4_54/Y NAND2X1_473/Y gnd NOR2X1_241/B vdd OAI21X1
XOAI21X1_529 NAND3X1_123/C INVX2_58/A OAI21X1_529/C gnd AND2X2_41/A vdd OAI21X1
XOAI21X1_518 BUFX4_229/Y MUX2X1_31/Y OAI21X1_518/C gnd INVX1_395/A vdd OAI21X1
XDFFPOSX1_421 BUFX2_85/A CLKBUF1_44/Y NOR3X1_28/Y gnd vdd DFFPOSX1
XDFFPOSX1_410 NOR2X1_18/A CLKBUF1_20/Y NOR3X1_18/Y gnd vdd DFFPOSX1
XDFFPOSX1_443 NAND3X1_12/A CLKBUF1_54/Y BUFX2_42/A gnd vdd DFFPOSX1
XDFFPOSX1_454 NAND3X1_34/A CLKBUF1_26/Y BUFX2_53/A gnd vdd DFFPOSX1
XDFFPOSX1_465 NAND3X1_56/A CLKBUF1_47/Y BUFX2_64/A gnd vdd DFFPOSX1
XDFFPOSX1_432 BUFX2_91/A CLKBUF1_13/Y NOR3X1_39/Y gnd vdd DFFPOSX1
XNAND2X1_502 INVX8_4/A NAND2X1_472/B gnd NAND2X1_502/Y vdd NAND2X1
XDFFPOSX1_476 BUFX2_43/A CLKBUF1_33/Y NAND3X1_15/Y gnd vdd DFFPOSX1
XDFFPOSX1_487 BUFX2_54/A CLKBUF1_41/Y NAND3X1_37/Y gnd vdd DFFPOSX1
XDFFPOSX1_498 BUFX2_65/A CLKBUF1_6/Y NAND3X1_59/Y gnd vdd DFFPOSX1
XNAND2X1_535 AND2X2_52/A AOI21X1_185/B gnd OAI21X1_604/C vdd NAND2X1
XNAND2X1_524 INVX2_38/Y MUX2X1_39/A gnd AOI22X1_99/A vdd NAND2X1
XNAND2X1_513 INVX1_394/Y NOR2X1_283/Y gnd OAI22X1_30/C vdd NAND2X1
XNAND2X1_546 INVX8_3/A MUX2X1_34/A gnd OAI21X1_634/C vdd NAND2X1
XNAND2X1_557 BUFX4_228/Y MUX2X1_47/B gnd NAND2X1_557/Y vdd NAND2X1
XNAND2X1_579 INVX8_3/A OAI21X1_719/A gnd NAND2X1_579/Y vdd NAND2X1
XNAND2X1_568 OAI21X1_689/Y AOI22X1_103/Y gnd AOI21X1_174/C vdd NAND2X1
XAOI21X1_170 AOI21X1_170/A AOI21X1_170/B INVX2_65/Y gnd NOR3X1_60/A vdd AOI21X1
XAOI21X1_192 INVX2_18/A OAI21X1_722/Y BUFX4_276/Y gnd OAI21X1_723/C vdd AOI21X1
XAOI21X1_181 NOR2X1_81/Y OAI21X1_698/B BUFX4_88/Y gnd AOI21X1_181/Y vdd AOI21X1
XNAND3X1_141 OAI21X1_591/Y OAI21X1_595/Y NOR2X1_300/Y gnd INVX1_82/A vdd NAND3X1
XNAND3X1_130 INVX8_11/Y NAND3X1_129/Y NAND3X1_130/C gnd NAND3X1_130/Y vdd NAND3X1
XNAND3X1_152 NAND3X1_152/A AOI21X1_165/Y OAI21X1_665/Y gnd NAND3X1_152/Y vdd NAND3X1
XNAND3X1_163 NAND3X1_163/A NAND3X1_161/Y AOI21X1_189/Y gnd NAND3X1_163/Y vdd NAND3X1
XNAND3X1_174 INVX2_26/Y INVX1_430/Y NAND3X1_174/C gnd NAND3X1_175/B vdd NAND3X1
XFILL_30_0_1 gnd vdd FILL
XNAND3X1_185 INVX1_491/Y INVX1_492/Y NOR3X1_66/Y gnd NOR2X1_398/B vdd NAND3X1
XNAND3X1_196 INVX1_510/Y BUFX4_207/Y BUFX4_35/Y gnd NAND3X1_197/B vdd NAND3X1
XFILL_38_1_1 gnd vdd FILL
XOAI21X1_304 NOR2X1_101/Y NOR2X1_102/Y INVX1_411/A gnd OAI21X1_305/B vdd OAI21X1
XFILL_21_0_1 gnd vdd FILL
XOAI21X1_315 INVX1_338/Y INVX4_4/A NAND2X1_266/Y gnd MUX2X1_24/B vdd OAI21X1
XOAI21X1_326 AOI21X1_40/Y NAND3X1_91/Y AOI21X1_41/Y gnd AOI21X1_43/B vdd OAI21X1
XOAI21X1_337 INVX1_315/Y INVX2_27/A INVX2_26/Y gnd AOI21X1_45/C vdd OAI21X1
XOAI21X1_348 BUFX4_42/Y MUX2X1_6/Y OAI21X1_348/C gnd INVX1_353/A vdd OAI21X1
XOAI21X1_359 MUX2X1_19/Y MUX2X1_20/S OAI21X1_359/C gnd AND2X2_38/A vdd OAI21X1
XDFFPOSX1_240 OAI21X1_133/C CLKBUF1_23/Y INVX1_84/A gnd vdd DFFPOSX1
XBUFX4_2 CLK gnd BUFX4_2/Y vdd BUFX4
XDFFPOSX1_262 MUX2X1_10/A CLKBUF1_14/Y NAND3X1_22/A gnd vdd DFFPOSX1
XDFFPOSX1_273 MUX2X1_1/A CLKBUF1_52/Y NAND3X1_44/A gnd vdd DFFPOSX1
XDFFPOSX1_251 OAI21X1_155/C CLKBUF1_23/Y INVX1_95/A gnd vdd DFFPOSX1
XNAND2X1_310 INVX1_346/Y AND2X2_20/Y gnd OR2X2_16/A vdd NAND2X1
XDFFPOSX1_284 AOI22X1_67/A CLKBUF1_17/Y NAND3X1_66/A gnd vdd DFFPOSX1
XDFFPOSX1_295 AND2X2_93/B CLKBUF1_13/Y NOR3X1_11/Y gnd vdd DFFPOSX1
XXOR2X1_15 OR2X2_52/B INVX2_2/A gnd XOR2X1_15/Y vdd XOR2X1
XNAND2X1_332 BUFX4_42/Y NOR2X1_123/B gnd OAI21X1_350/C vdd NAND2X1
XNAND2X1_321 INVX4_4/Y INVX1_339/Y gnd AOI21X1_48/B vdd NAND2X1
XNAND2X1_343 NOR2X1_165/Y NOR2X1_171/Y gnd BUFX4_175/A vdd NAND2X1
XNAND2X1_354 MUX2X1_13/A INVX4_4/A gnd OAI21X1_372/C vdd NAND2X1
XNAND2X1_387 BUFX4_43/Y MUX2X1_37/A gnd OAI21X1_403/C vdd NAND2X1
XNAND2X1_376 BUFX4_82/Y OAI21X1_391/Y gnd NOR2X1_311/B vdd NAND2X1
XNAND2X1_365 INVX8_8/A INVX2_17/A gnd NAND2X1_365/Y vdd NAND2X1
XFILL_4_1_1 gnd vdd FILL
XNAND2X1_398 BUFX4_58/Y AND2X2_44/A gnd NAND2X1_398/Y vdd NAND2X1
XFILL_29_1_1 gnd vdd FILL
XNOR3X1_50 NOR3X1_50/A AOI21X1_4/C NOR3X1_49/C gnd NOR3X1_50/Y vdd NOR3X1
XNOR3X1_61 AND2X2_60/Y NOR3X1_61/B NOR3X1_61/C gnd NOR3X1_61/Y vdd NOR3X1
XNOR3X1_72 NOR3X1_72/A NOR3X1_72/B NOR3X1_72/C gnd NOR3X1_72/Y vdd NOR3X1
XFILL_12_0_1 gnd vdd FILL
XINVX4_2 INVX4_2/A gnd INVX4_2/Y vdd INVX4
XOAI21X1_860 NAND2X1_689/Y INVX1_491/A INVX8_13/Y gnd OAI21X1_860/Y vdd OAI21X1
XOAI21X1_871 INVX2_73/Y DFFPOSX1_41/Q OAI21X1_871/C gnd NOR2X1_404/B vdd OAI21X1
XOAI21X1_893 INVX8_14/Y AOI21X1_231/Y OAI21X1_893/C gnd OAI21X1_893/Y vdd OAI21X1
XOAI21X1_882 OAI22X1_6/Y INVX2_79/Y INVX4_11/A gnd OAI21X1_882/Y vdd OAI21X1
XNAND3X1_5 INVX4_1/Y INVX1_149/Y NAND3X1_7/C gnd NAND3X1_5/Y vdd NAND3X1
XOAI21X1_101 BUFX4_273/Y BUFX4_193/Y OAI21X1_101/C gnd OAI21X1_102/C vdd OAI21X1
XOAI21X1_112 BUFX4_184/Y INVX1_106/Y OAI21X1_111/Y gnd INVX1_591/A vdd OAI21X1
XOAI21X1_123 BUFX4_273/Y BUFX4_193/Y OAI21X1_123/C gnd OAI21X1_123/Y vdd OAI21X1
XOAI21X1_145 BUFX4_269/Y BUFX4_192/Y OAI21X1_145/C gnd OAI21X1_145/Y vdd OAI21X1
XOAI21X1_134 BUFX4_185/Y INVX1_117/Y OAI21X1_133/Y gnd INVX1_613/A vdd OAI21X1
XOAI21X1_156 BUFX4_186/Y INVX1_128/Y OAI21X1_155/Y gnd INVX1_635/A vdd OAI21X1
XOAI21X1_167 BUFX4_12/Y BUFX4_199/Y OAI21X1_167/C gnd NAND3X1_19/C vdd OAI21X1
XOAI21X1_178 BUFX4_14/Y BUFX4_197/Y OAI21X1_178/C gnd NAND3X1_41/C vdd OAI21X1
XOAI21X1_189 BUFX4_13/Y BUFX4_196/Y OAI21X1_862/Y gnd NAND3X1_63/C vdd OAI21X1
XINVX1_209 INVX1_209/A gnd INVX1_209/Y vdd INVX1
XNAND2X1_140 INVX1_253/Y AOI21X1_15/Y gnd NAND2X1_140/Y vdd NAND2X1
XNAND2X1_151 INVX2_14/Y NOR2X1_41/B gnd AOI21X1_24/A vdd NAND2X1
XNAND2X1_162 MUX2X1_1/B BUFX4_146/Y gnd NAND3X1_84/C vdd NAND2X1
XNAND2X1_173 INVX1_276/A INVX1_275/Y gnd AND2X2_16/B vdd NAND2X1
XNAND2X1_195 NOR2X1_6/A NOR2X1_70/Y gnd NOR2X1_71/B vdd NAND2X1
XNAND2X1_184 AOI21X1_30/A INVX1_284/Y gnd NOR2X1_57/A vdd NAND2X1
XAOI22X1_18 AOI22X1_18/A BUFX4_236/Y BUFX4_258/Y AOI22X1_18/D gnd AOI22X1_18/Y vdd
+ AOI22X1
XAOI22X1_29 AOI22X1_29/A OR2X2_3/B BUFX4_257/Y AOI22X1_29/D gnd AOI22X1_29/Y vdd AOI22X1
XOAI21X1_690 OR2X2_40/A INVX1_382/A OAI21X1_690/C gnd NOR3X1_61/C vdd OAI21X1
XINVX1_710 INVX1_710/A gnd INVX1_710/Y vdd INVX1
XNOR3X1_8 INVX4_1/A NOR3X1_8/B NOR3X1_8/C gnd NOR3X1_8/Y vdd NOR3X1
XINVX1_721 INVX1_721/A gnd INVX1_721/Y vdd INVX1
XINVX1_743 data_memory_interface_data[3] gnd INVX1_743/Y vdd INVX1
XINVX1_732 INVX1_732/A gnd INVX1_732/Y vdd INVX1
XINVX1_754 data_memory_interface_data[30] gnd INVX1_754/Y vdd INVX1
XFILL_5_2 gnd vdd FILL
XXNOR2X1_40 INVX1_272/A NOR2X1_45/A gnd XNOR2X1_40/Y vdd XNOR2X1
XXNOR2X1_51 XNOR2X1_51/A BUFX2_53/A gnd XNOR2X1_51/Y vdd XNOR2X1
XBUFX2_72 vdd gnd instruction_memory_interface_frame_mask[0] vdd BUFX2
XBUFX2_50 BUFX2_50/A gnd instruction_memory_interface_address[11] vdd BUFX2
XBUFX2_61 BUFX2_61/A gnd instruction_memory_interface_address[22] vdd BUFX2
XBUFX2_94 BUFX2_94/A gnd BUFX2_94/Y vdd BUFX2
XBUFX2_83 BUFX2_83/A gnd BUFX2_83/Y vdd BUFX2
XAOI21X1_40 AOI21X1_77/A AOI21X1_40/B AOI21X1_40/C gnd AOI21X1_40/Y vdd AOI21X1
XAOI21X1_51 BUFX4_41/Y MUX2X1_30/B AOI21X1_93/C gnd AOI21X1_51/Y vdd AOI21X1
XAOI21X1_62 AOI21X1_48/A AOI21X1_48/B BUFX4_213/Y gnd AOI21X1_62/Y vdd AOI21X1
XAOI21X1_95 INVX1_387/Y INVX4_6/Y AOI21X1_95/C gnd AOI21X1_95/Y vdd AOI21X1
XAOI21X1_73 INVX1_374/Y INVX4_6/Y AOI21X1_73/C gnd AOI21X1_73/Y vdd AOI21X1
XAOI21X1_84 INVX2_47/A OR2X2_28/A BUFX4_86/Y gnd AOI21X1_84/Y vdd AOI21X1
XOAI21X1_2 INVX1_2/Y BUFX4_23/Y OAI21X1_2/C gnd OAI21X1_2/Y vdd OAI21X1
XFILL_9_0_1 gnd vdd FILL
XNOR2X1_419 NOR2X1_419/A NOR2X1_419/B gnd INVX1_714/A vdd NOR2X1
XNOR2X1_408 NOR2X1_408/A NOR2X1_408/B gnd BUFX4_164/A vdd NOR2X1
XINVX1_551 INVX1_551/A gnd INVX1_551/Y vdd INVX1
XINVX1_540 INVX1_613/A gnd INVX1_540/Y vdd INVX1
XINVX1_562 INVX1_635/A gnd INVX1_562/Y vdd INVX1
XNAND2X1_909 OAI21X1_95/Y BUFX4_61/Y gnd NAND2X1_909/Y vdd NAND2X1
XINVX1_595 INVX1_595/A gnd INVX1_595/Y vdd INVX1
XINVX1_573 INVX1_500/A gnd INVX1_573/Y vdd INVX1
XINVX1_584 INVX1_511/A gnd INVX1_584/Y vdd INVX1
XFILL_37_7_0 gnd vdd FILL
XFILL_20_6_0 gnd vdd FILL
XFILL_3_7_0 gnd vdd FILL
XXOR2X1_5 XOR2X1_5/A XOR2X1_5/B gnd XOR2X1_5/Y vdd XOR2X1
XFILL_28_7_0 gnd vdd FILL
XMUX2X1_6 MUX2X1_6/A MUX2X1_6/B INVX4_4/A gnd MUX2X1_6/Y vdd MUX2X1
XFILL_11_6_0 gnd vdd FILL
XCLKBUF1_7 BUFX4_3/Y gnd CLKBUF1_7/Y vdd CLKBUF1
XBUFX4_112 NOR2X1_7/Y gnd AND2X2_2/B vdd BUFX4
XAOI22X1_161 data_memory_interface_data[25] BUFX4_109/Y BUFX4_170/Y BUFX4_251/Y gnd
+ AOI22X1_161/Y vdd AOI22X1
XAOI22X1_150 data_memory_interface_data[14] BUFX4_105/Y AOI22X1_150/C BUFX4_10/Y gnd
+ AOI22X1_150/Y vdd AOI22X1
XBUFX4_101 BUFX4_99/A gnd BUFX4_101/Y vdd BUFX4
XFILL_19_7_0 gnd vdd FILL
XBUFX4_134 AND2X2_79/Y gnd BUFX4_134/Y vdd BUFX4
XBUFX4_145 OR2X2_3/Y gnd BUFX4_145/Y vdd BUFX4
XBUFX4_123 BUFX4_122/A gnd BUFX4_123/Y vdd BUFX4
XNOR2X1_216 INVX8_3/A OR2X2_30/B gnd INVX2_55/A vdd NOR2X1
XNOR2X1_205 INVX8_3/A NOR2X1_205/B gnd NOR2X1_205/Y vdd NOR2X1
XBUFX4_178 BUFX4_178/A gnd BUFX4_178/Y vdd BUFX4
XBUFX4_156 NOR2X1_2/Y gnd BUFX4_156/Y vdd BUFX4
XBUFX4_167 BUFX4_164/A gnd BUFX4_167/Y vdd BUFX4
XNOR2X1_249 INVX2_44/A NOR2X1_249/B gnd NOR2X1_249/Y vdd NOR2X1
XNOR2X1_238 INVX8_3/A NOR2X1_238/B gnd NOR2X1_238/Y vdd NOR2X1
XBUFX4_189 BUFX4_188/A gnd BUFX4_189/Y vdd BUFX4
XNOR2X1_227 NOR2X1_229/B INVX4_6/A gnd NOR2X1_227/Y vdd NOR2X1
XOAI21X1_1002 AOI21X1_263/Y OAI21X1_994/B AOI22X1_142/Y gnd OAI21X1_1002/Y vdd OAI21X1
XOAI21X1_1013 OAI21X1_1009/A NOR3X1_81/Y OAI22X1_60/C gnd AOI21X1_266/B vdd OAI21X1
XOAI21X1_1035 BUFX4_67/Y BUFX4_70/Y AOI22X1_151/Y gnd OAI21X1_1035/Y vdd OAI21X1
XOAI21X1_1046 BUFX4_67/Y BUFX4_70/Y AOI22X1_162/Y gnd OAI21X1_1046/Y vdd OAI21X1
XOAI21X1_1024 BUFX4_65/Y BUFX4_69/Y AOI22X1_147/Y gnd OAI21X1_1024/Y vdd OAI21X1
XOAI21X1_1057 INVX4_13/A INVX2_90/Y INVX1_753/A gnd OAI21X1_1057/Y vdd OAI21X1
XOAI21X1_1068 INVX1_759/Y INVX2_90/Y INVX1_757/A gnd OAI21X1_1069/B vdd OAI21X1
XINVX1_370 INVX1_370/A gnd INVX1_370/Y vdd INVX1
XINVX1_392 INVX1_392/A gnd INVX1_392/Y vdd INVX1
XINVX1_381 INVX1_381/A gnd INVX1_381/Y vdd INVX1
XNAND2X1_717 NAND2X1_717/A NAND2X1_717/B gnd NAND2X1_3/B vdd NAND2X1
XNAND2X1_706 INVX1_500/Y BUFX4_205/Y gnd NAND3X1_191/C vdd NAND2X1
XNAND2X1_728 INVX1_515/Y BUFX4_202/Y gnd NAND3X1_203/C vdd NAND2X1
XNAND2X1_739 OAI21X1_75/Y BUFX4_132/Y gnd NAND2X1_739/Y vdd NAND2X1
XINVX8_9 INVX8_9/A gnd INVX8_9/Y vdd INVX8
XDFFPOSX1_51 AOI22X1_13/A CLKBUF1_51/Y INVX1_104/A gnd vdd DFFPOSX1
XDFFPOSX1_40 INVX1_640/A CLKBUF1_43/Y INVX2_75/A gnd vdd DFFPOSX1
XDFFPOSX1_62 AOI22X1_24/A CLKBUF1_19/Y INVX1_115/A gnd vdd DFFPOSX1
XDFFPOSX1_84 INVX1_197/A CLKBUF1_55/Y OAI21X1_109/C gnd vdd DFFPOSX1
XDFFPOSX1_73 AOI22X1_35/A CLKBUF1_30/Y INVX1_126/A gnd vdd DFFPOSX1
XDFFPOSX1_95 INVX1_208/A CLKBUF1_19/Y DFFPOSX1_95/D gnd vdd DFFPOSX1
XBUFX4_18 BUFX4_22/A gnd BUFX4_18/Y vdd BUFX4
XBUFX4_29 BUFX4_27/A gnd BUFX4_29/Y vdd BUFX4
XFILL_43_5_0 gnd vdd FILL
XNAND3X1_323 BUFX4_122/Y NAND3X1_322/Y NAND3X1_323/C gnd NAND2X1_914/B vdd NAND3X1
XNAND3X1_301 BUFX4_122/Y NAND3X1_300/Y NAND3X1_301/C gnd NAND2X1_881/B vdd NAND3X1
XNAND3X1_312 INVX1_629/Y BUFX4_99/Y BUFX4_167/Y gnd NAND3X1_312/Y vdd NAND3X1
XNAND3X1_334 AOI22X1_130/Y NAND3X1_334/B AND2X2_87/Y gnd NOR2X1_432/A vdd NAND3X1
XNAND3X1_356 NOR2X1_466/Y NOR2X1_467/Y BUFX4_11/Y gnd NAND3X1_356/Y vdd NAND3X1
XNAND3X1_345 NOR2X1_466/Y INVX2_90/A NOR2X1_467/Y gnd NOR3X1_80/C vdd NAND3X1
XFILL_34_5_0 gnd vdd FILL
XFILL_22_1 gnd vdd FILL
XOAI21X1_519 BUFX4_214/Y NAND2X1_438/B NAND2X1_479/Y gnd OAI21X1_520/A vdd OAI21X1
XOAI21X1_508 AND2X2_38/Y BUFX4_128/Y INVX4_5/Y gnd OAI21X1_509/B vdd OAI21X1
XDFFPOSX1_422 BUFX2_86/A CLKBUF1_44/Y NOR3X1_29/Y gnd vdd DFFPOSX1
XDFFPOSX1_411 NOR2X1_14/A CLKBUF1_20/Y NOR3X1_19/Y gnd vdd DFFPOSX1
XDFFPOSX1_400 INVX1_460/A CLKBUF1_62/Y OAI21X1_57/Y gnd vdd DFFPOSX1
XDFFPOSX1_444 NAND3X1_14/A CLKBUF1_54/Y BUFX2_43/A gnd vdd DFFPOSX1
XDFFPOSX1_455 NAND3X1_36/A CLKBUF1_41/Y BUFX2_54/A gnd vdd DFFPOSX1
XDFFPOSX1_433 BUFX2_92/A CLKBUF1_44/Y NOR3X1_40/Y gnd vdd DFFPOSX1
XDFFPOSX1_488 BUFX2_55/A CLKBUF1_10/Y NAND3X1_39/Y gnd vdd DFFPOSX1
XDFFPOSX1_477 BUFX2_44/A CLKBUF1_33/Y NAND3X1_17/Y gnd vdd DFFPOSX1
XNAND2X1_503 INVX8_5/A OAI21X1_531/Y gnd NAND2X1_503/Y vdd NAND2X1
XDFFPOSX1_499 BUFX2_66/A CLKBUF1_6/Y NAND3X1_61/Y gnd vdd DFFPOSX1
XDFFPOSX1_466 NAND3X1_58/A CLKBUF1_36/Y BUFX2_65/A gnd vdd DFFPOSX1
XNAND2X1_514 BUFX4_214/Y MUX2X1_36/Y gnd OAI21X1_569/C vdd NAND2X1
XNAND2X1_525 AOI22X1_99/B AOI22X1_99/A gnd INVX2_64/A vdd NAND2X1
XNAND2X1_536 INVX2_36/Y INVX2_53/A gnd INVX1_401/A vdd NAND2X1
XNAND2X1_547 INVX8_4/A NAND2X1_547/B gnd NAND2X1_547/Y vdd NAND2X1
XNAND2X1_558 MUX2X1_20/S MUX2X1_49/B gnd NAND2X1_559/B vdd NAND2X1
XNAND2X1_569 OR2X2_38/B NOR2X1_335/Y gnd NAND2X1_569/Y vdd NAND2X1
XFILL_0_5_0 gnd vdd FILL
XFILL_25_5_0 gnd vdd FILL
XAOI21X1_160 AOI21X1_160/A AOI21X1_160/B INVX2_65/Y gnd NOR3X1_59/A vdd AOI21X1
XAOI21X1_182 INVX8_7/A OR2X2_29/A OAI21X1_703/Y gnd NOR3X1_62/A vdd AOI21X1
XAOI21X1_171 INVX4_7/A MUX2X1_29/Y AOI21X1_171/C gnd OAI21X1_678/C vdd AOI21X1
XAOI21X1_193 INVX2_55/A AND2X2_66/A OAI21X1_730/Y gnd NOR2X1_348/A vdd AOI21X1
XFILL_8_6_0 gnd vdd FILL
XFILL_16_5_0 gnd vdd FILL
XNAND3X1_131 NAND3X1_130/Y OAI21X1_541/Y NAND3X1_131/C gnd INVX1_77/A vdd NAND3X1
XNAND3X1_120 NAND3X1_117/Y OAI21X1_494/Y AOI21X1_90/Y gnd INVX1_73/A vdd NAND3X1
XNAND3X1_142 OAI21X1_605/Y OAI21X1_611/Y NOR3X1_57/Y gnd INVX1_83/A vdd NAND3X1
XNAND3X1_153 OAI21X1_677/Y NAND2X1_565/Y NAND3X1_153/C gnd AOI21X1_171/C vdd NAND3X1
XNAND3X1_164 OR2X2_40/Y NAND2X1_586/Y NOR2X1_347/Y gnd NOR3X1_63/C vdd NAND3X1
XNAND3X1_175 INVX8_11/Y NAND3X1_175/B NAND3X1_175/C gnd NAND3X1_178/B vdd NAND3X1
XNAND3X1_197 BUFX4_219/Y NAND3X1_197/B NAND3X1_197/C gnd NAND2X1_720/B vdd NAND3X1
XNAND3X1_186 NAND3X1_186/A NAND3X1_186/B NAND3X1_186/C gnd NOR2X1_400/A vdd NAND3X1
XOAI21X1_305 INVX1_328/Y OAI21X1_305/B AOI21X1_38/Y gnd AOI21X1_39/C vdd OAI21X1
XOAI21X1_316 INVX1_339/Y INVX4_4/A OAI21X1_316/C gnd MUX2X1_21/B vdd OAI21X1
XOAI21X1_327 NOR2X1_124/Y OAI22X1_24/C NAND2X1_297/Y gnd NOR2X1_126/A vdd OAI21X1
XOAI21X1_338 AOI21X1_45/Y AND2X2_21/Y NAND3X1_92/A gnd AOI21X1_46/C vdd OAI21X1
XOAI21X1_349 INVX1_353/Y INVX8_5/A NAND2X1_329/Y gnd NAND2X1_427/B vdd OAI21X1
XBUFX4_3 CLK gnd BUFX4_3/Y vdd BUFX4
XDFFPOSX1_230 OAI21X1_113/C CLKBUF1_21/Y INVX1_74/A gnd vdd DFFPOSX1
XDFFPOSX1_263 MUX2X1_9/A CLKBUF1_26/Y NAND3X1_24/A gnd vdd DFFPOSX1
XDFFPOSX1_252 OAI21X1_157/C CLKBUF1_21/Y INVX1_96/A gnd vdd DFFPOSX1
XDFFPOSX1_241 OAI21X1_135/C CLKBUF1_63/Y INVX1_85/A gnd vdd DFFPOSX1
XXOR2X1_16 BUFX2_91/A XOR2X1_12/B gnd XOR2X1_16/Y vdd XOR2X1
XNAND2X1_300 AOI22X1_96/B AOI22X1_96/A gnd INVX1_393/A vdd NAND2X1
XDFFPOSX1_274 AOI22X1_57/A CLKBUF1_52/Y NAND3X1_46/A gnd vdd DFFPOSX1
XDFFPOSX1_285 AOI22X1_68/A CLKBUF1_17/Y NAND3X1_68/A gnd vdd DFFPOSX1
XNAND2X1_311 NOR2X1_6/B NOR2X1_70/B gnd NOR2X1_131/A vdd NAND2X1
XDFFPOSX1_296 NOR2X1_134/B CLKBUF1_56/Y NOR3X1_1/Y gnd vdd DFFPOSX1
XNAND2X1_333 INVX8_8/A NOR2X1_249/B gnd OAI21X1_351/C vdd NAND2X1
XNAND2X1_322 INVX4_4/A INVX1_351/Y gnd AOI21X1_48/A vdd NAND2X1
XNAND2X1_344 AND2X2_93/B INVX2_49/Y gnd INVX1_356/A vdd NAND2X1
XNAND2X1_377 INVX8_7/A NOR2X1_311/B gnd NAND2X1_377/Y vdd NAND2X1
XNAND2X1_366 AND2X2_70/B OAI21X1_379/Y gnd NAND2X1_366/Y vdd NAND2X1
XNAND2X1_355 AND2X2_93/B INVX2_49/A gnd INVX2_56/A vdd NAND2X1
XNAND2X1_388 BUFX4_229/Y INVX1_368/Y gnd NAND2X1_388/Y vdd NAND2X1
XNAND2X1_399 BUFX4_85/Y NOR2X1_207/B gnd NAND2X1_399/Y vdd NAND2X1
XNOR3X1_51 INVX1_247/Y AOI21X1_4/C NOR3X1_49/C gnd NOR3X1_51/Y vdd NOR3X1
XNOR3X1_62 NOR3X1_62/A NOR3X1_62/B AND2X2_63/Y gnd NOR3X1_62/Y vdd NOR3X1
XNOR3X1_40 NOR3X1_4/A INVX1_181/Y NOR3X1_4/C gnd NOR3X1_40/Y vdd NOR3X1
XNOR3X1_73 NOR3X1_80/A NOR3X1_73/B NOR3X1_78/C gnd NOR3X1_73/Y vdd NOR3X1
XFILL_40_3_0 gnd vdd FILL
XINVX4_3 INVX4_3/A gnd INVX4_3/Y vdd INVX4
XOAI21X1_850 OR2X2_48/A INVX1_483/Y INVX1_484/Y gnd OAI21X1_851/C vdd OAI21X1
XOAI21X1_872 INVX2_74/Y DFFPOSX1_43/Q DFFPOSX1_45/Q gnd NOR2X1_404/A vdd OAI21X1
XOAI21X1_861 OAI21X1_860/Y AOI21X1_220/Y OAI21X1_861/C gnd OAI21X1_861/Y vdd OAI21X1
XOAI21X1_883 INVX1_654/Y OAI21X1_887/B INVX4_11/Y gnd OAI21X1_883/Y vdd OAI21X1
XOAI21X1_894 INVX8_14/Y AOI21X1_231/Y OAI21X1_894/C gnd OAI21X1_894/Y vdd OAI21X1
XFILL_31_3_0 gnd vdd FILL
XNAND3X1_6 INVX4_1/Y INVX1_150/Y NAND3X1_7/C gnd NAND3X1_6/Y vdd NAND3X1
XFILL_39_4_0 gnd vdd FILL
XFILL_22_3_0 gnd vdd FILL
XOAI21X1_102 BUFX4_182/Y INVX1_101/Y OAI21X1_102/C gnd INVX1_581/A vdd OAI21X1
XOAI21X1_113 BUFX4_272/Y BUFX4_195/Y OAI21X1_113/C gnd OAI21X1_113/Y vdd OAI21X1
XOAI21X1_146 BUFX4_182/Y INVX1_123/Y OAI21X1_145/Y gnd INVX1_625/A vdd OAI21X1
XOAI21X1_124 BUFX4_182/Y INVX1_112/Y OAI21X1_123/Y gnd INVX1_603/A vdd OAI21X1
XOAI21X1_135 BUFX4_269/Y BUFX4_192/Y OAI21X1_135/C gnd OAI21X1_135/Y vdd OAI21X1
XOAI21X1_179 BUFX4_12/Y BUFX4_199/Y OAI21X1_845/Y gnd NAND3X1_43/C vdd OAI21X1
XOAI21X1_168 BUFX4_14/Y BUFX4_197/Y OAI21X1_168/C gnd NAND3X1_21/C vdd OAI21X1
XOAI21X1_157 BUFX4_273/Y BUFX4_193/Y OAI21X1_157/C gnd OAI21X1_157/Y vdd OAI21X1
XNAND2X1_152 AOI21X1_24/A INVX1_259/Y gnd NOR2X1_43/B vdd NAND2X1
XNAND2X1_141 OAI21X1_244/Y NAND2X1_140/Y gnd NOR2X1_33/B vdd NAND2X1
XNAND2X1_130 NAND3X1_80/Y NAND2X1_130/B gnd NOR2X1_29/B vdd NAND2X1
XFILL_5_4_0 gnd vdd FILL
XNAND2X1_163 INVX1_268/A NAND2X1_163/B gnd NAND2X1_163/Y vdd NAND2X1
XNAND2X1_174 INVX1_276/Y INVX1_275/A gnd NAND2X1_175/A vdd NAND2X1
XNAND2X1_196 INVX4_4/A AOI22X1_63/A gnd NAND2X1_196/Y vdd NAND2X1
XNAND2X1_185 INVX1_285/Y NOR2X1_56/B gnd NAND2X1_186/A vdd NAND2X1
XFILL_13_3_0 gnd vdd FILL
XAOI22X1_19 AOI22X1_19/A AOI22X1_9/B OR2X2_3/A AOI22X1_19/D gnd AOI22X1_19/Y vdd AOI22X1
XOAI21X1_680 NOR2X1_325/B NOR2X1_325/A INVX1_413/Y gnd AND2X2_58/A vdd OAI21X1
XOAI21X1_691 AND2X2_58/Y NOR2X1_333/Y AOI21X1_38/B gnd NAND3X1_156/B vdd OAI21X1
XINVX1_711 INVX1_711/A gnd INVX1_711/Y vdd INVX1
XINVX1_700 INVX1_700/A gnd INVX1_700/Y vdd INVX1
XNOR3X1_9 NOR3X1_9/A NOR3X1_9/B NOR3X1_9/C gnd NOR3X1_9/Y vdd NOR3X1
XINVX1_722 INVX1_722/A gnd INVX1_722/Y vdd INVX1
XINVX1_733 INVX1_733/A gnd INVX1_733/Y vdd INVX1
XINVX1_744 data_memory_interface_data[20] gnd INVX1_744/Y vdd INVX1
XINVX1_755 data_memory_interface_data[15] gnd INVX1_755/Y vdd INVX1
XFILL_5_3 gnd vdd FILL
XXNOR2X1_30 XNOR2X1_30/A NOR2X1_46/B gnd XNOR2X1_30/Y vdd XNOR2X1
XXNOR2X1_41 XNOR2X1_41/A NOR2X1_45/B gnd XNOR2X1_41/Y vdd XNOR2X1
XXNOR2X1_52 NOR3X1_66/Y BUFX2_65/A gnd XNOR2X1_52/Y vdd XNOR2X1
XBUFX2_51 BUFX2_51/A gnd instruction_memory_interface_address[12] vdd BUFX2
XBUFX2_62 BUFX2_62/A gnd instruction_memory_interface_address[23] vdd BUFX2
XBUFX2_40 BUFX2_40/A gnd instruction_memory_interface_address[1] vdd BUFX2
XBUFX2_73 vdd gnd instruction_memory_interface_frame_mask[1] vdd BUFX2
XBUFX2_84 BUFX2_84/A gnd BUFX2_84/Y vdd BUFX2
XBUFX2_95 BUFX2_95/A gnd BUFX2_95/Y vdd BUFX2
XAOI21X1_52 INVX8_3/A AOI21X1_52/B INVX8_7/A gnd AOI21X1_52/Y vdd AOI21X1
XAOI21X1_41 NAND3X1_91/C AOI21X1_41/B AOI21X1_41/C gnd AOI21X1_41/Y vdd AOI21X1
XAOI21X1_30 AOI21X1_30/A XNOR2X1_46/A NOR2X1_55/Y gnd XOR2X1_7/A vdd AOI21X1
XAOI21X1_74 AOI21X1_74/A NOR2X1_210/B AOI21X1_74/C gnd AOI21X1_74/Y vdd AOI21X1
XAOI21X1_85 AOI21X1_85/A AOI21X1_85/B BUFX4_77/Y gnd OAI22X1_17/B vdd AOI21X1
XAOI21X1_63 AOI21X1_63/A NOR2X1_195/A AOI21X1_63/C gnd AOI21X1_63/Y vdd AOI21X1
XAOI21X1_96 AOI21X1_96/A AOI21X1_96/B AOI21X1_96/C gnd AOI21X1_96/Y vdd AOI21X1
XOAI21X1_3 INVX1_3/Y BUFX4_21/Y OAI21X1_3/C gnd OAI21X1_3/Y vdd OAI21X1
XNOR2X1_409 XOR2X1_16/Y XOR2X1_17/Y gnd NOR2X1_409/Y vdd NOR2X1
XOAI22X1_60 INVX2_92/Y INVX4_14/Y OAI22X1_60/C OAI22X1_60/D gnd OAI22X1_60/Y vdd OAI22X1
XINVX1_541 INVX1_614/A gnd INVX1_541/Y vdd INVX1
XINVX1_563 INVX1_636/A gnd INVX1_563/Y vdd INVX1
XINVX1_552 INVX1_625/A gnd INVX1_552/Y vdd INVX1
XINVX1_530 INVX1_603/A gnd INVX1_530/Y vdd INVX1
XINVX1_585 INVX1_585/A gnd INVX1_585/Y vdd INVX1
XINVX1_596 INVX1_523/A gnd INVX1_596/Y vdd INVX1
XINVX1_574 INVX1_501/A gnd INVX1_574/Y vdd INVX1
XFILL_37_7_1 gnd vdd FILL
XFILL_36_2_0 gnd vdd FILL
XFILL_20_6_1 gnd vdd FILL
XFILL_3_7_1 gnd vdd FILL
XXOR2X1_6 XOR2X1_6/A XOR2X1_6/B gnd XOR2X1_6/Y vdd XOR2X1
XFILL_28_7_1 gnd vdd FILL
XFILL_2_2_0 gnd vdd FILL
XFILL_27_2_0 gnd vdd FILL
XMUX2X1_7 MUX2X1_7/A MUX2X1_7/B INVX4_4/A gnd MUX2X1_7/Y vdd MUX2X1
XFILL_11_6_1 gnd vdd FILL
XFILL_10_1_0 gnd vdd FILL
XCLKBUF1_8 BUFX4_2/Y gnd CLKBUF1_8/Y vdd CLKBUF1
XAOI22X1_140 data_memory_interface_data[3] BUFX4_105/Y AOI22X1_140/C BUFX4_8/Y gnd
+ AOI22X1_140/Y vdd AOI22X1
XAOI22X1_151 data_memory_interface_data[15] BUFX4_109/Y BUFX4_169/Y BUFX4_10/Y gnd
+ AOI22X1_151/Y vdd AOI22X1
XBUFX4_102 BUFX4_99/A gnd BUFX4_102/Y vdd BUFX4
XAOI22X1_162 data_memory_interface_data[26] BUFX4_109/Y BUFX4_171/Y BUFX4_251/Y gnd
+ AOI22X1_162/Y vdd AOI22X1
XBUFX4_113 NOR2X1_7/Y gnd INVX8_2/A vdd BUFX4
XBUFX4_124 INVX8_7/Y gnd BUFX4_124/Y vdd BUFX4
XBUFX4_146 BUFX4_148/A gnd BUFX4_146/Y vdd BUFX4
XFILL_19_7_1 gnd vdd FILL
XBUFX4_135 AND2X2_79/Y gnd BUFX4_135/Y vdd BUFX4
XNOR2X1_206 BUFX4_58/Y AND2X2_29/A gnd NOR2X1_206/Y vdd NOR2X1
XFILL_18_2_0 gnd vdd FILL
XBUFX4_179 BUFX4_178/A gnd BUFX4_179/Y vdd BUFX4
XBUFX4_157 NOR2X1_2/Y gnd BUFX4_157/Y vdd BUFX4
XBUFX4_168 BUFX4_164/A gnd BUFX4_168/Y vdd BUFX4
XNOR2X1_228 INVX2_57/Y NOR2X1_228/B gnd NOR2X1_228/Y vdd NOR2X1
XNOR2X1_239 BUFX4_57/Y NOR2X1_239/B gnd NOR2X1_239/Y vdd NOR2X1
XNOR2X1_217 INVX8_9/A OR2X2_27/B gnd NOR2X1_217/Y vdd NOR2X1
XOAI21X1_1003 INVX4_13/Y INVX8_16/Y data_memory_interface_data[30] gnd OAI21X1_1003/Y
+ vdd OAI21X1
XOAI21X1_1025 NOR2X1_481/Y INVX4_12/A data_memory_interface_data[28] gnd OAI21X1_1025/Y
+ vdd OAI21X1
XOAI21X1_1036 BUFX4_64/Y BUFX4_68/Y AOI22X1_152/Y gnd OAI21X1_1036/Y vdd OAI21X1
XOAI21X1_1014 OAI21X1_993/B data_memory_interface_data[24] BUFX4_10/Y gnd AOI21X1_267/C
+ vdd OAI21X1
XOAI21X1_1058 AOI21X1_270/Y OAI21X1_1057/Y INVX1_756/Y gnd OAI21X1_1058/Y vdd OAI21X1
XOAI21X1_1047 BUFX4_67/Y BUFX4_70/Y AOI22X1_163/Y gnd OAI21X1_1047/Y vdd OAI21X1
XOAI21X1_1069 AOI21X1_271/Y OAI21X1_1069/B NOR2X1_487/Y gnd OAI21X1_1069/Y vdd OAI21X1
XINVX1_371 INVX1_371/A gnd INVX1_371/Y vdd INVX1
XINVX1_360 OR2X2_29/B gnd INVX1_360/Y vdd INVX1
XINVX1_393 INVX1_393/A gnd INVX1_393/Y vdd INVX1
XINVX1_382 INVX1_382/A gnd INVX1_382/Y vdd INVX1
XNAND2X1_718 OAI21X1_68/Y BUFX4_133/Y gnd NAND2X1_718/Y vdd NAND2X1
XNAND2X1_707 INVX1_501/A INVX2_73/Y gnd NAND3X1_189/A vdd NAND2X1
XNAND2X1_729 NAND2X1_727/Y NAND2X1_729/B gnd NAND2X1_7/B vdd NAND2X1
XDFFPOSX1_41 DFFPOSX1_41/Q CLKBUF1_43/Y INVX1_501/A gnd vdd DFFPOSX1
XDFFPOSX1_30 AOI22X1_30/D CLKBUF1_32/Y DFFPOSX1_30/D gnd vdd DFFPOSX1
XDFFPOSX1_52 AOI22X1_14/A CLKBUF1_55/Y INVX1_105/A gnd vdd DFFPOSX1
XDFFPOSX1_63 AOI22X1_25/A CLKBUF1_19/Y INVX1_116/A gnd vdd DFFPOSX1
XDFFPOSX1_85 INVX1_198/A CLKBUF1_11/Y OAI21X1_111/C gnd vdd DFFPOSX1
XDFFPOSX1_96 INVX1_209/A CLKBUF1_30/Y OAI21X1_133/C gnd vdd DFFPOSX1
XDFFPOSX1_74 AOI22X1_36/A CLKBUF1_61/Y INVX1_127/A gnd vdd DFFPOSX1
XBUFX4_19 BUFX4_22/A gnd BUFX4_19/Y vdd BUFX4
XFILL_43_5_1 gnd vdd FILL
XNAND3X1_324 NOR2X1_409/Y NOR2X1_410/Y NAND3X1_324/C gnd NAND3X1_325/B vdd NAND3X1
XFILL_42_0_0 gnd vdd FILL
XNAND3X1_313 BUFX4_123/Y NAND3X1_312/Y NAND3X1_313/C gnd NAND2X1_899/B vdd NAND3X1
XNAND3X1_302 INVX1_619/Y BUFX4_100/Y BUFX4_165/Y gnd NAND3X1_302/Y vdd NAND3X1
XNAND3X1_335 AND2X2_95/A AND2X2_95/B AOI22X1_131/Y gnd OR2X2_68/A vdd NAND3X1
XNAND3X1_346 INVX4_12/Y INVX2_87/Y INVX4_13/A gnd OAI22X1_58/C vdd NAND3X1
XNAND3X1_357 data_memory_interface_data[14] NOR2X1_477/Y INVX4_13/A gnd NAND3X1_357/Y
+ vdd NAND3X1
XFILL_34_5_1 gnd vdd FILL
XFILL_22_2 gnd vdd FILL
XFILL_33_0_0 gnd vdd FILL
XOAI21X1_509 NOR2X1_241/Y OAI21X1_509/B AOI21X1_94/Y gnd AOI21X1_95/C vdd OAI21X1
XFILL_15_1 gnd vdd FILL
XDFFPOSX1_401 INVX2_81/A CLKBUF1_37/Y OAI21X1_58/Y gnd vdd DFFPOSX1
XDFFPOSX1_412 INVX1_228/A CLKBUF1_20/Y NAND3X1_72/Y gnd vdd DFFPOSX1
XDFFPOSX1_456 NAND3X1_38/A CLKBUF1_35/Y BUFX2_55/A gnd vdd DFFPOSX1
XDFFPOSX1_445 NAND3X1_16/A CLKBUF1_33/Y BUFX2_44/A gnd vdd DFFPOSX1
XDFFPOSX1_434 BUFX2_93/A CLKBUF1_13/Y NOR3X1_41/Y gnd vdd DFFPOSX1
XDFFPOSX1_423 INVX1_495/A CLKBUF1_59/Y NOR3X1_30/Y gnd vdd DFFPOSX1
XDFFPOSX1_489 BUFX2_56/A CLKBUF1_10/Y NAND3X1_41/Y gnd vdd DFFPOSX1
XDFFPOSX1_478 INVX2_72/A CLKBUF1_10/Y NAND3X1_19/Y gnd vdd DFFPOSX1
XDFFPOSX1_467 NAND3X1_60/A CLKBUF1_6/Y BUFX2_66/A gnd vdd DFFPOSX1
XINVX1_190 NOR2X1_11/A gnd INVX1_190/Y vdd INVX1
XNAND2X1_515 BUFX4_52/Y NAND2X1_561/B gnd OAI21X1_570/C vdd NAND2X1
XNAND2X1_526 INVX8_5/A MUX2X1_36/A gnd NAND2X1_526/Y vdd NAND2X1
XNAND2X1_504 BUFX4_56/Y NOR2X1_323/B gnd NAND2X1_505/B vdd NAND2X1
XNAND2X1_548 INVX8_5/A MUX2X1_41/Y gnd NAND2X1_548/Y vdd NAND2X1
XNAND2X1_537 MUX2X1_40/S MUX2X1_41/Y gnd NAND2X1_537/Y vdd NAND2X1
XNAND2X1_559 NAND2X1_556/Y NAND2X1_559/B gnd NOR2X1_328/B vdd NAND2X1
XFILL_0_5_1 gnd vdd FILL
XFILL_25_5_1 gnd vdd FILL
XFILL_24_0_0 gnd vdd FILL
XAOI21X1_150 AOI21X1_150/A NAND2X1_543/Y OAI22X1_30/C gnd NOR3X1_58/C vdd AOI21X1
XAOI21X1_172 INVX8_3/A MUX2X1_38/A INVX8_7/A gnd OAI21X1_686/C vdd AOI21X1
XAOI21X1_161 INVX8_3/A NOR2X1_323/B INVX8_7/A gnd OAI21X1_652/C vdd AOI21X1
XAOI21X1_183 INVX1_416/Y INVX8_12/A OAI21X1_707/Y gnd NAND3X1_158/B vdd AOI21X1
XAOI21X1_194 NAND2X1_318/Y INVX1_419/A NOR2X1_349/Y gnd OAI21X1_750/B vdd AOI21X1
XFILL_8_6_1 gnd vdd FILL
XFILL_7_1_0 gnd vdd FILL
XFILL_16_5_1 gnd vdd FILL
XFILL_15_0_0 gnd vdd FILL
XNAND3X1_132 BUFX4_91/Y NOR2X1_281/B OR2X2_32/Y gnd NAND3X1_132/Y vdd NAND3X1
XNAND3X1_121 NAND3X1_121/A OR2X2_29/Y NAND3X1_121/C gnd AOI22X1_90/C vdd NAND3X1
XNAND3X1_110 NAND3X1_110/A NAND3X1_110/B AOI21X1_66/Y gnd INVX1_68/A vdd NAND3X1
XNAND3X1_143 NAND3X1_143/A NAND2X1_544/Y OAI21X1_625/Y gnd NAND3X1_143/Y vdd NAND3X1
XNAND3X1_154 NAND3X1_154/A OAI21X1_681/Y NOR3X1_60/Y gnd INVX1_88/A vdd NAND3X1
XNAND3X1_165 NAND3X1_165/A NAND3X1_165/B NOR3X1_63/Y gnd INVX1_92/A vdd NAND3X1
XNAND3X1_176 INVX2_26/A INVX1_434/Y NAND2X1_602/Y gnd NAND3X1_177/B vdd NAND3X1
XNAND3X1_198 INVX1_512/Y BUFX4_209/Y BUFX4_34/Y gnd NAND3X1_199/B vdd NAND3X1
XNAND3X1_187 NAND3X1_187/A NAND3X1_187/B AOI21X1_222/Y gnd NOR2X1_400/B vdd NAND3X1
XOAI21X1_328 INVX1_393/A AOI22X1_96/C AOI22X1_96/B gnd OAI21X1_329/B vdd OAI21X1
XOAI21X1_306 INVX1_329/Y NOR2X1_103/Y INVX2_67/A gnd OR2X2_39/A vdd OAI21X1
XOAI21X1_317 INVX1_340/Y INVX4_4/A NAND2X1_272/Y gnd MUX2X1_21/A vdd OAI21X1
XOAI21X1_339 INVX8_8/A MUX2X1_13/Y NOR2X1_152/Y gnd NOR2X1_153/A vdd OAI21X1
XDFFPOSX1_231 OAI21X1_115/C CLKBUF1_4/Y INVX1_75/A gnd vdd DFFPOSX1
XDFFPOSX1_220 AOI22X1_170/C CLKBUF1_28/Y INVX1_666/A gnd vdd DFFPOSX1
XBUFX4_4 CLK gnd BUFX4_4/Y vdd BUFX4
XDFFPOSX1_264 MUX2X1_8/A CLKBUF1_26/Y NAND3X1_26/A gnd vdd DFFPOSX1
XDFFPOSX1_253 OAI21X1_159/C CLKBUF1_23/Y INVX1_97/A gnd vdd DFFPOSX1
XDFFPOSX1_242 DFFPOSX1_98/D CLKBUF1_3/Y INVX1_86/A gnd vdd DFFPOSX1
XXOR2X1_17 OR2X2_52/B XOR2X1_13/B gnd XOR2X1_17/Y vdd XOR2X1
XNAND2X1_301 INVX2_43/A MUX2X1_8/Y gnd AOI22X1_96/C vdd NAND2X1
XDFFPOSX1_275 AOI22X1_58/A CLKBUF1_52/Y NAND3X1_48/A gnd vdd DFFPOSX1
XDFFPOSX1_297 NOR2X1_134/A CLKBUF1_56/Y NOR3X1_2/Y gnd vdd DFFPOSX1
XDFFPOSX1_286 AND2X2_1/B CLKBUF1_34/Y NAND3X1_5/Y gnd vdd DFFPOSX1
XNAND2X1_323 INVX8_8/A MUX2X1_21/A gnd AOI21X1_50/A vdd NAND2X1
XNAND2X1_345 AND2X2_23/Y AOI21X1_49/B gnd NOR2X1_203/B vdd NAND2X1
XNAND2X1_312 NOR2X1_129/Y NOR2X1_128/Y gnd INVX1_358/A vdd NAND2X1
XNAND2X1_334 BUFX4_40/Y INVX2_21/A gnd NAND2X1_334/Y vdd NAND2X1
XNAND2X1_378 INVX8_8/A MUX2X1_21/B gnd OAI21X1_392/C vdd NAND2X1
XNAND2X1_356 INVX8_8/A MUX2X1_13/Y gnd NOR2X1_195/A vdd NAND2X1
XNAND2X1_367 INVX8_4/A NOR2X1_223/B gnd OAI21X1_383/C vdd NAND2X1
XNAND2X1_389 INVX8_4/A OAI21X1_474/A gnd NAND2X1_389/Y vdd NAND2X1
XNOR3X1_52 INVX1_251/Y AOI21X1_4/C NOR3X1_49/C gnd NOR3X1_52/Y vdd NOR3X1
XNOR3X1_41 NOR3X1_3/A INVX1_182/Y BUFX4_49/Y gnd NOR3X1_41/Y vdd NOR3X1
XNOR3X1_30 NOR3X1_35/A INVX1_171/Y NOR3X1_8/C gnd NOR3X1_30/Y vdd NOR3X1
XNOR3X1_63 AND2X2_68/Y NOR3X1_63/B NOR3X1_63/C gnd NOR3X1_63/Y vdd NOR3X1
XNOR3X1_74 NOR3X1_78/C NOR3X1_73/B NOR3X1_79/A gnd NOR3X1_74/Y vdd NOR3X1
XFILL_40_3_1 gnd vdd FILL
XINVX4_4 INVX4_4/A gnd INVX4_4/Y vdd INVX4
XOAI21X1_840 NOR2X1_388/Y OAI21X1_839/Y OAI21X1_840/C gnd OAI21X1_840/Y vdd OAI21X1
XOAI21X1_851 OR2X2_48/A OR2X2_48/B OAI21X1_851/C gnd OAI21X1_851/Y vdd OAI21X1
XOAI21X1_862 XNOR2X1_53/Y NOR3X1_4/A OAI21X1_862/C gnd OAI21X1_862/Y vdd OAI21X1
XOAI21X1_884 INVX1_655/Y OAI21X1_887/B INVX4_11/Y gnd OAI21X1_884/Y vdd OAI21X1
XOAI21X1_873 INVX2_77/Y INVX1_502/A INVX1_504/A gnd NOR2X1_407/A vdd OAI21X1
XOAI21X1_895 INVX8_14/Y AOI21X1_231/Y AOI22X1_119/Y gnd OAI21X1_895/Y vdd OAI21X1
XNAND2X1_890 NAND2X1_890/A NAND2X1_890/B gnd NAND2X1_56/B vdd NAND2X1
XFILL_31_3_1 gnd vdd FILL
XNAND3X1_7 INVX4_1/Y INVX1_153/Y NAND3X1_7/C gnd NAND3X1_7/Y vdd NAND3X1
XFILL_39_4_1 gnd vdd FILL
XFILL_22_3_1 gnd vdd FILL
XOAI21X1_103 BUFX4_270/Y BUFX4_192/Y DFFPOSX1_81/D gnd OAI21X1_104/C vdd OAI21X1
XOAI21X1_147 BUFX4_272/Y BUFX4_195/Y OAI21X1_147/C gnd OAI21X1_147/Y vdd OAI21X1
XOAI21X1_114 BUFX4_183/Y INVX1_107/Y OAI21X1_113/Y gnd INVX1_593/A vdd OAI21X1
XOAI21X1_125 BUFX4_269/Y BUFX4_192/Y DFFPOSX1_92/D gnd OAI21X1_125/Y vdd OAI21X1
XOAI21X1_136 BUFX4_184/Y INVX1_118/Y OAI21X1_135/Y gnd INVX1_542/A vdd OAI21X1
XOAI21X1_169 BUFX4_14/Y BUFX4_197/Y OAI21X1_169/C gnd NAND3X1_23/C vdd OAI21X1
XOAI21X1_158 BUFX4_182/Y INVX1_129/Y OAI21X1_157/Y gnd INVX1_637/A vdd OAI21X1
XBUFX2_1 gnd gnd data_memory_interface_address[0] vdd BUFX2
XNAND2X1_142 NAND2X1_140/Y NAND2X1_142/B gnd NAND2X1_142/Y vdd NAND2X1
XNAND2X1_153 INVX1_261/A INVX1_260/Y gnd NAND2X1_153/Y vdd NAND2X1
XNAND2X1_131 NAND3X1_80/Y NAND2X1_131/B gnd INVX1_244/A vdd NAND2X1
XNAND2X1_120 INVX2_5/Y OR2X2_9/A gnd AOI21X1_6/B vdd NAND2X1
XFILL_5_4_1 gnd vdd FILL
XNAND2X1_175 NAND2X1_175/A AND2X2_16/B gnd NOR2X1_49/B vdd NAND2X1
XNAND2X1_164 MUX2X1_1/A BUFX4_232/Y gnd NAND3X1_84/B vdd NAND2X1
XNAND2X1_186 NAND2X1_186/A INVX1_286/Y gnd XOR2X1_7/B vdd NAND2X1
XNAND2X1_197 INVX4_4/A AOI22X1_64/A gnd NAND2X1_197/Y vdd NAND2X1
XFILL_13_3_1 gnd vdd FILL
XINVX2_1 INVX2_1/A gnd INVX2_1/Y vdd INVX2
XAOI21X1_1 AOI21X1_1/A AOI21X1_1/B reset gnd AOI21X1_1/Y vdd AOI21X1
XOAI21X1_692 AOI21X1_38/A NOR2X1_333/Y OR2X2_38/B gnd NOR2X1_336/B vdd OAI21X1
XOAI21X1_681 INVX2_70/A AND2X2_58/A NOR2X1_331/Y gnd OAI21X1_681/Y vdd OAI21X1
XOAI21X1_670 INVX2_70/Y AOI21X1_168/B OAI21X1_670/C gnd NAND3X1_154/A vdd OAI21X1
XINVX1_701 OR2X2_56/A gnd INVX1_701/Y vdd INVX1
XINVX1_712 INVX1_712/A gnd INVX1_712/Y vdd INVX1
XINVX1_723 INVX1_723/A gnd INVX1_723/Y vdd INVX1
XINVX1_745 data_memory_interface_data[11] gnd INVX1_745/Y vdd INVX1
XINVX1_734 data_memory_interface_data[16] gnd INVX1_734/Y vdd INVX1
XINVX1_756 INVX1_756/A gnd INVX1_756/Y vdd INVX1
XXNOR2X1_20 AOI21X1_15/Y INVX1_253/A gnd XNOR2X1_20/Y vdd XNOR2X1
XXNOR2X1_31 NOR2X1_37/B INVX2_12/Y gnd NOR2X1_47/A vdd XNOR2X1
XXNOR2X1_42 XNOR2X1_42/A NOR2X1_49/B gnd XNOR2X1_42/Y vdd XNOR2X1
XXNOR2X1_53 NOR3X1_67/Y BUFX2_67/A gnd XNOR2X1_53/Y vdd XNOR2X1
XBUFX2_41 BUFX2_41/A gnd instruction_memory_interface_address[2] vdd BUFX2
XBUFX2_52 BUFX2_52/A gnd instruction_memory_interface_address[13] vdd BUFX2
XBUFX2_63 BUFX2_63/A gnd instruction_memory_interface_address[24] vdd BUFX2
XBUFX2_30 BUFX2_30/A gnd data_memory_interface_address[29] vdd BUFX2
XBUFX2_74 vdd gnd instruction_memory_interface_frame_mask[2] vdd BUFX2
XBUFX2_85 BUFX2_85/A gnd BUFX2_85/Y vdd BUFX2
XBUFX2_96 BUFX2_96/A gnd BUFX2_96/Y vdd BUFX2
XAOI21X1_20 MUX2X1_6/B BUFX4_150/Y NOR3X1_54/Y gnd AOI21X1_20/Y vdd AOI21X1
XAOI21X1_42 AOI22X1_70/Y AOI21X1_42/B AOI21X1_42/C gnd AOI21X1_42/Y vdd AOI21X1
XAOI21X1_31 NOR2X1_57/Y INVX1_281/A AOI21X1_31/C gnd INVX1_293/A vdd AOI21X1
XAOI21X1_53 BUFX4_38/Y INVX2_17/A AOI21X1_53/C gnd AOI21X1_53/Y vdd AOI21X1
XAOI21X1_64 AOI21X1_64/A AOI21X1_63/Y BUFX4_87/Y gnd AOI21X1_64/Y vdd AOI21X1
XAOI21X1_75 INVX4_7/A AOI21X1_75/B AOI21X1_75/C gnd AOI21X1_75/Y vdd AOI21X1
XAOI21X1_86 AOI21X1_86/A NOR2X1_150/Y NOR2X1_148/Y gnd AOI21X1_86/Y vdd AOI21X1
XAOI21X1_97 AOI21X1_97/A AOI22X1_79/D AOI22X1_80/A gnd AOI21X1_97/Y vdd AOI21X1
XOAI21X1_4 INVX1_4/Y BUFX4_18/Y OAI21X1_4/C gnd OAI21X1_4/Y vdd OAI21X1
XOAI22X1_50 AND2X2_84/Y NOR2X1_426/Y AND2X2_85/Y INVX1_697/A gnd NOR3X1_70/B vdd OAI22X1
XINVX1_520 INVX1_593/A gnd INVX1_520/Y vdd INVX1
XINVX1_553 INVX1_553/A gnd INVX1_553/Y vdd INVX1
XINVX1_531 INVX1_604/A gnd INVX1_531/Y vdd INVX1
XINVX1_542 INVX1_542/A gnd INVX1_542/Y vdd INVX1
XINVX1_564 INVX1_637/A gnd INVX1_564/Y vdd INVX1
XINVX1_575 INVX1_502/A gnd INVX1_575/Y vdd INVX1
XINVX1_586 INVX1_513/A gnd INVX1_586/Y vdd INVX1
XFILL_3_1 gnd vdd FILL
XINVX1_597 INVX1_524/A gnd INVX1_597/Y vdd INVX1
XFILL_36_2_1 gnd vdd FILL
XXOR2X1_7 XOR2X1_7/A XOR2X1_7/B gnd XOR2X1_7/Y vdd XOR2X1
XFILL_2_2_1 gnd vdd FILL
XFILL_27_2_1 gnd vdd FILL
XMUX2X1_8 MUX2X1_8/A OR2X2_59/A INVX4_4/A gnd MUX2X1_8/Y vdd MUX2X1
XFILL_10_1_1 gnd vdd FILL
XCLKBUF1_9 BUFX4_1/Y gnd CLKBUF1_9/Y vdd CLKBUF1
XAOI22X1_130 OR2X2_58/Y AOI22X1_130/B NAND2X1_951/Y OR2X2_59/Y gnd AOI22X1_130/Y vdd
+ AOI22X1
XBUFX4_103 BUFX4_99/A gnd BUFX4_103/Y vdd BUFX4
XAOI22X1_152 data_memory_interface_data[16] INVX4_14/A BUFX4_169/Y BUFX4_253/Y gnd
+ AOI22X1_152/Y vdd AOI22X1
XAOI22X1_163 data_memory_interface_data[27] BUFX4_109/Y BUFX4_171/Y BUFX4_251/Y gnd
+ AOI22X1_163/Y vdd AOI22X1
XAOI22X1_141 data_memory_interface_data[4] BUFX4_107/Y AOI22X1_141/C BUFX4_10/Y gnd
+ OAI21X1_998/C vdd AOI22X1
XBUFX4_125 INVX8_7/Y gnd BUFX4_125/Y vdd BUFX4
XBUFX4_136 OAI22X1_1/Y gnd BUFX4_136/Y vdd BUFX4
XBUFX4_114 NOR2X1_7/Y gnd BUFX4_114/Y vdd BUFX4
XBUFX4_147 BUFX4_148/A gnd BUFX4_147/Y vdd BUFX4
XNOR2X1_207 BUFX4_124/Y NOR2X1_207/B gnd NOR2X1_207/Y vdd NOR2X1
XFILL_18_2_1 gnd vdd FILL
XBUFX4_158 NOR2X1_2/Y gnd BUFX4_158/Y vdd BUFX4
XBUFX4_169 BUFX4_171/A gnd BUFX4_169/Y vdd BUFX4
XNOR2X1_229 INVX8_9/A NOR2X1_229/B gnd NOR2X1_229/Y vdd NOR2X1
XNOR2X1_218 INVX8_4/A MUX2X1_19/Y gnd NOR2X1_218/Y vdd NOR2X1
XOAI21X1_1004 INVX1_750/Y OAI21X1_992/B OAI21X1_1003/Y gnd AOI21X1_264/B vdd OAI21X1
XOAI21X1_1026 INVX1_748/Y INVX2_93/A OAI21X1_1025/Y gnd AOI22X1_148/C vdd OAI21X1
XOAI21X1_1015 BUFX4_64/Y BUFX4_68/Y NOR2X1_485/Y gnd OAI21X1_1015/Y vdd OAI21X1
XOAI21X1_1037 BUFX4_66/Y BUFX4_71/Y AOI22X1_153/Y gnd OAI21X1_1037/Y vdd OAI21X1
XOAI21X1_1059 NOR3X1_73/B INVX2_88/A INVX8_17/Y gnd INVX1_757/A vdd OAI21X1
XOAI21X1_1048 BUFX4_65/Y BUFX4_69/Y AOI22X1_164/Y gnd OAI21X1_1048/Y vdd OAI21X1
XINVX1_350 INVX1_350/A gnd INVX1_350/Y vdd INVX1
XINVX1_361 INVX1_361/A gnd INVX1_361/Y vdd INVX1
XINVX1_383 INVX1_383/A gnd INVX1_383/Y vdd INVX1
XINVX1_372 INVX1_372/A gnd INVX1_372/Y vdd INVX1
XINVX1_394 INVX1_394/A gnd INVX1_394/Y vdd INVX1
XNAND2X1_719 INVX1_509/Y BUFX4_202/Y gnd NAND3X1_197/C vdd NAND2X1
XNAND2X1_708 INVX1_495/A INVX2_75/Y gnd NAND2X1_708/Y vdd NAND2X1
XDFFPOSX1_20 AOI22X1_20/D CLKBUF1_12/Y DFFPOSX1_20/D gnd vdd DFFPOSX1
XNAND2X1_1020 data_memory_interface_data[14] INVX2_93/Y gnd NAND2X1_1020/Y vdd NAND2X1
XDFFPOSX1_42 XOR2X1_13/B CLKBUF1_39/Y OR2X2_50/A gnd vdd DFFPOSX1
XDFFPOSX1_31 AOI22X1_31/D CLKBUF1_49/Y DFFPOSX1_31/D gnd vdd DFFPOSX1
XDFFPOSX1_53 AOI22X1_15/A CLKBUF1_30/Y INVX1_106/A gnd vdd DFFPOSX1
XDFFPOSX1_86 INVX1_199/A CLKBUF1_15/Y OAI21X1_113/C gnd vdd DFFPOSX1
XDFFPOSX1_64 AOI22X1_26/A CLKBUF1_43/Y INVX1_117/A gnd vdd DFFPOSX1
XDFFPOSX1_75 AOI22X1_37/A CLKBUF1_51/Y INVX1_128/A gnd vdd DFFPOSX1
XDFFPOSX1_97 INVX1_210/A CLKBUF1_30/Y OAI21X1_135/C gnd vdd DFFPOSX1
XFILL_42_0_1 gnd vdd FILL
XNAND3X1_314 INVX1_631/Y BUFX4_101/Y BUFX4_166/Y gnd NAND3X1_315/B vdd NAND3X1
XNAND3X1_303 BUFX4_119/Y NAND3X1_302/Y NAND2X1_883/Y gnd NAND2X1_884/B vdd NAND3X1
XNAND3X1_336 NOR2X1_442/Y AOI22X1_126/Y NOR3X1_71/Y gnd NOR2X1_462/A vdd NAND3X1
XNAND3X1_325 BUFX4_96/Y NAND3X1_325/B BUFX4_119/Y gnd BUFX4_27/A vdd NAND3X1
XNAND3X1_347 INVX1_715/A INVX1_716/Y NOR2X1_466/Y gnd NOR3X1_78/C vdd NAND3X1
XNAND3X1_358 data_memory_interface_data[15] NOR2X1_477/Y INVX4_13/A gnd OAI22X1_60/C
+ vdd NAND3X1
XFILL_33_0_1 gnd vdd FILL
XFILL_15_2 gnd vdd FILL
XDFFPOSX1_402 OR2X2_55/B CLKBUF1_46/Y OAI21X1_59/Y gnd vdd DFFPOSX1
XDFFPOSX1_413 INVX1_225/A CLKBUF1_20/Y NOR3X1_20/Y gnd vdd DFFPOSX1
XDFFPOSX1_424 INVX2_73/A CLKBUF1_39/Y NOR3X1_31/Y gnd vdd DFFPOSX1
XDFFPOSX1_446 NAND3X1_18/A CLKBUF1_10/Y INVX2_72/A gnd vdd DFFPOSX1
XDFFPOSX1_435 BUFX2_94/A CLKBUF1_13/Y NOR3X1_42/Y gnd vdd DFFPOSX1
XDFFPOSX1_457 NAND3X1_40/A CLKBUF1_10/Y BUFX2_56/A gnd vdd DFFPOSX1
XDFFPOSX1_479 BUFX2_46/A CLKBUF1_7/Y NAND3X1_21/Y gnd vdd DFFPOSX1
XDFFPOSX1_468 NAND3X1_62/A CLKBUF1_47/Y BUFX2_67/A gnd vdd DFFPOSX1
XINVX1_191 NOR2X1_11/Y gnd INVX1_191/Y vdd INVX1
XNAND2X1_527 BUFX4_214/Y NAND2X1_547/B gnd NAND2X1_527/Y vdd NAND2X1
XNAND2X1_516 BUFX4_127/Y NOR2X1_368/B gnd OAI22X1_30/D vdd NAND2X1
XNAND2X1_505 NAND2X1_501/Y NAND2X1_505/B gnd OR2X2_33/A vdd NAND2X1
XINVX1_180 instruction_memory_interface_data[24] gnd INVX1_180/Y vdd INVX1
XNAND2X1_549 BUFX4_125/Y NAND2X1_549/B gnd OAI21X1_635/C vdd NAND2X1
XNAND2X1_538 BUFX4_214/Y NAND2X1_556/B gnd NAND2X1_538/Y vdd NAND2X1
XFILL_24_0_1 gnd vdd FILL
XAOI21X1_140 AOI21X1_54/B AOI21X1_89/A OAI21X1_598/Y gnd AOI21X1_140/Y vdd AOI21X1
XAOI21X1_151 INVX4_7/A NOR2X1_207/B NAND3X1_143/Y gnd AOI21X1_151/Y vdd AOI21X1
XAOI21X1_173 AOI21X1_173/A NAND2X1_567/Y INVX2_65/Y gnd NOR3X1_61/B vdd AOI21X1
XAOI21X1_184 INVX1_417/Y NOR2X1_341/Y INVX1_418/Y gnd OAI21X1_708/C vdd AOI21X1
XAOI21X1_162 INVX4_7/A AOI22X1_83/A NAND3X1_150/Y gnd AOI21X1_162/Y vdd AOI21X1
XAOI21X1_195 OAI21X1_750/B NAND2X1_578/Y INVX2_18/A gnd NOR2X1_355/B vdd AOI21X1
XFILL_7_1_1 gnd vdd FILL
XFILL_15_0_1 gnd vdd FILL
XNAND3X1_111 NAND3X1_111/A OAI21X1_448/Y AOI21X1_73/Y gnd INVX1_69/A vdd NAND3X1
XNAND3X1_122 NAND3X1_122/A AOI22X1_90/Y AOI21X1_95/Y gnd INVX1_74/A vdd NAND3X1
XNAND3X1_100 INVX2_41/Y INVX2_40/Y NOR2X1_170/Y gnd OR2X2_21/B vdd NAND3X1
XNAND3X1_133 INVX2_58/A INVX4_8/A AOI22X1_96/Y gnd NOR2X1_296/A vdd NAND3X1
XNAND3X1_144 INVX8_11/Y NAND3X1_146/C NAND3X1_144/C gnd NAND3X1_144/Y vdd NAND3X1
XNAND3X1_155 INVX8_11/Y NAND3X1_155/B OR2X2_38/Y gnd NAND3X1_155/Y vdd NAND3X1
XNAND3X1_166 BUFX4_93/Y OAI21X1_741/Y NAND3X1_166/C gnd NAND3X1_167/B vdd NAND3X1
XNAND3X1_188 BUFX4_208/Y NOR2X1_401/Y AOI21X1_223/Y gnd BUFX4_204/A vdd NAND3X1
XNAND3X1_177 BUFX4_93/Y NAND3X1_177/B NAND3X1_177/C gnd NAND3X1_178/C vdd NAND3X1
XNAND3X1_199 BUFX4_218/Y NAND3X1_199/B NAND3X1_199/C gnd NAND2X1_723/B vdd NAND3X1
XOAI21X1_329 NOR2X1_126/Y OAI21X1_329/B NAND3X1_93/C gnd NAND2X1_308/B vdd OAI21X1
XOAI21X1_307 INVX1_330/Y INVX4_4/A OAI21X1_307/C gnd MUX2X1_39/A vdd OAI21X1
XOAI21X1_318 INVX1_369/A INVX2_52/A AOI21X1_63/A gnd AOI21X1_40/B vdd OAI21X1
XBUFX4_5 CLK gnd BUFX4_5/Y vdd BUFX4
XDFFPOSX1_210 INVX1_722/A CLKBUF1_8/Y OR2X2_56/B gnd vdd DFFPOSX1
XDFFPOSX1_221 AOI22X1_171/C CLKBUF1_38/Y INVX1_467/A gnd vdd DFFPOSX1
XDFFPOSX1_254 MUX2X1_13/A CLKBUF1_17/Y NAND3X1_8/A gnd vdd DFFPOSX1
XDFFPOSX1_232 OAI21X1_117/C CLKBUF1_53/Y INVX1_76/A gnd vdd DFFPOSX1
XDFFPOSX1_243 OAI21X1_139/C CLKBUF1_63/Y INVX1_87/A gnd vdd DFFPOSX1
XDFFPOSX1_265 MUX2X1_7/A CLKBUF1_54/Y NAND3X1_28/A gnd vdd DFFPOSX1
XNAND2X1_302 INVX2_40/A MUX2X1_5/Y gnd NAND2X1_500/A vdd NAND2X1
XDFFPOSX1_276 AOI22X1_59/A CLKBUF1_27/Y NAND3X1_50/A gnd vdd DFFPOSX1
XDFFPOSX1_298 OR2X2_17/B CLKBUF1_44/Y NOR3X1_3/Y gnd vdd DFFPOSX1
XDFFPOSX1_287 AND2X2_1/A CLKBUF1_34/Y NAND3X1_6/Y gnd vdd DFFPOSX1
XNAND2X1_324 BUFX4_44/Y MUX2X1_12/Y gnd OAI21X1_342/C vdd NAND2X1
XNAND2X1_313 NOR2X1_6/A OR2X2_44/A gnd NOR2X1_132/B vdd NAND2X1
XNAND2X1_335 BUFX4_40/Y INVX2_27/A gnd NAND2X1_335/Y vdd NAND2X1
XNAND2X1_368 BUFX4_39/Y NOR2X1_94/B gnd OAI21X1_631/C vdd NAND2X1
XNAND2X1_357 NOR2X1_195/A INVX2_52/Y gnd OAI21X1_375/C vdd NAND2X1
XNAND2X1_346 INVX1_377/A AND2X2_23/Y gnd INVX4_5/A vdd NAND2X1
XNAND2X1_379 BUFX4_44/Y MUX2X1_11/Y gnd OAI21X1_393/C vdd NAND2X1
XNOR3X1_53 INVX1_254/Y AOI21X1_4/C NOR3X1_49/C gnd NOR3X1_53/Y vdd NOR3X1
XNOR3X1_42 NOR3X1_3/A INVX1_183/Y BUFX4_49/Y gnd NOR3X1_42/Y vdd NOR3X1
XNOR3X1_20 INVX4_1/A INVX1_161/Y NOR3X1_8/C gnd NOR3X1_20/Y vdd NOR3X1
XNOR3X1_31 NOR3X1_35/A INVX1_172/Y BUFX4_48/Y gnd NOR3X1_31/Y vdd NOR3X1
XNOR3X1_64 NOR3X1_64/A NOR3X1_64/B NOR3X1_64/C gnd NOR3X1_64/Y vdd NOR3X1
XNOR3X1_75 INVX2_88/A INVX2_89/A NOR3X1_75/C gnd NOR3X1_75/Y vdd NOR3X1
XNOR2X1_390 INVX1_480/A NOR2X1_390/B gnd AND2X2_78/A vdd NOR2X1
XINVX4_5 INVX4_5/A gnd INVX4_5/Y vdd INVX4
XOAI21X1_841 NOR3X1_66/C INVX1_478/Y INVX1_479/Y gnd OAI21X1_841/Y vdd OAI21X1
XOAI21X1_830 NAND2X1_654/Y INVX1_474/Y INVX1_475/Y gnd OAI21X1_830/Y vdd OAI21X1
XOAI21X1_874 BUFX2_87/A INVX1_640/Y NAND2X1_915/Y gnd OAI21X1_874/Y vdd OAI21X1
XOAI21X1_852 OAI21X1_851/Y INVX8_13/A OAI21X1_852/C gnd OAI21X1_182/C vdd OAI21X1
XOAI21X1_863 NOR3X1_68/C INVX1_488/Y INVX1_489/Y gnd OAI21X1_863/Y vdd OAI21X1
XOAI21X1_885 INVX1_656/Y OAI21X1_887/B INVX4_11/Y gnd OAI21X1_885/Y vdd OAI21X1
XOAI21X1_896 INVX8_14/Y AOI21X1_231/Y AOI22X1_120/Y gnd OAI21X1_896/Y vdd OAI21X1
XNAND2X1_880 INVX1_616/Y BUFX4_98/Y gnd NAND3X1_301/C vdd NAND2X1
XNAND2X1_891 OAI21X1_89/Y BUFX4_63/Y gnd NAND2X1_891/Y vdd NAND2X1
XNAND3X1_8 NAND3X1_8/A AND2X2_2/B AND2X2_2/A gnd AOI21X1_1/A vdd NAND3X1
XOAI21X1_104 BUFX4_184/Y INVX1_102/Y OAI21X1_104/C gnd INVX1_583/A vdd OAI21X1
XOAI21X1_115 BUFX4_273/Y BUFX4_193/Y OAI21X1_115/C gnd OAI21X1_115/Y vdd OAI21X1
XOAI21X1_126 BUFX4_184/Y INVX1_113/Y OAI21X1_125/Y gnd INVX1_532/A vdd OAI21X1
XOAI21X1_137 BUFX4_270/Y OR2X2_2/B DFFPOSX1_98/D gnd OAI21X1_137/Y vdd OAI21X1
XOAI21X1_148 BUFX4_183/Y INVX1_124/Y OAI21X1_147/Y gnd INVX1_554/A vdd OAI21X1
XOAI21X1_159 OR2X2_2/A BUFX4_194/Y OAI21X1_159/C gnd OAI21X1_159/Y vdd OAI21X1
XBUFX2_2 gnd gnd data_memory_interface_address[1] vdd BUFX2
XNAND2X1_110 INVX1_226/Y INVX1_227/Y gnd NOR2X1_16/B vdd NAND2X1
XNAND2X1_143 XNOR2X1_17/Y XNOR2X1_20/Y gnd NOR2X1_38/B vdd NAND2X1
XNAND2X1_132 INVX1_690/A BUFX4_147/Y gnd NAND3X1_81/C vdd NAND2X1
XNAND2X1_121 AOI21X1_6/B OR2X2_9/Y gnd XNOR2X1_5/A vdd NAND2X1
XNAND2X1_154 INVX1_261/Y INVX1_260/A gnd NAND2X1_155/A vdd NAND2X1
XNAND2X1_176 NOR2X1_47/Y NOR2X1_46/Y gnd NOR2X1_48/B vdd NAND2X1
XNAND2X1_165 NAND3X1_84/Y NAND2X1_163/Y gnd OR2X2_11/A vdd NAND2X1
XNAND2X1_187 INVX1_282/A NOR2X1_57/Y gnd INVX1_287/A vdd NAND2X1
XNAND2X1_198 INVX4_4/A AOI22X1_62/A gnd NAND2X1_198/Y vdd NAND2X1
XFILL_41_6_0 gnd vdd FILL
XINVX2_2 INVX2_2/A gnd INVX2_2/Y vdd INVX2
XOAI21X1_660 INVX1_410/Y INVX2_69/Y NAND3X1_89/B gnd NOR2X1_325/A vdd OAI21X1
XOAI21X1_693 NOR2X1_336/B INVX1_417/A INVX1_418/A gnd AOI21X1_176/C vdd OAI21X1
XOAI21X1_682 AOI21X1_38/A NOR2X1_333/Y AOI21X1_168/B gnd OAI21X1_682/Y vdd OAI21X1
XOAI21X1_671 OAI21X1_700/A INVX8_5/A NAND2X1_564/Y gnd MUX2X1_45/A vdd OAI21X1
XAOI21X1_2 NAND3X1_9/Y AOI21X1_2/B reset gnd AOI21X1_2/Y vdd AOI21X1
XINVX1_702 OR2X2_54/B gnd INVX1_702/Y vdd INVX1
XINVX1_735 data_memory_interface_data[0] gnd INVX1_735/Y vdd INVX1
XINVX1_713 AND2X2_93/B gnd INVX1_713/Y vdd INVX1
XINVX1_724 INVX1_724/A gnd INVX1_724/Y vdd INVX1
XINVX1_757 INVX1_757/A gnd INVX1_757/Y vdd INVX1
XINVX1_746 data_memory_interface_data[4] gnd INVX1_746/Y vdd INVX1
XXNOR2X1_21 NOR2X1_31/B INVX2_9/Y gnd NOR2X1_34/A vdd XNOR2X1
XXNOR2X1_32 XNOR2X1_32/A NOR2X1_47/A gnd XNOR2X1_32/Y vdd XNOR2X1
XXNOR2X1_10 XNOR2X1_10/A XNOR2X1_9/Y gnd XNOR2X1_10/Y vdd XNOR2X1
XXNOR2X1_43 XNOR2X1_28/A INVX2_11/Y gnd NOR2X1_46/A vdd XNOR2X1
XXNOR2X1_54 INVX1_689/A INVX1_443/A gnd AND2X2_95/A vdd XNOR2X1
XBUFX2_20 BUFX2_20/A gnd data_memory_interface_address[19] vdd BUFX2
XBUFX2_53 BUFX2_53/A gnd instruction_memory_interface_address[14] vdd BUFX2
XBUFX2_42 BUFX2_42/A gnd instruction_memory_interface_address[3] vdd BUFX2
XBUFX2_31 BUFX2_31/A gnd data_memory_interface_address[30] vdd BUFX2
XBUFX2_75 vdd gnd instruction_memory_interface_frame_mask[3] vdd BUFX2
XBUFX2_64 BUFX2_64/A gnd instruction_memory_interface_address[25] vdd BUFX2
XBUFX2_86 BUFX2_86/A gnd BUFX2_86/Y vdd BUFX2
XBUFX2_97 BUFX2_97/A gnd BUFX2_97/Y vdd BUFX2
XFILL_32_6_0 gnd vdd FILL
XFILL_23_6_0 gnd vdd FILL
XAOI21X1_10 NOR2X1_29/Y INVX1_240/A INVX1_244/Y gnd AOI21X1_10/Y vdd AOI21X1
XAOI21X1_43 NOR2X1_108/Y AOI21X1_43/B AOI21X1_43/C gnd AOI21X1_43/Y vdd AOI21X1
XAOI21X1_21 XNOR2X1_33/Y XNOR2X1_32/A NOR2X1_37/Y gnd XNOR2X1_35/A vdd AOI21X1
XAOI21X1_32 INVX1_293/A AOI21X1_32/B NOR2X1_64/A gnd NOR2X1_61/B vdd AOI21X1
XAOI21X1_76 OR2X2_18/Y AOI21X1_47/B BUFX4_54/Y gnd OAI22X1_21/A vdd AOI21X1
XAOI21X1_65 NOR2X1_194/Y INVX1_372/Y AOI21X1_65/C gnd AOI21X1_65/Y vdd AOI21X1
XAOI21X1_54 BUFX4_83/Y AOI21X1_54/B BUFX4_124/Y gnd AOI21X1_54/Y vdd AOI21X1
XAOI21X1_87 OAI22X1_15/B AOI21X1_87/B INVX2_57/Y gnd AOI21X1_87/Y vdd AOI21X1
XAOI21X1_98 AOI21X1_98/A NOR2X1_232/A AOI22X1_86/A gnd AOI21X1_98/Y vdd AOI21X1
XOAI21X1_5 INVX1_5/Y BUFX4_21/Y OAI21X1_5/C gnd OAI21X1_5/Y vdd OAI21X1
XFILL_6_7_0 gnd vdd FILL
XFILL_14_6_0 gnd vdd FILL
XOAI22X1_40 MUX2X1_50/B OAI22X1_40/B MUX2X1_52/Y OR2X2_33/B gnd OAI22X1_40/Y vdd OAI22X1
XOAI22X1_51 AND2X2_89/Y OAI22X1_51/B AND2X2_90/Y OAI22X1_51/D gnd NOR3X1_71/B vdd
+ OAI22X1
XOAI21X1_490 NOR2X1_228/Y NAND2X1_460/Y NOR2X1_230/Y gnd NOR2X1_231/B vdd OAI21X1
XINVX1_510 INVX1_583/A gnd INVX1_510/Y vdd INVX1
XINVX1_543 INVX1_543/A gnd INVX1_543/Y vdd INVX1
XINVX1_554 INVX1_554/A gnd INVX1_554/Y vdd INVX1
XINVX1_532 INVX1_532/A gnd INVX1_532/Y vdd INVX1
XINVX1_521 INVX1_521/A gnd INVX1_521/Y vdd INVX1
XINVX1_565 INVX1_565/A gnd INVX1_565/Y vdd INVX1
XINVX1_576 INVX1_503/A gnd INVX1_576/Y vdd INVX1
XINVX1_587 INVX1_514/A gnd INVX1_587/Y vdd INVX1
XINVX1_598 INVX1_525/A gnd INVX1_598/Y vdd INVX1
XFILL_3_2 gnd vdd FILL
XFILL_38_1 gnd vdd FILL
XXOR2X1_8 XOR2X1_8/A XOR2X1_8/B gnd XOR2X1_8/Y vdd XOR2X1
XMUX2X1_9 MUX2X1_9/A MUX2X1_9/B INVX4_4/A gnd MUX2X1_9/Y vdd MUX2X1
XAOI22X1_120 OAI22X1_49/A INVX4_11/A BUFX4_263/Y BUFX2_92/A gnd AOI22X1_120/Y vdd
+ AOI22X1
XAOI22X1_142 data_memory_interface_data[5] BUFX4_107/Y AOI22X1_142/C BUFX4_9/Y gnd
+ AOI22X1_142/Y vdd AOI22X1
XAOI22X1_131 OR2X2_60/Y AOI22X1_131/B AOI22X1_131/C OR2X2_61/Y gnd AOI22X1_131/Y vdd
+ AOI22X1
XAOI22X1_153 data_memory_interface_data[17] BUFX4_108/Y BUFX4_172/Y BUFX4_251/Y gnd
+ AOI22X1_153/Y vdd AOI22X1
XAOI22X1_164 data_memory_interface_data[28] BUFX4_108/Y BUFX4_172/Y BUFX4_250/Y gnd
+ AOI22X1_164/Y vdd AOI22X1
XBUFX4_115 BUFX4_118/A gnd BUFX4_115/Y vdd BUFX4
XBUFX4_126 INVX8_7/Y gnd BUFX4_126/Y vdd BUFX4
XBUFX4_137 OAI22X1_1/Y gnd BUFX4_137/Y vdd BUFX4
XBUFX4_104 BUFX4_107/A gnd INVX4_14/A vdd BUFX4
XBUFX4_148 BUFX4_148/A gnd BUFX4_148/Y vdd BUFX4
XBUFX4_159 NOR2X1_2/Y gnd BUFX4_159/Y vdd BUFX4
XNOR2X1_219 INVX1_378/A AOI21X1_74/Y gnd NOR2X1_220/A vdd NOR2X1
XNOR2X1_208 INVX4_5/A NOR2X1_207/Y gnd NOR2X1_208/Y vdd NOR2X1
XOAI21X1_1027 BUFX4_65/Y BUFX4_69/Y AOI22X1_148/Y gnd OAI21X1_1027/Y vdd OAI21X1
XOAI21X1_1005 INVX1_750/Y OAI21X1_993/B NAND2X1_1017/Y gnd AOI22X1_143/C vdd OAI21X1
XOAI21X1_1016 NOR2X1_481/Y INVX4_12/A data_memory_interface_data[25] gnd OAI21X1_1016/Y
+ vdd OAI21X1
XOAI21X1_1038 BUFX4_66/Y BUFX4_71/Y AOI22X1_154/Y gnd OAI21X1_1038/Y vdd OAI21X1
XOAI21X1_1049 BUFX4_67/Y BUFX4_70/Y AOI22X1_165/Y gnd OAI21X1_1049/Y vdd OAI21X1
XINVX1_362 INVX1_362/A gnd INVX1_362/Y vdd INVX1
XINVX1_351 INVX1_351/A gnd INVX1_351/Y vdd INVX1
XINVX1_340 OR2X2_64/A gnd INVX1_340/Y vdd INVX1
XINVX1_373 INVX1_373/A gnd INVX1_373/Y vdd INVX1
XINVX1_384 INVX1_384/A gnd INVX1_384/Y vdd INVX1
XINVX1_395 INVX1_395/A gnd INVX1_395/Y vdd INVX1
XNAND2X1_709 INVX2_75/A INVX1_495/Y gnd NAND2X1_709/Y vdd NAND2X1
XFILL_37_5_0 gnd vdd FILL
XFILL_20_4_0 gnd vdd FILL
XNAND2X1_1010 NAND3X1_352/Y NOR2X1_480/Y gnd BUFX2_38/A vdd NAND2X1
XDFFPOSX1_10 AOI22X1_10/D CLKBUF1_49/Y DFFPOSX1_10/D gnd vdd DFFPOSX1
XDFFPOSX1_43 DFFPOSX1_43/Q CLKBUF1_43/Y INVX1_502/A gnd vdd DFFPOSX1
XDFFPOSX1_21 AOI22X1_21/D CLKBUF1_18/Y DFFPOSX1_21/D gnd vdd DFFPOSX1
XDFFPOSX1_54 AOI22X1_16/A CLKBUF1_15/Y INVX1_107/A gnd vdd DFFPOSX1
XDFFPOSX1_32 AOI22X1_32/D CLKBUF1_24/Y DFFPOSX1_32/D gnd vdd DFFPOSX1
XNAND2X1_1021 BUFX2_77/A BUFX4_118/Y gnd NAND3X1_359/C vdd NAND2X1
XDFFPOSX1_87 INVX1_200/A CLKBUF1_2/Y OAI21X1_115/C gnd vdd DFFPOSX1
XDFFPOSX1_76 AOI22X1_38/A CLKBUF1_50/Y INVX1_129/A gnd vdd DFFPOSX1
XDFFPOSX1_65 AOI22X1_27/A CLKBUF1_55/Y INVX1_118/A gnd vdd DFFPOSX1
XDFFPOSX1_98 INVX1_211/A CLKBUF1_3/Y DFFPOSX1_98/D gnd vdd DFFPOSX1
XFILL_3_5_0 gnd vdd FILL
XFILL_28_5_0 gnd vdd FILL
XNAND3X1_315 BUFX4_121/Y NAND3X1_315/B NAND3X1_315/C gnd NAND2X1_902/B vdd NAND3X1
XNAND3X1_304 INVX1_621/Y BUFX4_99/Y BUFX4_167/Y gnd NAND3X1_305/B vdd NAND3X1
XNAND3X1_337 NAND3X1_337/A AOI22X1_135/Y INVX1_699/Y gnd NAND3X1_337/Y vdd NAND3X1
XNAND3X1_326 OAI22X1_6/Y BUFX2_87/A NOR2X1_412/Y gnd NAND3X1_327/C vdd NAND3X1
XNAND3X1_348 INVX2_88/Y NAND3X1_1/B NOR2X1_470/Y gnd NOR2X1_471/B vdd NAND3X1
XFILL_11_4_0 gnd vdd FILL
XNAND3X1_359 NAND3X1_359/A NAND3X1_359/B NAND3X1_359/C gnd NAND3X1_359/Y vdd NAND3X1
XFILL_19_5_0 gnd vdd FILL
XDFFPOSX1_403 OR2X2_54/B CLKBUF1_46/Y OAI21X1_60/Y gnd vdd DFFPOSX1
XDFFPOSX1_447 NAND3X1_20/A CLKBUF1_33/Y BUFX2_46/A gnd vdd DFFPOSX1
XDFFPOSX1_436 BUFX2_95/A CLKBUF1_13/Y NOR3X1_43/Y gnd vdd DFFPOSX1
XDFFPOSX1_414 INVX2_4/A CLKBUF1_20/Y NOR3X1_21/Y gnd vdd DFFPOSX1
XDFFPOSX1_425 OR2X2_50/B CLKBUF1_9/Y NOR3X1_32/Y gnd vdd DFFPOSX1
XDFFPOSX1_458 NAND3X1_42/A CLKBUF1_45/Y BUFX2_57/A gnd vdd DFFPOSX1
XDFFPOSX1_469 NAND3X1_64/A CLKBUF1_36/Y BUFX2_68/A gnd vdd DFFPOSX1
XINVX1_170 instruction_memory_interface_data[14] gnd INVX1_170/Y vdd INVX1
XINVX1_192 INVX1_192/A gnd INVX1_192/Y vdd INVX1
XNAND2X1_517 BUFX4_84/Y NOR2X1_368/B gnd MUX2X1_55/A vdd NAND2X1
XNAND2X1_506 BUFX4_56/Y NOR2X1_218/Y gnd OR2X2_42/B vdd NAND2X1
XINVX1_181 instruction_memory_interface_data[25] gnd INVX1_181/Y vdd INVX1
XNAND2X1_539 BUFX4_51/Y OAI21X1_719/A gnd OAI21X1_614/C vdd NAND2X1
XNAND2X1_528 BUFX4_56/Y NOR2X1_236/Y gnd INVX1_397/A vdd NAND2X1
XAOI21X1_141 AOI22X1_72/B NOR2X1_305/Y NOR2X1_248/Y gnd OAI21X1_601/B vdd AOI21X1
XAOI21X1_130 NOR2X1_296/Y OAI21X1_513/C AOI21X1_130/C gnd OAI21X1_694/A vdd AOI21X1
XAOI21X1_152 INVX4_9/A MUX2X1_34/A AOI21X1_152/C gnd NOR2X1_318/A vdd AOI21X1
XAOI21X1_185 NOR2X1_342/Y AOI21X1_185/B OAI21X1_708/Y gnd OAI21X1_743/A vdd AOI21X1
XAOI21X1_163 NAND2X1_561/Y AOI21X1_163/B INVX8_7/A gnd OAI21X1_663/A vdd AOI21X1
XAOI21X1_174 INVX4_7/A AOI22X1_87/B AOI21X1_174/C gnd OAI21X1_690/C vdd AOI21X1
XAOI21X1_196 INVX1_422/A OAI21X1_734/Y BUFX4_276/Y gnd OAI21X1_735/C vdd AOI21X1
XFILL_43_3_0 gnd vdd FILL
XNAND3X1_123 INVX2_58/A OAI21X1_526/B NAND3X1_123/C gnd AOI22X1_92/D vdd NAND3X1
XNAND3X1_112 NAND3X1_112/A OR2X2_27/Y AOI21X1_80/Y gnd INVX1_70/A vdd NAND3X1
XNAND3X1_101 AND2X2_20/Y NOR2X1_177/Y NOR2X1_129/Y gnd NAND3X1_101/Y vdd NAND3X1
XNAND3X1_145 OAI21X1_620/Y NAND3X1_144/Y NOR3X1_58/Y gnd INVX1_84/A vdd NAND3X1
XNAND3X1_134 NAND3X1_134/A NAND3X1_134/B AOI21X1_115/Y gnd AOI21X1_116/C vdd NAND3X1
XNAND3X1_156 BUFX4_90/Y NAND3X1_156/B NAND2X1_569/Y gnd NAND3X1_157/A vdd NAND3X1
XNAND3X1_167 NAND3X1_167/A NAND3X1_167/B AOI21X1_198/Y gnd INVX1_93/A vdd NAND3X1
XNAND3X1_178 AOI21X1_213/Y NAND3X1_178/B NAND3X1_178/C gnd INVX1_97/A vdd NAND3X1
XNAND3X1_189 NAND3X1_189/A NAND2X1_708/Y NAND2X1_709/Y gnd NOR2X1_402/A vdd NAND3X1
XFILL_34_3_0 gnd vdd FILL
XFILL_20_1 gnd vdd FILL
XOAI21X1_319 NOR2X1_110/Y AOI22X1_81/C AOI22X1_81/B gnd AOI21X1_40/C vdd OAI21X1
XOAI21X1_308 INVX1_331/Y INVX4_4/A NAND2X1_244/Y gnd MUX2X1_37/B vdd OAI21X1
XBUFX4_6 CLK gnd BUFX4_6/Y vdd BUFX4
XDFFPOSX1_222 OAI21X1_97/C CLKBUF1_21/Y INVX1_65/A gnd vdd DFFPOSX1
XDFFPOSX1_211 INVX1_723/A CLKBUF1_28/Y INVX1_457/A gnd vdd DFFPOSX1
XDFFPOSX1_200 INVX1_728/A CLKBUF1_28/Y OR2X2_59/B gnd vdd DFFPOSX1
XDFFPOSX1_255 MUX2X1_14/A CLKBUF1_47/Y NAND3X1_9/A gnd vdd DFFPOSX1
XDFFPOSX1_244 OAI21X1_141/C CLKBUF1_2/Y INVX1_88/A gnd vdd DFFPOSX1
XDFFPOSX1_233 OAI21X1_119/C CLKBUF1_21/Y INVX1_77/A gnd vdd DFFPOSX1
XDFFPOSX1_266 MUX2X1_5/A CLKBUF1_14/Y NAND3X1_30/A gnd vdd DFFPOSX1
XDFFPOSX1_277 AOI22X1_60/A CLKBUF1_17/Y NAND3X1_52/A gnd vdd DFFPOSX1
XDFFPOSX1_288 INVX1_66/A CLKBUF1_34/Y NOR3X1_12/Y gnd vdd DFFPOSX1
XNAND2X1_325 BUFX4_39/Y NOR2X1_151/B gnd OAI21X1_452/C vdd NAND2X1
XNAND2X1_303 INVX2_41/A MUX2X1_6/Y gnd OAI21X1_330/C vdd NAND2X1
XNAND2X1_336 MUX2X1_20/S MUX2X1_26/A gnd OAI21X1_359/C vdd NAND2X1
XNAND2X1_314 INVX1_347/Y INVX1_355/A gnd NOR2X1_135/B vdd NAND2X1
XDFFPOSX1_299 OR2X2_17/A CLKBUF1_56/Y NOR3X1_4/Y gnd vdd DFFPOSX1
XNAND2X1_369 BUFX4_39/Y MUX2X1_42/A gnd OAI21X1_385/C vdd NAND2X1
XNAND2X1_358 NOR2X1_182/Y BUFX4_85/Y gnd NOR2X1_299/B vdd NAND2X1
XNAND2X1_347 INVX2_51/Y AND2X2_24/Y gnd NOR2X1_176/B vdd NAND2X1
XNOR3X1_10 NOR3X1_9/A INVX1_147/Y NOR3X1_9/C gnd NOR3X1_10/Y vdd NOR3X1
XNOR3X1_43 NOR3X1_3/A INVX1_184/Y BUFX4_49/Y gnd NOR3X1_43/Y vdd NOR3X1
XNOR3X1_21 INVX4_1/A INVX1_162/Y BUFX4_45/Y gnd NOR3X1_21/Y vdd NOR3X1
XNOR3X1_32 NOR3X1_35/A INVX1_173/Y NOR3X1_8/C gnd NOR3X1_32/Y vdd NOR3X1
XNOR3X1_54 INVX1_257/Y AOI21X1_4/C NOR3X1_49/C gnd NOR3X1_54/Y vdd NOR3X1
XNOR3X1_65 OR2X2_46/Y OR2X2_47/Y NOR3X1_65/C gnd NOR3X1_65/Y vdd NOR3X1
XNOR3X1_76 NOR3X1_76/A NOR2X1_3/B OR2X2_69/Y gnd NOR3X1_76/Y vdd NOR3X1
XFILL_0_3_0 gnd vdd FILL
XFILL_25_3_0 gnd vdd FILL
XNOR2X1_380 BUFX2_41/A BUFX2_42/A gnd NOR2X1_380/Y vdd NOR2X1
XNOR2X1_391 OR2X2_48/B OR2X2_48/A gnd NOR2X1_392/B vdd NOR2X1
XINVX4_6 INVX4_6/A gnd INVX4_6/Y vdd INVX4
XOAI21X1_842 NOR3X1_66/C INVX1_480/A OAI21X1_841/Y gnd OAI21X1_843/A vdd OAI21X1
XOAI21X1_820 INVX1_471/Y BUFX2_44/A INVX8_13/Y gnd OAI21X1_820/Y vdd OAI21X1
XOAI21X1_831 NOR3X1_65/C OR2X2_46/Y OAI21X1_830/Y gnd OAI21X1_831/Y vdd OAI21X1
XOAI21X1_875 INVX2_76/Y DFFPOSX1_41/Q OAI21X1_875/C gnd NOR2X1_410/B vdd OAI21X1
XOAI21X1_853 OR2X2_48/Y INVX1_485/Y INVX8_13/Y gnd OAI21X1_853/Y vdd OAI21X1
XOAI21X1_864 NOR3X1_68/C INVX1_490/Y OAI21X1_863/Y gnd OAI21X1_864/Y vdd OAI21X1
XOAI21X1_897 INVX8_14/Y AOI21X1_231/Y AOI22X1_121/Y gnd OAI21X1_897/Y vdd OAI21X1
XOAI21X1_886 INVX1_657/Y OAI21X1_887/B INVX4_11/Y gnd OAI21X1_886/Y vdd OAI21X1
XFILL_8_4_0 gnd vdd FILL
XNAND2X1_870 OAI21X1_82/Y BUFX4_60/Y gnd NAND2X1_870/Y vdd NAND2X1
XNAND2X1_881 NAND2X1_879/Y NAND2X1_881/B gnd NAND2X1_53/B vdd NAND2X1
XNAND2X1_892 INVX1_624/Y BUFX4_97/Y gnd NAND3X1_309/C vdd NAND2X1
XFILL_16_3_0 gnd vdd FILL
XNAND3X1_9 NAND3X1_9/A AND2X2_2/B AND2X2_2/A gnd NAND3X1_9/Y vdd NAND3X1
XOAI21X1_116 BUFX4_183/Y INVX1_108/Y OAI21X1_115/Y gnd INVX1_595/A vdd OAI21X1
XOAI21X1_127 BUFX4_272/Y BUFX4_195/Y OAI21X1_127/C gnd OAI21X1_128/C vdd OAI21X1
XOAI21X1_105 BUFX4_269/Y BUFX4_193/Y OAI21X1_105/C gnd OAI21X1_106/C vdd OAI21X1
XOAI21X1_138 BUFX4_185/Y INVX1_119/Y OAI21X1_137/Y gnd INVX1_617/A vdd OAI21X1
XOAI21X1_149 BUFX4_270/Y OR2X2_2/B OAI21X1_149/C gnd OAI21X1_150/C vdd OAI21X1
XBUFX2_3 BUFX2_3/A gnd data_memory_interface_address[2] vdd BUFX2
XNAND2X1_100 AND2X2_3/B AND2X2_3/A gnd OAI22X1_1/B vdd NAND2X1
XNAND2X1_133 INVX1_247/A BUFX4_231/Y gnd NAND3X1_81/B vdd NAND2X1
XNAND2X1_144 AOI21X1_17/A XNOR2X1_24/Y gnd NOR2X1_38/A vdd NAND2X1
XNAND2X1_122 AOI21X1_7/Y NAND3X1_78/Y gnd INVX1_240/A vdd NAND2X1
XNAND2X1_111 INVX1_225/A INVX1_228/Y gnd OR2X2_6/A vdd NAND2X1
XNAND2X1_155 NAND2X1_155/A NAND2X1_153/Y gnd XOR2X1_3/B vdd NAND2X1
XNAND2X1_177 AND2X2_15/Y AND2X2_14/Y gnd AOI21X1_29/C vdd NAND2X1
XNAND2X1_166 INVX1_270/Y OAI21X1_263/Y gnd INVX1_272/A vdd NAND2X1
XNAND2X1_199 INVX4_4/A AOI22X1_61/A gnd NAND2X1_199/Y vdd NAND2X1
XNAND2X1_188 INVX1_288/Y NOR2X1_58/B gnd AND2X2_17/B vdd NAND2X1
XFILL_41_6_1 gnd vdd FILL
XFILL_40_1_0 gnd vdd FILL
XINVX2_3 INVX2_3/A gnd INVX2_3/Y vdd INVX2
XOAI21X1_650 NAND2X1_572/B INVX8_4/A NAND2X1_551/Y gnd MUX2X1_54/B vdd OAI21X1
XOAI21X1_661 INVX4_10/Y INVX1_409/A BUFX4_90/Y gnd NOR2X1_326/A vdd OAI21X1
XOAI21X1_672 MUX2X1_45/Y OR2X2_33/B BUFX4_55/Y gnd AND2X2_56/A vdd OAI21X1
XOAI21X1_683 INVX2_29/Y INVX2_30/Y OAI21X1_682/Y gnd OR2X2_38/A vdd OAI21X1
XINVX1_703 OR2X2_55/B gnd INVX1_703/Y vdd INVX1
XAOI21X1_3 NOR2X1_22/Y AOI21X1_3/B INVX2_79/A gnd INVX1_145/A vdd AOI21X1
XOAI21X1_694 OAI21X1_694/A NAND2X1_570/Y AOI21X1_176/Y gnd AOI21X1_200/B vdd OAI21X1
XINVX1_714 INVX1_714/A gnd INVX1_714/Y vdd INVX1
XINVX1_725 INVX1_725/A gnd INVX1_725/Y vdd INVX1
XINVX1_736 data_memory_interface_data[17] gnd INVX1_736/Y vdd INVX1
XINVX1_758 BUFX4_253/Y gnd INVX1_758/Y vdd INVX1
XINVX1_747 data_memory_interface_data[21] gnd INVX1_747/Y vdd INVX1
XXNOR2X1_22 AOI21X1_17/B NOR2X1_34/A gnd XNOR2X1_22/Y vdd XNOR2X1
XXNOR2X1_11 XNOR2X1_9/A INVX2_7/A gnd AOI21X1_7/B vdd XNOR2X1
XXNOR2X1_33 NOR2X1_37/B INVX2_12/A gnd XNOR2X1_33/Y vdd XNOR2X1
XXNOR2X1_44 NOR2X1_40/B INVX2_13/Y gnd NOR2X1_47/B vdd XNOR2X1
XXNOR2X1_55 INVX1_690/A INVX1_442/A gnd AND2X2_95/B vdd XNOR2X1
XBUFX2_10 BUFX2_10/A gnd data_memory_interface_address[9] vdd BUFX2
XINVX1_90 INVX1_90/A gnd INVX1_90/Y vdd INVX1
XBUFX2_43 BUFX2_43/A gnd instruction_memory_interface_address[4] vdd BUFX2
XBUFX2_54 BUFX2_54/A gnd instruction_memory_interface_address[15] vdd BUFX2
XBUFX2_21 BUFX2_21/A gnd data_memory_interface_address[20] vdd BUFX2
XBUFX2_32 BUFX2_32/A gnd data_memory_interface_address[31] vdd BUFX2
XBUFX2_76 gnd gnd instruction_memory_interface_state vdd BUFX2
XBUFX2_65 BUFX2_65/A gnd instruction_memory_interface_address[26] vdd BUFX2
XBUFX2_87 BUFX2_87/A gnd BUFX2_87/Y vdd BUFX2
XBUFX2_98 INVX8_14/A gnd BUFX2_98/Y vdd BUFX2
XFILL_32_6_1 gnd vdd FILL
XFILL_31_1_0 gnd vdd FILL
XNOR2X1_1 NOR2X1_1/A INVX1_66/Y gnd NOR2X1_1/Y vdd NOR2X1
XFILL_39_2_0 gnd vdd FILL
XFILL_23_6_1 gnd vdd FILL
XFILL_22_1_0 gnd vdd FILL
XAOI21X1_22 NOR2X1_37/Y XNOR2X1_34/Y NOR2X1_40/Y gnd AOI21X1_22/Y vdd AOI21X1
XAOI21X1_11 AOI21X1_8/A AOI21X1_8/B INVX1_246/Y gnd AOI21X1_11/Y vdd AOI21X1
XAOI21X1_33 INVX1_270/A AND2X2_15/Y AOI21X1_33/C gnd AOI21X1_33/Y vdd AOI21X1
XAOI21X1_44 INVX1_376/A AND2X2_42/A AND2X2_26/A gnd INVX1_348/A vdd AOI21X1
XAOI21X1_77 AOI21X1_77/A AOI21X1_77/B AOI21X1_77/C gnd AOI21X1_77/Y vdd AOI21X1
XAOI21X1_66 NOR2X1_209/Y INVX4_6/Y AOI21X1_66/C gnd AOI21X1_66/Y vdd AOI21X1
XAOI21X1_55 INVX1_348/A NOR2X1_185/B INVX2_49/Y gnd INVX1_394/A vdd AOI21X1
XAOI21X1_99 NOR2X1_246/Y AOI21X1_99/B AOI21X1_99/C gnd NOR2X1_253/B vdd AOI21X1
XAOI21X1_88 AOI21X1_88/A OAI22X1_17/D AOI21X1_88/C gnd AOI21X1_88/Y vdd AOI21X1
XOAI21X1_6 INVX1_6/Y BUFX4_24/Y OAI21X1_6/C gnd OAI21X1_6/Y vdd OAI21X1
XFILL_6_7_1 gnd vdd FILL
XFILL_5_2_0 gnd vdd FILL
XOAI22X1_30 OAI22X1_30/A MUX2X1_55/A OAI22X1_30/C OAI22X1_30/D gnd NOR2X1_284/B vdd
+ OAI22X1
XFILL_13_1_0 gnd vdd FILL
XFILL_14_6_1 gnd vdd FILL
XOAI22X1_41 INVX4_7/Y OR2X2_42/B OAI22X1_43/B INVX2_22/Y gnd OAI22X1_41/Y vdd OAI22X1
XOAI22X1_52 AND2X2_96/Y NOR2X1_463/Y AND2X2_97/Y OAI22X1_52/D gnd NOR3X1_72/B vdd
+ OAI22X1
XOAI21X1_480 INVX2_57/A OAI21X1_480/B OAI22X1_18/Y gnd OAI21X1_480/Y vdd OAI21X1
XOAI21X1_491 AOI21X1_87/Y NOR2X1_232/A AND2X2_35/B gnd OAI21X1_491/Y vdd OAI21X1
XINVX1_500 INVX1_500/A gnd INVX1_500/Y vdd INVX1
XINVX1_511 INVX1_511/A gnd INVX1_511/Y vdd INVX1
XINVX1_544 INVX1_617/A gnd INVX1_544/Y vdd INVX1
XINVX1_533 INVX1_533/A gnd INVX1_533/Y vdd INVX1
XINVX1_522 INVX1_595/A gnd INVX1_522/Y vdd INVX1
XINVX1_555 INVX1_628/A gnd INVX1_555/Y vdd INVX1
XINVX1_566 INVX1_639/A gnd INVX1_566/Y vdd INVX1
XINVX1_577 INVX1_504/A gnd INVX1_577/Y vdd INVX1
XINVX1_588 INVX1_515/A gnd INVX1_588/Y vdd INVX1
XINVX1_599 INVX1_599/A gnd INVX1_599/Y vdd INVX1
XFILL_3_3 gnd vdd FILL
XFILL_38_2 gnd vdd FILL
XXOR2X1_9 XOR2X1_9/A BUFX2_64/A gnd XOR2X1_9/Y vdd XOR2X1
XAOI22X1_110 OR2X2_49/Y NAND2X1_704/Y NAND2X1_705/Y OR2X2_50/Y gnd BUFX4_210/A vdd
+ AOI22X1
XAOI22X1_121 OAI22X1_49/A INVX4_11/A BUFX4_261/Y BUFX2_93/A gnd AOI22X1_121/Y vdd
+ AOI22X1
XAOI22X1_143 data_memory_interface_data[6] BUFX4_105/Y AOI22X1_143/C BUFX4_8/Y gnd
+ AOI22X1_143/Y vdd AOI22X1
XAOI22X1_132 OR2X2_62/Y NAND2X1_956/Y AOI22X1_132/C OR2X2_63/Y gnd OAI21X1_907/C vdd
+ AOI22X1
XAOI22X1_154 data_memory_interface_data[18] BUFX4_108/Y BUFX4_170/Y BUFX4_250/Y gnd
+ AOI22X1_154/Y vdd AOI22X1
XBUFX4_127 INVX8_7/Y gnd BUFX4_127/Y vdd BUFX4
XBUFX4_116 BUFX4_118/A gnd BUFX4_116/Y vdd BUFX4
XBUFX4_105 BUFX4_107/A gnd BUFX4_105/Y vdd BUFX4
XAOI22X1_165 data_memory_interface_data[29] BUFX4_109/Y BUFX4_171/Y BUFX4_251/Y gnd
+ AOI22X1_165/Y vdd AOI22X1
XBUFX4_138 OAI22X1_1/Y gnd BUFX4_138/Y vdd BUFX4
XBUFX4_149 BUFX4_148/A gnd AND2X2_11/A vdd BUFX4
XNOR2X1_209 INVX8_3/A INVX1_389/A gnd NOR2X1_209/Y vdd NOR2X1
XOAI21X1_1028 NOR2X1_481/Y INVX4_12/A data_memory_interface_data[29] gnd OAI21X1_1029/C
+ vdd OAI21X1
XOAI21X1_1006 AOI21X1_264/Y OAI21X1_994/B AOI22X1_143/Y gnd OAI21X1_1006/Y vdd OAI21X1
XOAI21X1_1017 INVX1_739/Y INVX2_93/A OAI21X1_1016/Y gnd AOI22X1_145/C vdd OAI21X1
XOAI21X1_1039 BUFX4_66/Y BUFX4_71/Y AOI22X1_155/Y gnd OAI21X1_1039/Y vdd OAI21X1
XINVX1_330 MUX2X1_3/B gnd INVX1_330/Y vdd INVX1
XINVX1_341 INVX1_689/A gnd INVX1_341/Y vdd INVX1
XINVX1_352 INVX1_352/A gnd INVX1_352/Y vdd INVX1
XINVX1_374 INVX1_374/A gnd INVX1_374/Y vdd INVX1
XINVX1_396 INVX1_396/A gnd INVX1_396/Y vdd INVX1
XINVX1_385 INVX1_385/A gnd INVX1_385/Y vdd INVX1
XINVX1_363 INVX1_363/A gnd INVX1_363/Y vdd INVX1
XFILL_37_5_1 gnd vdd FILL
XFILL_36_0_0 gnd vdd FILL
XFILL_20_4_1 gnd vdd FILL
XNAND2X1_1011 INVX4_12/Y OAI21X1_979/Y gnd OAI21X1_981/B vdd NAND2X1
XNAND2X1_1000 AND2X2_100/Y NOR3X1_76/Y gnd INVX1_756/A vdd NAND2X1
XDFFPOSX1_11 AOI22X1_11/D CLKBUF1_55/Y DFFPOSX1_11/D gnd vdd DFFPOSX1
XDFFPOSX1_44 XOR2X1_12/B CLKBUF1_39/Y OR2X2_49/A gnd vdd DFFPOSX1
XDFFPOSX1_33 AOI22X1_33/D CLKBUF1_32/Y DFFPOSX1_33/D gnd vdd DFFPOSX1
XDFFPOSX1_22 AOI22X1_22/D CLKBUF1_42/Y DFFPOSX1_22/D gnd vdd DFFPOSX1
XNAND2X1_1022 DFFPOSX1_214/Q INVX4_14/A gnd NAND3X1_359/A vdd NAND2X1
XDFFPOSX1_77 AOI22X1_39/A CLKBUF1_31/Y INVX1_130/A gnd vdd DFFPOSX1
XDFFPOSX1_55 AOI22X1_17/A CLKBUF1_63/Y INVX1_108/A gnd vdd DFFPOSX1
XDFFPOSX1_66 AOI22X1_28/A CLKBUF1_51/Y INVX1_119/A gnd vdd DFFPOSX1
XDFFPOSX1_88 INVX1_201/A CLKBUF1_18/Y OAI21X1_117/C gnd vdd DFFPOSX1
XDFFPOSX1_99 INVX1_212/A CLKBUF1_19/Y OAI21X1_139/C gnd vdd DFFPOSX1
XFILL_28_5_1 gnd vdd FILL
XFILL_3_5_1 gnd vdd FILL
XFILL_2_0_0 gnd vdd FILL
XFILL_27_0_0 gnd vdd FILL
XNAND3X1_305 BUFX4_123/Y NAND3X1_305/B NAND3X1_305/C gnd NAND2X1_887/B vdd NAND3X1
XNAND3X1_338 AOI21X1_245/A AND2X2_93/Y OAI21X1_925/Y gnd NAND3X1_343/C vdd NAND3X1
XNAND3X1_327 NAND2X1_926/Y OAI21X1_882/Y NAND3X1_327/C gnd NAND3X1_327/Y vdd NAND3X1
XNAND3X1_316 INVX1_633/Y BUFX4_101/Y BUFX4_164/Y gnd NAND3X1_316/Y vdd NAND3X1
XNAND3X1_349 NAND3X1_349/A INVX2_93/A OAI22X1_58/C gnd BUFX2_37/A vdd NAND3X1
XFILL_11_4_1 gnd vdd FILL
XFILL_19_5_1 gnd vdd FILL
XFILL_18_0_0 gnd vdd FILL
XDFFPOSX1_404 OR2X2_53/B CLKBUF1_37/Y OAI21X1_61/Y gnd vdd DFFPOSX1
XDFFPOSX1_437 BUFX2_96/A CLKBUF1_44/Y NOR3X1_44/Y gnd vdd DFFPOSX1
XDFFPOSX1_415 NOR2X1_22/B CLKBUF1_34/Y NOR3X1_22/Y gnd vdd DFFPOSX1
XDFFPOSX1_426 INVX2_74/A CLKBUF1_9/Y NOR3X1_33/Y gnd vdd DFFPOSX1
XDFFPOSX1_448 NAND3X1_22/A CLKBUF1_7/Y BUFX2_47/A gnd vdd DFFPOSX1
XDFFPOSX1_459 NAND3X1_44/A CLKBUF1_45/Y BUFX2_58/A gnd vdd DFFPOSX1
XINVX1_160 instruction_memory_interface_data[4] gnd INVX1_160/Y vdd INVX1
XNAND2X1_518 INVX2_39/Y MUX2X1_37/B gnd AOI22X1_99/D vdd NAND2X1
XNAND2X1_507 NOR2X1_277/Y NOR3X1_56/Y gnd NAND3X1_134/B vdd NAND2X1
XINVX1_182 instruction_memory_interface_data[26] gnd INVX1_182/Y vdd INVX1
XINVX1_193 INVX1_193/A gnd INVX1_193/Y vdd INVX1
XINVX1_171 instruction_memory_interface_data[15] gnd INVX1_171/Y vdd INVX1
XNAND2X1_529 BUFX4_84/Y MUX2X1_38/Y gnd OAI21X1_779/A vdd NAND2X1
XAOI21X1_131 INVX1_399/A OAI21X1_694/A BUFX4_275/Y gnd AOI21X1_131/Y vdd AOI21X1
XAOI21X1_142 AOI22X1_71/B OAI22X1_9/C OAI22X1_9/B gnd OAI21X1_601/C vdd AOI21X1
XAOI21X1_120 BUFX4_43/Y MUX2X1_37/A NOR2X1_192/Y gnd MUX2X1_36/A vdd AOI21X1
XAOI21X1_164 BUFX4_51/Y NOR2X1_328/B AOI21X1_164/C gnd OAI21X1_665/A vdd AOI21X1
XAOI21X1_153 AOI21X1_153/A BUFX4_190/Y OAI22X1_39/Y gnd AOI21X1_153/Y vdd AOI21X1
XAOI21X1_175 AND2X2_59/A INVX1_412/Y INVX1_414/Y gnd INVX1_418/A vdd AOI21X1
XAOI21X1_186 INVX2_33/Y OAI21X1_646/Y AOI21X1_186/C gnd AOI21X1_186/Y vdd AOI21X1
XAOI21X1_197 INVX4_7/Y OR2X2_42/A OR2X2_41/Y gnd NOR2X1_352/A vdd AOI21X1
XFILL_43_3_1 gnd vdd FILL
XNAND3X1_113 BUFX4_80/Y BUFX4_83/Y INVX1_371/A gnd OR2X2_42/A vdd NAND3X1
XNAND3X1_102 NAND3X1_101/Y OAI21X1_371/Y NAND3X1_102/C gnd NOR2X1_178/A vdd NAND3X1
XNAND3X1_124 AOI22X1_91/Y AOI22X1_92/Y NOR2X1_250/Y gnd INVX1_75/A vdd NAND3X1
XNAND3X1_135 NAND3X1_132/Y OAI21X1_555/Y NAND3X1_135/C gnd INVX1_78/A vdd NAND3X1
XNAND3X1_146 AOI21X1_37/B INVX1_402/A NAND3X1_146/C gnd NAND3X1_147/B vdd NAND3X1
XNAND3X1_157 NAND3X1_157/A NAND3X1_155/Y NOR3X1_61/Y gnd INVX1_89/A vdd NAND3X1
XNAND3X1_179 BUFX2_41/A BUFX2_42/A BUFX2_43/A gnd INVX1_471/A vdd NAND3X1
XNAND3X1_168 OR2X2_42/Y NOR2X1_361/Y OAI21X1_748/Y gnd AOI21X1_201/C vdd NAND3X1
XFILL_34_3_1 gnd vdd FILL
XFILL_20_2 gnd vdd FILL
XOAI21X1_309 INVX1_332/Y INVX4_4/A OAI21X1_309/C gnd MUX2X1_35/B vdd OAI21X1
XBUFX4_7 CLK gnd BUFX4_7/Y vdd BUFX4
XDFFPOSX1_201 INVX1_729/A CLKBUF1_28/Y OR2X2_58/B gnd vdd DFFPOSX1
XDFFPOSX1_212 INVX1_724/A CLKBUF1_29/Y INVX1_458/A gnd vdd DFFPOSX1
XDFFPOSX1_234 OAI21X1_121/C CLKBUF1_57/Y INVX1_78/A gnd vdd DFFPOSX1
XDFFPOSX1_245 OAI21X1_143/C CLKBUF1_63/Y INVX1_89/A gnd vdd DFFPOSX1
XDFFPOSX1_223 OAI21X1_99/C CLKBUF1_23/Y INVX1_67/A gnd vdd DFFPOSX1
XDFFPOSX1_256 INVX1_351/A CLKBUF1_52/Y NAND3X1_10/A gnd vdd DFFPOSX1
XDFFPOSX1_267 MUX2X1_6/A CLKBUF1_14/Y NAND3X1_32/A gnd vdd DFFPOSX1
XDFFPOSX1_278 AOI22X1_61/A CLKBUF1_17/Y NAND3X1_54/A gnd vdd DFFPOSX1
XDFFPOSX1_289 NOR2X1_1/A CLKBUF1_13/Y NOR3X1_13/Y gnd vdd DFFPOSX1
XNAND2X1_326 INVX8_5/A AOI21X1_51/Y gnd NAND2X1_326/Y vdd NAND2X1
XNAND2X1_304 INVX2_41/Y MUX2X1_37/A gnd OAI21X1_606/C vdd NAND2X1
XNAND2X1_315 INVX2_48/Y INVX1_390/A gnd NOR2X1_135/A vdd NAND2X1
XNAND2X1_337 INVX8_3/A AND2X2_38/A gnd OAI21X1_367/C vdd NAND2X1
XNAND2X1_359 BUFX4_124/Y NOR2X1_186/Y gnd OR2X2_29/B vdd NAND2X1
XNAND2X1_348 INVX1_390/A AND2X2_25/A gnd NOR2X1_175/B vdd NAND2X1
XNOR3X1_44 NOR3X1_3/A INVX1_185/Y BUFX4_49/Y gnd NOR3X1_44/Y vdd NOR3X1
XNOR3X1_11 NOR3X1_4/A INVX1_148/Y NOR3X1_4/C gnd NOR3X1_11/Y vdd NOR3X1
XNOR3X1_22 INVX4_1/A INVX1_163/Y BUFX4_45/Y gnd NOR3X1_22/Y vdd NOR3X1
XNOR3X1_33 NOR3X1_35/A INVX1_174/Y BUFX4_48/Y gnd NOR3X1_33/Y vdd NOR3X1
XNOR3X1_66 NOR3X1_66/A NOR3X1_66/B NOR3X1_66/C gnd NOR3X1_66/Y vdd NOR3X1
XNOR3X1_55 XNOR2X1_8/Y XNOR2X1_9/Y AOI21X1_6/Y gnd NOR3X1_55/Y vdd NOR3X1
XNOR3X1_77 NOR3X1_78/C INVX2_90/Y NOR3X1_79/A gnd NOR3X1_77/Y vdd NOR3X1
XFILL_25_3_1 gnd vdd FILL
XFILL_0_3_1 gnd vdd FILL
XNOR2X1_370 BUFX4_276/Y NOR2X1_370/B gnd NOR2X1_370/Y vdd NOR2X1
XNOR2X1_381 BUFX2_43/A OR2X2_45/A gnd NOR2X1_381/Y vdd NOR2X1
XNOR2X1_392 BUFX2_61/A NOR2X1_392/B gnd NOR2X1_392/Y vdd NOR2X1
XINVX4_7 INVX4_7/A gnd INVX4_7/Y vdd INVX4
XOAI21X1_821 OAI21X1_820/Y INVX1_470/Y OAI21X1_821/C gnd OAI21X1_821/Y vdd OAI21X1
XOAI21X1_832 OAI21X1_831/Y OR2X2_45/B OAI21X1_832/C gnd OAI21X1_832/Y vdd OAI21X1
XOAI21X1_810 BUFX4_178/Y INVX1_463/Y NAND2X1_633/Y gnd OAI21X1_810/Y vdd OAI21X1
XOAI21X1_876 INVX2_77/Y DFFPOSX1_43/Q DFFPOSX1_45/Q gnd NOR2X1_410/A vdd OAI21X1
XOAI21X1_843 OAI21X1_843/A OR2X2_45/B OAI21X1_843/C gnd OAI21X1_178/C vdd OAI21X1
XOAI21X1_854 OAI21X1_853/Y NOR2X1_392/Y OAI21X1_854/C gnd OAI21X1_854/Y vdd OAI21X1
XOAI21X1_865 OAI21X1_864/Y BUFX4_241/Y OAI21X1_865/C gnd OAI21X1_865/Y vdd OAI21X1
XOAI21X1_898 INVX8_14/Y AOI21X1_231/Y AOI22X1_122/Y gnd OAI21X1_898/Y vdd OAI21X1
XOAI21X1_887 INVX1_658/Y OAI21X1_887/B INVX4_11/Y gnd OAI21X1_887/Y vdd OAI21X1
XFILL_8_4_1 gnd vdd FILL
XNAND2X1_882 OAI21X1_86/Y BUFX4_59/Y gnd NAND2X1_882/Y vdd NAND2X1
XNAND2X1_860 NAND2X1_858/Y NAND2X1_860/B gnd NAND2X1_46/B vdd NAND2X1
XNAND2X1_871 INVX1_610/Y BUFX4_95/Y gnd NAND2X1_871/Y vdd NAND2X1
XNAND2X1_893 NAND2X1_891/Y NAND2X1_893/B gnd NAND2X1_57/B vdd NAND2X1
XFILL_16_3_1 gnd vdd FILL
XOAI21X1_117 BUFX4_272/Y BUFX4_195/Y OAI21X1_117/C gnd OAI21X1_118/C vdd OAI21X1
XOAI21X1_128 BUFX4_183/Y INVX1_114/Y OAI21X1_128/C gnd INVX1_607/A vdd OAI21X1
XOAI21X1_106 BUFX4_182/Y INVX1_103/Y OAI21X1_106/C gnd INVX1_585/A vdd OAI21X1
XOAI21X1_139 BUFX4_270/Y OR2X2_2/B OAI21X1_139/C gnd OAI21X1_139/Y vdd OAI21X1
XBUFX2_4 BUFX2_4/A gnd data_memory_interface_address[3] vdd BUFX2
XNAND2X1_101 AND2X2_4/B AND2X2_4/A gnd OAI22X1_1/C vdd NAND2X1
XNAND2X1_134 NAND3X1_81/Y AOI21X1_13/B gnd INVX1_248/A vdd NAND2X1
XNAND2X1_123 OR2X2_61/A BUFX4_146/Y gnd NAND3X1_79/C vdd NAND2X1
XNAND2X1_112 NOR2X1_17/Y NOR2X1_16/Y gnd NAND2X1_112/Y vdd NAND2X1
XNAND2X1_145 NOR2X1_34/Y NOR2X1_33/Y gnd NOR2X1_48/A vdd NAND2X1
XNAND2X1_178 AOI21X1_28/C NOR2X1_49/Y gnd AND2X2_16/A vdd NAND2X1
XNAND2X1_156 XNOR2X1_37/Y XNOR2X1_38/Y gnd NOR2X1_42/B vdd NAND2X1
XNAND2X1_167 OR2X2_12/B OR2X2_12/A gnd NAND2X1_168/A vdd NAND2X1
XNAND2X1_189 NOR2X1_62/A INVX1_291/Y gnd INVX1_292/A vdd NAND2X1
XFILL_40_1_1 gnd vdd FILL
XINVX2_4 INVX2_4/A gnd OR2X2_6/B vdd INVX2
XOAI21X1_640 NOR2X1_317/Y NOR2X1_94/Y NOR2X1_320/Y gnd OAI21X1_640/Y vdd OAI21X1
XOAI21X1_651 NOR2X1_323/Y NOR2X1_322/Y BUFX4_129/Y gnd AOI21X1_160/A vdd OAI21X1
XOAI21X1_673 BUFX4_55/Y AOI22X1_98/C AND2X2_56/Y gnd AOI21X1_170/B vdd OAI21X1
XOAI21X1_662 OAI21X1_662/A BUFX4_228/Y NAND2X1_557/Y gnd MUX2X1_49/B vdd OAI21X1
XAOI21X1_4 AOI21X1_4/A AOI21X1_4/B AOI21X1_4/C gnd BUFX4_233/A vdd AOI21X1
XOAI21X1_684 NOR2X1_332/Y NOR2X1_99/Y OR2X2_38/A gnd NAND3X1_155/B vdd OAI21X1
XOAI21X1_695 NOR2X1_81/Y AOI21X1_200/B OAI21X1_695/C gnd NAND3X1_159/A vdd OAI21X1
XINVX1_704 OR2X2_53/A gnd INVX1_704/Y vdd INVX1
XINVX1_726 INVX1_726/A gnd INVX1_726/Y vdd INVX1
XINVX1_715 INVX1_715/A gnd NOR3X1_76/A vdd INVX1
XINVX1_748 data_memory_interface_data[12] gnd INVX1_748/Y vdd INVX1
XINVX1_759 INVX1_759/A gnd INVX1_759/Y vdd INVX1
XINVX1_737 data_memory_interface_data[1] gnd INVX1_737/Y vdd INVX1
XXNOR2X1_23 NOR2X1_31/B INVX2_9/A gnd AOI21X1_17/A vdd XNOR2X1
XXNOR2X1_12 INVX1_240/A NOR2X1_29/A gnd XNOR2X1_12/Y vdd XNOR2X1
XXNOR2X1_34 NOR2X1_40/B INVX2_13/A gnd XNOR2X1_34/Y vdd XNOR2X1
XXNOR2X1_45 XNOR2X1_45/A NOR2X1_54/B gnd XNOR2X1_45/Y vdd XNOR2X1
XNAND2X1_690 BUFX2_65/A BUFX2_66/A gnd INVX1_491/A vdd NAND2X1
XBUFX2_11 BUFX2_11/A gnd data_memory_interface_address[10] vdd BUFX2
XINVX1_91 INVX1_91/A gnd INVX1_91/Y vdd INVX1
XINVX1_80 INVX1_80/A gnd INVX1_80/Y vdd INVX1
XBUFX2_33 BUFX2_33/A gnd data_memory_interface_enable vdd BUFX2
XBUFX2_44 BUFX2_44/A gnd instruction_memory_interface_address[5] vdd BUFX2
XBUFX2_22 BUFX2_22/A gnd data_memory_interface_address[21] vdd BUFX2
XBUFX2_55 BUFX2_55/A gnd instruction_memory_interface_address[16] vdd BUFX2
XBUFX2_66 BUFX2_66/A gnd instruction_memory_interface_address[27] vdd BUFX2
XBUFX2_77 BUFX2_77/A gnd BUFX2_77/Y vdd BUFX2
XBUFX2_99 INVX8_14/A gnd BUFX2_99/Y vdd BUFX2
XBUFX2_88 INVX2_76/A gnd BUFX2_88/Y vdd BUFX2
XFILL_31_1_1 gnd vdd FILL
XNOR2X1_2 OR2X2_1/Y NOR2X1_2/B gnd NOR2X1_2/Y vdd NOR2X1
XFILL_39_2_1 gnd vdd FILL
XFILL_22_1_1 gnd vdd FILL
XAOI21X1_23 NOR2X1_36/A NOR2X1_39/Y INVX1_263/A gnd AOI21X1_29/A vdd AOI21X1
XAOI21X1_12 AOI21X1_8/A AOI21X1_8/B INVX1_250/Y gnd AOI21X1_12/Y vdd AOI21X1
XAOI21X1_34 AOI21X1_33/Y AOI21X1_34/B INVX1_287/A gnd AOI21X1_34/Y vdd AOI21X1
XAOI21X1_67 INVX8_3/A NOR2X1_270/B INVX8_7/A gnd AOI21X1_67/Y vdd AOI21X1
XAOI21X1_56 AOI21X1_56/A BUFX4_152/Y AOI21X1_56/C gnd AOI21X1_56/Y vdd AOI21X1
XAOI21X1_45 INVX2_28/Y AOI21X1_45/B AOI21X1_45/C gnd AOI21X1_45/Y vdd AOI21X1
XAOI21X1_78 AOI22X1_81/B AOI21X1_78/B NOR2X1_110/Y gnd AOI21X1_78/Y vdd AOI21X1
XAOI21X1_89 AOI21X1_89/A AOI21X1_89/B AOI21X1_89/C gnd AOI21X1_89/Y vdd AOI21X1
XOAI21X1_7 INVX1_7/Y BUFX4_24/Y OAI21X1_7/C gnd OAI21X1_7/Y vdd OAI21X1
XFILL_5_2_1 gnd vdd FILL
XOAI22X1_20 OAI22X1_20/A AND2X2_36/A INVX4_8/Y OAI22X1_43/B gnd AOI21X1_94/C vdd OAI22X1
XOAI22X1_31 OAI22X1_31/A OAI22X1_31/B OAI22X1_31/C NOR2X1_285/Y gnd NOR2X1_304/A vdd
+ OAI22X1
XFILL_13_1_1 gnd vdd FILL
XOAI22X1_42 AND2X2_70/Y OAI22X1_42/B MUX2X1_49/A MUX2X1_49/S gnd OAI22X1_42/Y vdd
+ OAI22X1
XOAI22X1_53 INVX2_91/Y OAI22X1_58/B OAI22X1_58/C INVX1_735/Y gnd OAI22X1_53/Y vdd
+ OAI22X1
XOAI21X1_470 OAI21X1_470/A INVX8_5/A OAI21X1_470/C gnd NAND2X1_438/B vdd OAI21X1
XOAI21X1_481 OAI21X1_416/A BUFX4_215/Y NAND2X1_454/Y gnd NOR2X1_225/B vdd OAI21X1
XOAI21X1_492 AOI22X1_86/A OAI22X1_11/A NOR2X1_232/Y gnd NAND3X1_117/C vdd OAI21X1
XINVX1_501 INVX1_501/A gnd INVX1_501/Y vdd INVX1
XINVX1_534 INVX1_607/A gnd INVX1_534/Y vdd INVX1
XINVX1_512 INVX1_585/A gnd INVX1_512/Y vdd INVX1
XINVX1_523 INVX1_523/A gnd INVX1_523/Y vdd INVX1
XINVX1_545 INVX1_545/A gnd INVX1_545/Y vdd INVX1
XINVX1_578 INVX1_578/A gnd INVX1_578/Y vdd INVX1
XINVX1_567 INVX1_640/A gnd INVX1_567/Y vdd INVX1
XINVX1_556 INVX1_556/A gnd INVX1_556/Y vdd INVX1
XINVX1_589 INVX1_589/A gnd INVX1_589/Y vdd INVX1
XAOI22X1_100 INVX1_329/Y BUFX4_154/Y OR2X2_24/Y INVX1_399/Y gnd AOI22X1_100/Y vdd
+ AOI22X1
XAOI22X1_111 INVX1_501/Y INVX2_73/A INVX1_502/A INVX2_74/Y gnd NAND2X1_710/B vdd AOI22X1
XAOI22X1_144 data_memory_interface_data[7] BUFX4_105/Y AOI22X1_144/C BUFX4_8/Y gnd
+ AOI22X1_144/Y vdd AOI22X1
XAOI22X1_155 data_memory_interface_data[19] BUFX4_108/Y BUFX4_170/Y BUFX4_250/Y gnd
+ AOI22X1_155/Y vdd AOI22X1
XAOI22X1_133 INVX1_685/Y INVX1_435/A OR2X2_64/Y NAND2X1_959/Y gnd AOI22X1_133/Y vdd
+ AOI22X1
XAOI22X1_122 OAI22X1_49/A INVX4_11/A BUFX4_263/Y BUFX2_94/A gnd AOI22X1_122/Y vdd
+ AOI22X1
XBUFX4_117 BUFX4_118/A gnd BUFX4_117/Y vdd BUFX4
XBUFX4_128 INVX8_7/Y gnd BUFX4_128/Y vdd BUFX4
XBUFX4_106 BUFX4_107/A gnd BUFX4_106/Y vdd BUFX4
XAOI22X1_166 data_memory_interface_data[30] INVX4_14/A BUFX4_169/Y BUFX4_253/Y gnd
+ AOI22X1_166/Y vdd AOI22X1
XBUFX4_139 OAI22X1_1/Y gnd BUFX4_139/Y vdd BUFX4
XOAI21X1_1018 BUFX4_65/Y BUFX4_69/Y AOI22X1_145/Y gnd OAI21X1_1018/Y vdd OAI21X1
XOAI21X1_1007 NOR3X1_77/Y NOR3X1_78/Y INVX8_16/A gnd OAI21X1_1007/Y vdd OAI21X1
XOAI21X1_1029 INVX1_751/Y INVX2_93/A OAI21X1_1029/C gnd AOI22X1_149/C vdd OAI21X1
XINVX1_342 INVX1_342/A gnd INVX1_342/Y vdd INVX1
XINVX1_331 MUX2X1_4/B gnd INVX1_331/Y vdd INVX1
XINVX1_353 INVX1_353/A gnd INVX1_353/Y vdd INVX1
XINVX1_320 INVX1_672/A gnd INVX1_320/Y vdd INVX1
XINVX1_375 INVX1_375/A gnd INVX1_375/Y vdd INVX1
XINVX1_386 MUX2X1_30/Y gnd INVX1_386/Y vdd INVX1
XINVX1_364 INVX1_364/A gnd INVX1_364/Y vdd INVX1
XINVX1_397 INVX1_397/A gnd INVX1_397/Y vdd INVX1
XFILL_1_1 gnd vdd FILL
XFILL_43_1 gnd vdd FILL
XFILL_36_0_1 gnd vdd FILL
XNAND2X1_1001 OAI21X1_966/C OAI21X1_951/Y gnd OAI21X1_952/C vdd NAND2X1
XDFFPOSX1_45 DFFPOSX1_45/Q CLKBUF1_43/Y INVX1_504/A gnd vdd DFFPOSX1
XDFFPOSX1_23 AOI22X1_23/D CLKBUF1_50/Y DFFPOSX1_23/D gnd vdd DFFPOSX1
XDFFPOSX1_34 AOI22X1_34/D CLKBUF1_24/Y DFFPOSX1_34/D gnd vdd DFFPOSX1
XDFFPOSX1_12 AOI22X1_12/D CLKBUF1_55/Y DFFPOSX1_12/D gnd vdd DFFPOSX1
XNAND2X1_1023 INVX1_726/A BUFX4_252/Y gnd NAND3X1_359/B vdd NAND2X1
XNAND2X1_1012 data_memory_interface_data[1] OAI21X1_993/B gnd OAI21X1_985/C vdd NAND2X1
XDFFPOSX1_56 AOI22X1_18/A CLKBUF1_18/Y INVX1_109/A gnd vdd DFFPOSX1
XDFFPOSX1_78 INVX1_188/A CLKBUF1_21/Y OAI21X1_97/C gnd vdd DFFPOSX1
XDFFPOSX1_67 AOI22X1_29/A CLKBUF1_61/Y INVX1_120/A gnd vdd DFFPOSX1
XDFFPOSX1_89 INVX1_202/A CLKBUF1_61/Y OAI21X1_119/C gnd vdd DFFPOSX1
XFILL_2_0_1 gnd vdd FILL
XFILL_27_0_1 gnd vdd FILL
XNAND3X1_306 INVX1_623/Y BUFX4_102/Y BUFX4_168/Y gnd NAND3X1_306/Y vdd NAND3X1
XNAND3X1_328 NOR2X1_6/A OR2X2_1/B INVX1_663/Y gnd NAND3X1_328/Y vdd NAND3X1
XNAND3X1_339 NAND2X1_991/Y AOI22X1_133/Y OAI21X1_907/C gnd OR2X2_68/B vdd NAND3X1
XNAND3X1_317 BUFX4_119/Y NAND3X1_316/Y NAND2X1_904/Y gnd NAND2X1_905/B vdd NAND3X1
XFILL_18_0_1 gnd vdd FILL
XFILL_30_7_0 gnd vdd FILL
XDFFPOSX1_427 OR2X2_49/B CLKBUF1_39/Y NOR3X1_34/Y gnd vdd DFFPOSX1
XDFFPOSX1_438 BUFX2_97/A CLKBUF1_44/Y NOR3X1_45/Y gnd vdd DFFPOSX1
XDFFPOSX1_405 INVX2_80/A CLKBUF1_22/Y OAI21X1_62/Y gnd vdd DFFPOSX1
XDFFPOSX1_416 NOR2X1_22/A CLKBUF1_9/Y NOR3X1_23/Y gnd vdd DFFPOSX1
XDFFPOSX1_449 NAND3X1_24/A CLKBUF1_33/Y XOR2X1_8/B gnd vdd DFFPOSX1
XINVX1_150 INVX1_150/A gnd INVX1_150/Y vdd INVX1
XINVX1_161 instruction_memory_interface_data[5] gnd INVX1_161/Y vdd INVX1
XNAND2X1_508 INVX8_3/A MUX2X1_26/Y gnd OAI21X1_558/C vdd NAND2X1
XINVX1_183 instruction_memory_interface_data[27] gnd INVX1_183/Y vdd INVX1
XINVX1_194 INVX1_194/A gnd INVX1_194/Y vdd INVX1
XINVX1_172 instruction_memory_interface_data[16] gnd INVX1_172/Y vdd INVX1
XNAND2X1_519 AOI22X1_99/C AOI22X1_99/D gnd INVX2_63/A vdd NAND2X1
XFILL_21_7_0 gnd vdd FILL
XAOI21X1_110 INVX2_60/Y AOI21X1_110/B OAI21X1_547/Y gnd NAND3X1_131/C vdd AOI21X1
XAOI21X1_132 AOI22X1_96/B NOR2X1_269/A OAI22X1_37/B gnd AOI21X1_132/Y vdd AOI21X1
XAOI21X1_121 OAI21X1_330/C OAI22X1_31/B NOR2X1_285/Y gnd OAI21X1_593/B vdd AOI21X1
XAOI21X1_154 NOR3X1_56/Y AOI21X1_154/B OR2X2_37/Y gnd NAND3X1_149/C vdd AOI21X1
XAOI21X1_143 AOI22X1_70/B OAI22X1_7/C OAI22X1_7/B gnd AOI21X1_143/Y vdd AOI21X1
XAOI21X1_165 INVX1_379/Y AOI21X1_89/A AOI21X1_165/C gnd AOI21X1_165/Y vdd AOI21X1
XAOI21X1_176 INVX1_405/Y NOR2X1_336/Y AOI21X1_176/C gnd AOI21X1_176/Y vdd AOI21X1
XAOI21X1_198 INVX2_65/A OAI22X1_40/Y AOI21X1_198/C gnd AOI21X1_198/Y vdd AOI21X1
XAOI21X1_187 AND2X2_65/Y OAI21X1_732/A AOI21X1_187/C gnd AOI21X1_190/B vdd AOI21X1
XNAND3X1_114 NAND3X1_114/A AOI21X1_82/Y NAND3X1_114/C gnd AOI21X1_83/C vdd NAND3X1
XNAND3X1_103 NOR2X1_203/B OR2X2_23/Y INVX8_11/A gnd NOR3X1_56/A vdd NAND3X1
XNAND3X1_147 INVX8_11/Y NAND3X1_147/B OAI21X1_630/Y gnd NAND3X1_147/Y vdd NAND3X1
XNAND3X1_136 OAI21X1_563/Y OAI21X1_565/Y NOR2X1_284/Y gnd INVX1_79/A vdd NAND3X1
XNAND3X1_125 INVX2_48/Y INVX1_355/A NOR2X1_257/Y gnd OR2X2_31/B vdd NAND3X1
XFILL_12_7_0 gnd vdd FILL
XNAND3X1_158 NAND3X1_158/A NAND3X1_158/B NAND2X1_575/Y gnd NOR3X1_62/B vdd NAND3X1
XNAND3X1_169 NAND3X1_169/A NAND3X1_169/B AOI21X1_201/Y gnd INVX1_94/A vdd NAND3X1
XDFFPOSX1_202 INVX1_730/A CLKBUF1_28/Y OR2X2_57/B gnd vdd DFFPOSX1
XDFFPOSX1_213 INVX1_725/A CLKBUF1_38/Y INVX1_459/A gnd vdd DFFPOSX1
XDFFPOSX1_235 OAI21X1_123/C CLKBUF1_53/Y INVX1_79/A gnd vdd DFFPOSX1
XDFFPOSX1_224 OAI21X1_101/C CLKBUF1_15/Y INVX1_68/A gnd vdd DFFPOSX1
XDFFPOSX1_246 OAI21X1_145/C CLKBUF1_63/Y INVX1_90/A gnd vdd DFFPOSX1
XBUFX4_8 BUFX4_9/A gnd BUFX4_8/Y vdd BUFX4
XDFFPOSX1_257 INVX1_350/A CLKBUF1_54/Y NAND3X1_12/A gnd vdd DFFPOSX1
XDFFPOSX1_268 MUX2X1_4/A CLKBUF1_14/Y NAND3X1_34/A gnd vdd DFFPOSX1
XDFFPOSX1_279 AOI22X1_62/A CLKBUF1_17/Y NAND3X1_56/A gnd vdd DFFPOSX1
XNAND2X1_327 INVX8_4/A INVX1_375/A gnd NAND2X1_327/Y vdd NAND2X1
XNAND2X1_305 OAI21X1_330/C OAI21X1_606/C gnd NOR2X1_281/A vdd NAND2X1
XNAND2X1_316 INVX2_23/Y INVX2_24/A gnd INVX1_428/A vdd NAND2X1
XNAND2X1_349 INVX1_355/A NOR2X1_175/Y gnd OR2X2_22/A vdd NAND2X1
XNAND2X1_338 INVX8_8/A NOR2X1_332/B gnd NAND2X1_338/Y vdd NAND2X1
XNOR3X1_34 NOR3X1_35/A INVX1_175/Y BUFX4_48/Y gnd NOR3X1_34/Y vdd NOR3X1
XNOR3X1_12 INVX4_1/A NOR3X1_12/B BUFX4_45/Y gnd NOR3X1_12/Y vdd NOR3X1
XNOR3X1_23 NOR3X1_35/A INVX1_164/Y BUFX4_48/Y gnd NOR3X1_23/Y vdd NOR3X1
XNOR3X1_67 NOR3X1_66/A NOR3X1_67/B NOR3X1_66/C gnd NOR3X1_67/Y vdd NOR3X1
XNOR3X1_56 NOR3X1_56/A INVX1_394/A NOR3X1_56/C gnd NOR3X1_56/Y vdd NOR3X1
XNOR3X1_45 NOR3X1_3/A INVX1_186/Y BUFX4_49/Y gnd NOR3X1_45/Y vdd NOR3X1
XNOR3X1_78 INVX2_90/Y NOR3X1_80/A NOR3X1_78/C gnd NOR3X1_78/Y vdd NOR3X1
XNOR2X1_360 AND2X2_56/B OR2X2_33/A gnd NOR2X1_360/Y vdd NOR2X1
XNOR2X1_382 INVX1_471/A NOR2X1_382/B gnd NOR2X1_382/Y vdd NOR2X1
XNOR2X1_393 OR2X2_48/B NOR2X1_393/B gnd AND2X2_78/B vdd NOR2X1
XNOR2X1_371 MUX2X1_45/Y INVX4_9/Y gnd NOR2X1_371/Y vdd NOR2X1
XINVX4_8 INVX4_8/A gnd INVX4_8/Y vdd INVX4
XOAI21X1_800 BUFX4_181/Y INVX1_453/Y NAND2X1_623/Y gnd OAI21X1_800/Y vdd OAI21X1
XOAI21X1_822 XNOR2X1_50/Y OR2X2_45/B OAI21X1_822/C gnd OAI21X1_167/C vdd OAI21X1
XOAI21X1_833 NOR2X1_385/Y OAI21X1_833/B NAND2X1_659/Y gnd OAI21X1_173/C vdd OAI21X1
XOAI21X1_811 BUFX4_178/Y INVX1_464/Y NAND2X1_634/Y gnd OAI21X1_811/Y vdd OAI21X1
XOAI21X1_844 OAI21X1_846/A INVX1_481/Y INVX8_13/Y gnd OAI21X1_844/Y vdd OAI21X1
XOAI21X1_855 NOR3X1_66/C NOR3X1_66/A INVX8_13/Y gnd OAI21X1_855/Y vdd OAI21X1
XOAI21X1_866 NAND2X1_695/Y OAI21X1_866/B OAI21X1_866/C gnd OAI21X1_866/Y vdd OAI21X1
XOAI21X1_899 INVX8_14/Y AOI21X1_231/Y AOI22X1_123/Y gnd OAI21X1_899/Y vdd OAI21X1
XOAI21X1_877 OAI21X1_877/A INVX1_644/Y NAND2X1_921/Y gnd OAI21X1_877/Y vdd OAI21X1
XOAI21X1_888 INVX1_659/Y OAI21X1_887/B INVX4_11/Y gnd OAI21X1_888/Y vdd OAI21X1
XNAND2X1_872 NAND2X1_870/Y NAND2X1_872/B gnd NAND2X1_50/B vdd NAND2X1
XNAND2X1_861 OAI21X1_79/Y BUFX4_60/Y gnd NAND2X1_861/Y vdd NAND2X1
XNAND2X1_850 INVX1_596/Y BUFX4_94/Y gnd NAND3X1_281/C vdd NAND2X1
XNAND2X1_894 OAI21X1_90/Y BUFX4_60/Y gnd NAND2X1_896/A vdd NAND2X1
XNAND2X1_883 INVX1_618/Y BUFX4_96/Y gnd NAND2X1_883/Y vdd NAND2X1
XFILL_35_6_0 gnd vdd FILL
XOAI21X1_118 BUFX4_183/Y INVX1_109/Y OAI21X1_118/C gnd INVX1_524/A vdd OAI21X1
XOAI21X1_129 BUFX4_270/Y OR2X2_2/B OAI21X1_129/C gnd OAI21X1_130/C vdd OAI21X1
XOAI21X1_107 OR2X2_2/A BUFX4_194/Y DFFPOSX1_83/D gnd OAI21X1_107/Y vdd OAI21X1
XBUFX2_5 BUFX2_5/A gnd data_memory_interface_address[4] vdd BUFX2
XNAND2X1_135 INVX1_689/A BUFX4_147/Y gnd NAND3X1_82/C vdd NAND2X1
XNAND2X1_124 INVX1_239/A BUFX4_232/Y gnd NAND3X1_79/B vdd NAND2X1
XNAND2X1_102 NOR2X1_5/Y AND2X2_1/Y gnd NOR2X1_7/A vdd NAND2X1
XNAND2X1_113 NOR2X1_14/A INVX1_227/Y gnd NAND3X1_74/B vdd NAND2X1
XNAND2X1_157 NOR2X1_36/A NOR2X1_39/Y gnd NAND2X1_158/B vdd NAND2X1
XNAND2X1_146 INVX1_258/Y AOI21X1_20/Y gnd NAND3X1_83/B vdd NAND2X1
XNAND2X1_168 NAND2X1_168/A OR2X2_12/Y gnd NOR2X1_45/A vdd NAND2X1
XNAND2X1_179 INVX1_278/Y NOR2X1_52/B gnd NAND2X1_180/A vdd NAND2X1
XFILL_26_6_0 gnd vdd FILL
XFILL_1_6_0 gnd vdd FILL
XNOR2X1_190 BUFX4_40/Y INVX2_27/Y gnd OR2X2_25/B vdd NOR2X1
XINVX2_5 INVX2_5/A gnd INVX2_5/Y vdd INVX2
XOAI21X1_630 NOR2X1_317/Y NOR2X1_94/Y OAI21X1_630/C gnd OAI21X1_630/Y vdd OAI21X1
XOAI21X1_641 NOR2X1_312/Y INVX1_329/A INVX2_68/A gnd OAI21X1_641/Y vdd OAI21X1
XOAI21X1_663 OAI21X1_663/A NOR2X1_327/Y INVX2_65/A gnd NAND3X1_152/A vdd OAI21X1
XOAI21X1_652 MUX2X1_54/B INVX8_3/A OAI21X1_652/C gnd OAI21X1_653/C vdd OAI21X1
XOAI21X1_674 NOR2X1_330/Y NOR2X1_329/Y BUFX4_128/Y gnd OAI21X1_675/C vdd OAI21X1
XAOI21X1_5 AOI21X1_5/A AOI21X1_5/B INVX1_230/Y gnd AOI21X1_5/Y vdd AOI21X1
XOAI21X1_685 INVX1_404/A BUFX4_217/Y OAI21X1_685/C gnd MUX2X1_56/B vdd OAI21X1
XOAI21X1_696 NOR2X1_98/Y INVX1_401/A INVX1_326/Y gnd OAI21X1_696/Y vdd OAI21X1
XINVX1_705 INVX1_705/A gnd INVX1_705/Y vdd INVX1
XINVX1_727 INVX1_727/A gnd INVX1_727/Y vdd INVX1
XINVX1_716 NOR2X1_3/B gnd INVX1_716/Y vdd INVX1
XINVX1_749 data_memory_interface_data[5] gnd INVX1_749/Y vdd INVX1
XINVX1_738 data_memory_interface_data[18] gnd INVX1_738/Y vdd INVX1
XFILL_9_7_0 gnd vdd FILL
XXNOR2X1_13 XNOR2X1_13/A NOR2X1_29/B gnd XNOR2X1_13/Y vdd XNOR2X1
XXNOR2X1_24 NOR2X1_32/B INVX2_10/A gnd XNOR2X1_24/Y vdd XNOR2X1
XXNOR2X1_35 XNOR2X1_35/A XNOR2X1_34/Y gnd XNOR2X1_35/Y vdd XNOR2X1
XXNOR2X1_46 XNOR2X1_46/A NOR2X1_57/A gnd XNOR2X1_46/Y vdd XNOR2X1
XNAND2X1_680 BUFX2_61/A BUFX2_62/A gnd NOR2X1_393/B vdd NAND2X1
XNAND2X1_691 NOR3X1_4/A NOR2X1_60/Y gnd OAI21X1_862/C vdd NAND2X1
XINVX1_70 INVX1_70/A gnd INVX1_70/Y vdd INVX1
XINVX1_81 INVX1_81/A gnd INVX1_81/Y vdd INVX1
XINVX1_92 INVX1_92/A gnd INVX1_92/Y vdd INVX1
XBUFX2_34 BUFX2_34/A gnd data_memory_interface_frame_mask[0] vdd BUFX2
XBUFX2_12 BUFX2_12/A gnd data_memory_interface_address[11] vdd BUFX2
XBUFX2_45 INVX2_72/A gnd instruction_memory_interface_address[6] vdd BUFX2
XBUFX2_23 BUFX2_23/A gnd data_memory_interface_address[22] vdd BUFX2
XBUFX2_56 BUFX2_56/A gnd instruction_memory_interface_address[17] vdd BUFX2
XFILL_17_6_0 gnd vdd FILL
XBUFX2_67 BUFX2_67/A gnd instruction_memory_interface_address[28] vdd BUFX2
XBUFX2_78 BUFX2_78/A gnd BUFX2_78/Y vdd BUFX2
XBUFX2_89 OR2X2_52/B gnd BUFX2_89/Y vdd BUFX2
XNOR2X1_3 NOR2X1_3/A NOR2X1_3/B gnd NOR2X1_3/Y vdd NOR2X1
XAOI21X1_24 AOI21X1_24/A XNOR2X1_36/A NOR2X1_41/Y gnd XOR2X1_3/A vdd AOI21X1
XAOI21X1_13 NAND3X1_81/Y AOI21X1_13/B AOI21X1_13/C gnd AOI21X1_13/Y vdd AOI21X1
XAOI21X1_35 INVX1_295/Y AOI21X1_35/B INVX1_298/Y gnd NOR2X1_67/A vdd AOI21X1
XAOI21X1_68 INVX8_7/A AOI21X1_68/B INVX4_5/A gnd AOI21X1_68/Y vdd AOI21X1
XAOI21X1_57 AOI21X1_57/A AOI21X1_57/B AOI21X1_57/C gnd AOI21X1_57/Y vdd AOI21X1
XAOI21X1_46 INVX1_316/Y AOI21X1_46/B AOI21X1_46/C gnd AOI21X1_46/Y vdd AOI21X1
XAOI21X1_79 INVX1_378/A AOI21X1_79/B BUFX4_86/Y gnd AOI21X1_79/Y vdd AOI21X1
XOAI21X1_8 INVX1_8/Y BUFX4_23/Y OAI21X1_8/C gnd OAI21X1_8/Y vdd OAI21X1
XOAI22X1_21 OAI22X1_21/A NOR2X1_110/Y AOI21X1_62/Y AOI21X1_78/B gnd OAI22X1_21/Y vdd
+ OAI22X1
XOAI22X1_10 OAI22X1_10/A AOI22X1_80/A AOI21X1_48/Y AOI22X1_79/D gnd OAI22X1_10/Y vdd
+ OAI22X1
XOAI22X1_32 INVX2_63/Y OAI22X1_43/B INVX8_12/Y OAI22X1_7/D gnd OAI22X1_32/Y vdd OAI22X1
XOAI22X1_43 INVX2_71/Y OAI22X1_43/B INVX8_12/Y NOR2X1_86/Y gnd NOR3X1_64/C vdd OAI22X1
XFILL_41_4_0 gnd vdd FILL
XOAI22X1_54 INVX2_92/Y OAI22X1_58/B OAI22X1_58/C INVX1_737/Y gnd OAI22X1_54/Y vdd
+ OAI22X1
XOAI21X1_471 BUFX4_217/Y NOR2X1_187/Y NAND2X1_438/Y gnd NOR2X1_222/B vdd OAI21X1
XOAI21X1_460 NOR2X1_150/Y NOR2X1_151/Y AOI21X1_74/Y gnd AOI21X1_80/A vdd OAI21X1
XOAI21X1_493 INVX2_46/A MUX2X1_16/Y NAND2X1_460/A gnd AND2X2_35/A vdd OAI21X1
XOAI21X1_482 OAI21X1_412/A BUFX4_213/Y NAND2X1_455/Y gnd AOI21X1_124/B vdd OAI21X1
XINVX1_502 INVX1_502/A gnd INVX1_502/Y vdd INVX1
XINVX1_524 INVX1_524/A gnd INVX1_524/Y vdd INVX1
XINVX1_513 INVX1_513/A gnd INVX1_513/Y vdd INVX1
XINVX1_535 INVX1_535/A gnd INVX1_535/Y vdd INVX1
XINVX1_557 INVX1_557/A gnd INVX1_557/Y vdd INVX1
XINVX1_546 INVX1_619/A gnd INVX1_546/Y vdd INVX1
XINVX1_568 BUFX2_87/A gnd INVX1_568/Y vdd INVX1
XINVX1_579 INVX1_579/A gnd INVX1_579/Y vdd INVX1
XFILL_32_4_0 gnd vdd FILL
XFILL_23_4_0 gnd vdd FILL
XAOI22X1_112 OR2X2_51/Y NAND2X1_814/Y AOI22X1_112/C OR2X2_52/Y gnd BUFX4_99/A vdd
+ AOI22X1
XAOI22X1_101 INVX2_68/Y BUFX4_154/Y OR2X2_24/Y INVX2_67/Y gnd AOI22X1_101/Y vdd AOI22X1
XAOI22X1_134 AOI22X1_134/A AOI22X1_134/B INVX1_697/Y NAND2X1_974/Y gnd AOI21X1_251/A
+ vdd AOI22X1
XAOI22X1_123 OAI22X1_49/A INVX4_11/A BUFX4_261/Y BUFX2_95/A gnd AOI22X1_123/Y vdd
+ AOI22X1
XAOI22X1_145 data_memory_interface_data[9] BUFX4_107/Y AOI22X1_145/C BUFX4_9/Y gnd
+ AOI22X1_145/Y vdd AOI22X1
XAOI22X1_156 data_memory_interface_data[20] BUFX4_108/Y BUFX4_172/Y BUFX4_250/Y gnd
+ AOI22X1_156/Y vdd AOI22X1
XFILL_6_5_0 gnd vdd FILL
XBUFX4_118 BUFX4_118/A gnd BUFX4_118/Y vdd BUFX4
XAOI22X1_167 data_memory_interface_data[31] BUFX4_108/Y BUFX4_170/Y BUFX4_250/Y gnd
+ AOI22X1_167/Y vdd AOI22X1
XBUFX4_107 BUFX4_107/A gnd BUFX4_107/Y vdd BUFX4
XBUFX4_129 INVX8_7/Y gnd BUFX4_129/Y vdd BUFX4
XFILL_14_4_0 gnd vdd FILL
XOAI21X1_1019 NOR2X1_481/Y INVX4_12/A data_memory_interface_data[26] gnd OAI21X1_1019/Y
+ vdd OAI21X1
XOAI21X1_1008 OAI21X1_1007/Y data_memory_interface_data[23] OAI22X1_58/B gnd OAI21X1_1009/A
+ vdd OAI21X1
XOAI21X1_290 INVX1_314/Y INVX4_4/A NAND2X1_205/Y gnd INVX2_27/A vdd OAI21X1
XINVX1_310 INVX1_668/A gnd INVX1_310/Y vdd INVX1
XINVX1_343 INVX1_690/A gnd INVX1_343/Y vdd INVX1
XINVX1_332 OR2X2_57/A gnd INVX1_332/Y vdd INVX1
XINVX1_321 MUX2X1_44/B gnd INVX1_321/Y vdd INVX1
XINVX1_365 INVX1_365/A gnd INVX1_365/Y vdd INVX1
XINVX1_354 INVX1_354/A gnd INVX1_354/Y vdd INVX1
XINVX1_387 INVX1_387/A gnd INVX1_387/Y vdd INVX1
XINVX1_376 INVX1_376/A gnd INVX1_376/Y vdd INVX1
XINVX1_398 INVX1_398/A gnd INVX1_398/Y vdd INVX1
XAND2X2_90 OR2X2_55/A OR2X2_55/B gnd AND2X2_90/Y vdd AND2X2
XFILL_1_2 gnd vdd FILL
XFILL_43_2 gnd vdd FILL
XNAND2X1_1002 DFFPOSX1_206/Q INVX4_14/A gnd OAI21X1_953/C vdd NAND2X1
XDFFPOSX1_13 AOI22X1_13/D CLKBUF1_51/Y DFFPOSX1_13/D gnd vdd DFFPOSX1
XDFFPOSX1_35 AOI22X1_35/D CLKBUF1_50/Y DFFPOSX1_35/D gnd vdd DFFPOSX1
XNAND2X1_1024 DFFPOSX1_215/Q BUFX4_106/Y gnd NAND3X1_360/A vdd NAND2X1
XDFFPOSX1_24 AOI22X1_24/D CLKBUF1_55/Y DFFPOSX1_24/D gnd vdd DFFPOSX1
XNAND2X1_1013 data_memory_interface_data[2] OAI21X1_993/B gnd OAI21X1_989/C vdd NAND2X1
XDFFPOSX1_46 AOI22X1_8/A CLKBUF1_50/Y INVX1_98/A gnd vdd DFFPOSX1
XDFFPOSX1_68 AOI22X1_30/A CLKBUF1_50/Y INVX1_121/A gnd vdd DFFPOSX1
XDFFPOSX1_57 AOI22X1_19/A CLKBUF1_61/Y INVX1_110/A gnd vdd DFFPOSX1
XDFFPOSX1_79 INVX1_192/A CLKBUF1_31/Y OAI21X1_99/C gnd vdd DFFPOSX1
XNAND3X1_318 INVX1_635/Y BUFX4_103/Y BUFX4_164/Y gnd NAND3X1_318/Y vdd NAND3X1
XNAND3X1_329 AND2X2_1/A AND2X2_1/B INVX1_66/A gnd OAI21X1_902/B vdd NAND3X1
XNAND3X1_307 BUFX4_120/Y NAND3X1_306/Y NAND3X1_307/C gnd NAND2X1_890/B vdd NAND3X1
XFILL_30_7_1 gnd vdd FILL
XDFFPOSX1_428 BUFX2_87/A CLKBUF1_39/Y NOR3X1_35/Y gnd vdd DFFPOSX1
XDFFPOSX1_406 INVX1_666/A CLKBUF1_46/Y OAI21X1_63/Y gnd vdd DFFPOSX1
XDFFPOSX1_417 OR2X2_8/B CLKBUF1_59/Y NOR3X1_24/Y gnd vdd DFFPOSX1
XDFFPOSX1_439 INVX8_14/A CLKBUF1_44/Y NOR3X1_46/Y gnd vdd DFFPOSX1
XINVX1_140 BUFX2_94/A gnd NOR3X1_3/B vdd INVX1
XINVX1_151 NOR2X1_18/A gnd NOR3X1_12/B vdd INVX1
XNAND2X1_509 BUFX4_80/Y INVX1_371/A gnd OR2X2_40/A vdd NAND2X1
XINVX1_184 instruction_memory_interface_data[28] gnd INVX1_184/Y vdd INVX1
XINVX1_162 instruction_memory_interface_data[6] gnd INVX1_162/Y vdd INVX1
XINVX1_195 INVX1_195/A gnd INVX1_195/Y vdd INVX1
XINVX1_173 instruction_memory_interface_data[17] gnd INVX1_173/Y vdd INVX1
XFILL_37_3_0 gnd vdd FILL
XAOI21X1_100 INVX4_8/Y NOR2X1_253/B BUFX4_274/Y gnd AOI22X1_90/B vdd AOI21X1
XAOI21X1_111 AOI22X1_89/B OAI22X1_22/D OAI22X1_22/B gnd AOI21X1_111/Y vdd AOI21X1
XAOI21X1_122 AOI21X1_122/A OAI22X1_8/B OAI22X1_8/C gnd OAI21X1_602/B vdd AOI21X1
XAOI21X1_133 AOI22X1_99/B NOR2X1_293/A OAI22X1_38/B gnd OAI21X1_593/C vdd AOI21X1
XFILL_20_2_0 gnd vdd FILL
XFILL_21_7_1 gnd vdd FILL
XAOI21X1_155 OAI21X1_641/Y AND2X2_52/B AOI21X1_155/C gnd INVX1_405/A vdd AOI21X1
XAOI21X1_144 NOR2X1_304/Y AOI21X1_144/B OAI21X1_602/Y gnd AOI21X1_144/Y vdd AOI21X1
XAOI21X1_166 OAI21X1_659/Y NOR2X1_326/Y NAND3X1_152/Y gnd OAI21X1_667/C vdd AOI21X1
XAOI21X1_188 MUX2X1_49/Y INVX2_55/A INVX8_7/A gnd OAI21X1_719/C vdd AOI21X1
XAOI21X1_199 NOR2X1_72/Y INVX1_422/A NOR2X1_75/Y gnd AOI21X1_199/Y vdd AOI21X1
XAOI21X1_177 NOR2X1_81/Y AOI21X1_200/B BUFX4_276/Y gnd OAI21X1_695/C vdd AOI21X1
XFILL_28_3_0 gnd vdd FILL
XFILL_3_3_0 gnd vdd FILL
XNAND3X1_104 INVX4_5/A INVX8_10/A OAI22X1_43/B gnd NOR3X1_56/C vdd NAND3X1
XNAND3X1_115 OAI21X1_468/Y AOI22X1_84/Y AOI21X1_83/Y gnd INVX1_71/A vdd NAND3X1
XNAND3X1_148 BUFX4_91/Y OAI21X1_639/Y OAI21X1_640/Y gnd NAND3X1_148/Y vdd NAND3X1
XNAND3X1_137 OAI21X1_572/Y OR2X2_34/Y NOR2X1_290/Y gnd INVX1_80/A vdd NAND3X1
XNAND3X1_126 INVX2_48/Y INVX1_390/A INVX2_56/Y gnd NOR2X1_262/A vdd NAND3X1
XFILL_11_2_0 gnd vdd FILL
XFILL_12_7_1 gnd vdd FILL
XNAND3X1_159 NAND3X1_159/A OAI21X1_698/Y NOR3X1_62/Y gnd INVX1_90/A vdd NAND3X1
XFILL_19_3_0 gnd vdd FILL
XDFFPOSX1_203 INVX1_731/A CLKBUF1_16/Y INVX1_449/A gnd vdd DFFPOSX1
XDFFPOSX1_225 DFFPOSX1_81/D CLKBUF1_2/Y INVX1_69/A gnd vdd DFFPOSX1
XDFFPOSX1_236 DFFPOSX1_92/D CLKBUF1_23/Y INVX1_80/A gnd vdd DFFPOSX1
XDFFPOSX1_214 DFFPOSX1_214/Q CLKBUF1_16/Y INVX1_460/A gnd vdd DFFPOSX1
XBUFX4_9 BUFX4_9/A gnd BUFX4_9/Y vdd BUFX4
XDFFPOSX1_258 INVX1_239/A CLKBUF1_54/Y NAND3X1_14/A gnd vdd DFFPOSX1
XDFFPOSX1_269 MUX2X1_3/A CLKBUF1_14/Y NAND3X1_36/A gnd vdd DFFPOSX1
XDFFPOSX1_247 OAI21X1_147/C CLKBUF1_21/Y INVX1_91/A gnd vdd DFFPOSX1
XNAND2X1_306 INVX2_38/A MUX2X1_3/Y gnd AOI22X1_99/B vdd NAND2X1
XNAND2X1_317 NOR2X1_76/A INVX4_2/Y gnd OAI21X1_334/C vdd NAND2X1
XNAND2X1_339 INVX8_8/A NOR2X1_94/B gnd OAI21X1_648/C vdd NAND2X1
XNAND2X1_328 BUFX4_43/Y MUX2X1_37/B gnd NAND2X1_328/Y vdd NAND2X1
XNOR3X1_35 NOR3X1_35/A NOR3X1_35/B BUFX4_48/Y gnd NOR3X1_35/Y vdd NOR3X1
XNOR3X1_13 INVX4_1/A NOR3X1_13/B BUFX4_45/Y gnd NOR3X1_13/Y vdd NOR3X1
XNOR3X1_24 NOR3X1_35/A INVX1_165/Y NOR3X1_8/C gnd NOR3X1_24/Y vdd NOR3X1
XNOR3X1_57 NOR3X1_57/A NOR3X1_57/B NOR3X1_57/C gnd NOR3X1_57/Y vdd NOR3X1
XNOR3X1_68 NOR3X1_68/A INVX1_490/Y NOR3X1_68/C gnd NOR3X1_68/Y vdd NOR3X1
XNOR3X1_46 NOR3X1_4/A INVX1_187/Y NOR3X1_4/C gnd NOR3X1_46/Y vdd NOR3X1
XNOR3X1_79 NOR3X1_79/A INVX8_16/Y NOR3X1_80/C gnd NOR3X1_79/Y vdd NOR3X1
XNOR2X1_361 OAI22X1_41/Y NOR2X1_361/B gnd NOR2X1_361/Y vdd NOR2X1
XNOR2X1_350 BUFX4_88/Y NOR2X1_355/B gnd NOR2X1_350/Y vdd NOR2X1
XNOR2X1_383 BUFX2_47/A NOR2X1_382/Y gnd NOR2X1_383/Y vdd NOR2X1
XNOR2X1_394 NOR3X1_66/A NOR3X1_66/C gnd NOR2X1_395/B vdd NOR2X1
XNOR2X1_372 INVX8_5/A NOR2X1_372/B gnd NOR2X1_372/Y vdd NOR2X1
XOAI21X1_823 INVX1_470/A INVX2_72/Y INVX1_472/Y gnd OAI21X1_824/C vdd OAI21X1
XINVX4_9 INVX4_9/A gnd INVX4_9/Y vdd INVX4
XOAI21X1_801 BUFX4_180/Y INVX1_454/Y OAI21X1_801/C gnd OAI21X1_801/Y vdd OAI21X1
XOAI21X1_812 BUFX4_179/Y INVX1_465/Y NAND2X1_635/Y gnd OAI21X1_812/Y vdd OAI21X1
XOAI21X1_845 OAI21X1_844/Y AOI21X1_217/Y OAI21X1_845/C gnd OAI21X1_845/Y vdd OAI21X1
XOAI21X1_834 INVX1_476/Y OR2X2_47/A OAI21X1_834/C gnd OAI21X1_834/Y vdd OAI21X1
XOAI21X1_856 AOI21X1_219/Y OAI21X1_855/Y OAI21X1_856/C gnd OAI21X1_856/Y vdd OAI21X1
XOAI21X1_867 NOR3X1_68/Y BUFX2_70/A INVX8_13/Y gnd OAI21X1_867/Y vdd OAI21X1
XOAI21X1_878 OAI21X1_877/A INVX1_645/Y OAI21X1_878/C gnd OAI21X1_878/Y vdd OAI21X1
XOAI21X1_889 INVX1_660/Y OAI21X1_887/B INVX4_11/Y gnd OAI21X1_889/Y vdd OAI21X1
XNAND2X1_840 OAI21X1_72/Y BUFX4_62/Y gnd NAND2X1_840/Y vdd NAND2X1
XNAND2X1_851 NAND2X1_849/Y NAND2X1_851/B gnd NAND2X1_43/B vdd NAND2X1
XNAND2X1_873 OAI21X1_83/Y BUFX4_62/Y gnd NAND2X1_873/Y vdd NAND2X1
XNAND2X1_862 INVX1_604/Y BUFX4_97/Y gnd NAND3X1_289/C vdd NAND2X1
XNAND2X1_884 NAND2X1_882/Y NAND2X1_884/B gnd NAND2X1_54/B vdd NAND2X1
XNAND2X1_895 INVX1_626/Y BUFX4_95/Y gnd NAND3X1_311/C vdd NAND2X1
XFILL_43_1_0 gnd vdd FILL
XNAND3X1_90 OAI22X1_29/A OR2X2_32/B AOI22X1_70/Y gnd NOR2X1_108/B vdd NAND3X1
XNOR2X1_90 INVX1_433/A INVX1_432/A gnd INVX2_26/A vdd NOR2X1
XFILL_34_1_0 gnd vdd FILL
XFILL_35_6_1 gnd vdd FILL
XOAI21X1_108 BUFX4_186/Y INVX1_104/Y OAI21X1_107/Y gnd INVX1_514/A vdd OAI21X1
XOAI21X1_119 OR2X2_2/A BUFX4_194/Y OAI21X1_119/C gnd OAI21X1_120/C vdd OAI21X1
XBUFX2_6 BUFX2_6/A gnd data_memory_interface_address[5] vdd BUFX2
XNAND2X1_125 AND2X2_1/A AND2X2_1/B gnd NOR3X1_48/C vdd NAND2X1
XNAND2X1_103 AND2X2_2/B AND2X2_2/A gnd NAND3X1_7/C vdd NAND2X1
XNAND2X1_114 NOR2X1_18/A INVX1_226/Y gnd OR2X2_5/A vdd NAND2X1
XNAND2X1_158 INVX1_263/Y NAND2X1_158/B gnd OAI21X1_276/B vdd NAND2X1
XNAND2X1_147 NAND3X1_83/A NAND3X1_83/B gnd NOR2X1_46/B vdd NAND2X1
XNAND2X1_136 INVX1_251/A BUFX4_231/Y gnd NAND3X1_82/B vdd NAND2X1
XNAND2X1_169 OR2X2_13/B OR2X2_13/A gnd NAND2X1_170/A vdd NAND2X1
XNAND2X1_1 NAND2X1_1/A BUFX4_20/Y gnd OAI21X1_1/C vdd NAND2X1
XFILL_0_1_0 gnd vdd FILL
XFILL_1_6_1 gnd vdd FILL
XFILL_25_1_0 gnd vdd FILL
XFILL_26_6_1 gnd vdd FILL
XNOR2X1_191 INVX8_8/A MUX2X1_7/Y gnd NOR2X1_191/Y vdd NOR2X1
XNOR2X1_180 NOR2X1_180/A NOR2X1_176/B gnd OR2X2_24/A vdd NOR2X1
XINVX2_6 INVX2_6/A gnd INVX2_6/Y vdd INVX2
XOAI21X1_631 MUX2X1_2/Y BUFX4_39/Y OAI21X1_631/C gnd OAI21X1_662/A vdd OAI21X1
XOAI21X1_620 INVX1_403/A AND2X2_48/A NOR2X1_313/Y gnd OAI21X1_620/Y vdd OAI21X1
XOAI21X1_642 AOI21X1_37/B INVX1_402/A OAI22X1_39/B gnd AOI21X1_155/C vdd OAI21X1
XOAI21X1_664 NAND2X1_561/B BUFX4_51/Y BUFX4_125/Y gnd AOI21X1_164/C vdd OAI21X1
XOAI21X1_653 BUFX4_129/Y OR2X2_27/B OAI21X1_653/C gnd AND2X2_53/B vdd OAI21X1
XOAI21X1_675 BUFX4_129/Y NOR2X1_229/B OAI21X1_675/C gnd AND2X2_57/B vdd OAI21X1
XAOI21X1_6 AOI21X1_5/Y AOI21X1_6/B AOI21X1_6/C gnd AOI21X1_6/Y vdd AOI21X1
XINVX1_717 NOR2X1_3/A gnd INVX1_717/Y vdd INVX1
XOAI21X1_697 AOI21X1_178/Y INVX2_33/A AND2X2_62/Y gnd AOI21X1_180/C vdd OAI21X1
XOAI21X1_686 MUX2X1_56/B INVX8_3/A OAI21X1_686/C gnd OAI21X1_687/C vdd OAI21X1
XINVX1_706 INVX2_51/A gnd OR2X2_66/B vdd INVX1
XINVX1_739 data_memory_interface_data[9] gnd INVX1_739/Y vdd INVX1
XINVX1_728 INVX1_728/A gnd INVX1_728/Y vdd INVX1
XFILL_9_7_1 gnd vdd FILL
XFILL_8_2_0 gnd vdd FILL
XXNOR2X1_14 AOI21X1_10/Y INVX1_248/A gnd XNOR2X1_14/Y vdd XNOR2X1
XXNOR2X1_36 XNOR2X1_36/A NOR2X1_43/B gnd XNOR2X1_36/Y vdd XNOR2X1
XXNOR2X1_25 XNOR2X1_25/A XNOR2X1_24/Y gnd XNOR2X1_25/Y vdd XNOR2X1
XXNOR2X1_47 NOR2X1_61/Y INVX1_294/A gnd XNOR2X1_47/Y vdd XNOR2X1
XNAND2X1_670 INVX8_13/A XNOR2X1_39/Y gnd OAI21X1_845/C vdd NAND2X1
XNAND2X1_681 AND2X2_78/A AND2X2_78/B gnd NOR3X1_66/A vdd NAND2X1
XINVX1_60 gnd gnd INVX1_60/Y vdd INVX1
XNAND2X1_692 BUFX4_241/Y XNOR2X1_47/Y gnd OAI21X1_865/C vdd NAND2X1
XINVX1_82 INVX1_82/A gnd INVX1_82/Y vdd INVX1
XINVX1_93 INVX1_93/A gnd INVX1_93/Y vdd INVX1
XINVX1_71 INVX1_71/A gnd INVX1_71/Y vdd INVX1
XBUFX2_35 BUFX2_35/A gnd data_memory_interface_frame_mask[1] vdd BUFX2
XBUFX2_13 BUFX2_13/A gnd data_memory_interface_address[12] vdd BUFX2
XBUFX2_24 BUFX2_24/A gnd data_memory_interface_address[23] vdd BUFX2
XBUFX2_57 BUFX2_57/A gnd instruction_memory_interface_address[18] vdd BUFX2
XBUFX2_46 BUFX2_46/A gnd instruction_memory_interface_address[7] vdd BUFX2
XFILL_16_1_0 gnd vdd FILL
XFILL_17_6_1 gnd vdd FILL
XBUFX2_68 BUFX2_68/A gnd instruction_memory_interface_address[29] vdd BUFX2
XDFFPOSX1_1 AND2X2_5/B CLKBUF1_60/Y NAND3X1_1/B gnd vdd DFFPOSX1
XBUFX2_79 BUFX2_79/A gnd BUFX2_79/Y vdd BUFX2
XNOR2X1_4 OR2X2_69/B OR2X2_69/A gnd NOR2X1_4/Y vdd NOR2X1
XAOI21X1_25 AOI21X1_13/Y INVX1_244/Y INVX1_252/A gnd AOI21X1_26/A vdd AOI21X1
XAOI21X1_14 NAND3X1_78/Y AOI21X1_7/Y AOI21X1_14/C gnd NOR2X1_30/B vdd AOI21X1
XAOI21X1_58 BUFX4_44/Y MUX2X1_21/A AOI21X1_56/A gnd MUX2X1_25/A vdd AOI21X1
XAOI21X1_47 OR2X2_18/Y AOI21X1_47/B INVX8_3/A gnd OAI22X1_10/A vdd AOI21X1
XAOI21X1_36 INVX1_293/A AOI21X1_32/B INVX1_299/Y gnd AOI21X1_36/Y vdd AOI21X1
XAOI21X1_69 AOI21X1_69/A AOI21X1_56/A AOI21X1_69/C gnd AOI21X1_69/Y vdd AOI21X1
XOAI21X1_9 INVX1_9/Y BUFX4_17/Y OAI21X1_9/C gnd OAI21X1_9/Y vdd OAI21X1
XOAI22X1_22 AND2X2_37/Y OAI22X1_22/B NOR2X1_244/Y OAI22X1_22/D gnd NOR2X1_246/B vdd
+ OAI22X1
XOAI22X1_11 OAI22X1_11/A AOI22X1_86/A NOR2X1_232/A NOR2X1_147/Y gnd NOR2X1_152/A vdd
+ OAI22X1
XOAI22X1_33 BUFX4_127/Y OAI22X1_33/B AND2X2_45/Y INVX4_5/Y gnd OAI22X1_34/C vdd OAI22X1
XFILL_41_4_1 gnd vdd FILL
XOAI22X1_44 NOR2X1_372/Y OAI22X1_44/B OAI22X1_44/C MUX2X1_20/S gnd AND2X2_71/A vdd
+ OAI22X1
XOAI22X1_55 INVX1_739/Y OAI22X1_58/B OAI22X1_58/C INVX1_740/Y gnd OAI22X1_55/Y vdd
+ OAI22X1
XOAI21X1_450 NAND2X1_342/B BUFX4_217/Y NAND2X1_427/Y gnd OAI21X1_558/B vdd OAI21X1
XOAI21X1_461 INVX8_3/A OAI22X1_14/A OAI21X1_461/C gnd AOI21X1_75/B vdd OAI21X1
XOAI21X1_483 AOI21X1_124/B BUFX4_57/Y INVX1_388/A gnd OAI22X1_19/C vdd OAI21X1
XOAI21X1_472 MUX2X1_49/S OAI21X1_380/Y OAI21X1_472/C gnd OAI21X1_472/Y vdd OAI21X1
XINVX1_514 INVX1_514/A gnd INVX1_514/Y vdd INVX1
XOAI21X1_494 AND2X2_35/Y NOR2X1_233/Y BUFX4_91/Y gnd OAI21X1_494/Y vdd OAI21X1
XINVX1_503 INVX1_503/A gnd INVX1_503/Y vdd INVX1
XINVX1_525 INVX1_525/A gnd INVX1_525/Y vdd INVX1
XINVX1_536 INVX1_609/A gnd INVX1_536/Y vdd INVX1
XINVX1_558 INVX1_558/A gnd INVX1_558/Y vdd INVX1
XINVX1_547 INVX1_547/A gnd INVX1_547/Y vdd INVX1
XINVX1_569 INVX2_1/A gnd INVX1_569/Y vdd INVX1
XFILL_32_4_1 gnd vdd FILL
XFILL_39_0_0 gnd vdd FILL
XFILL_23_4_1 gnd vdd FILL
XAOI22X1_102 INVX2_69/Y BUFX4_155/Y OR2X2_24/Y INVX4_10/Y gnd AOI22X1_102/Y vdd AOI22X1
XAOI22X1_146 data_memory_interface_data[10] BUFX4_107/Y AOI22X1_146/C BUFX4_9/Y gnd
+ AOI22X1_146/Y vdd AOI22X1
XAOI22X1_135 INVX2_82/Y INVX1_459/A INVX1_700/Y INVX1_458/A gnd AOI22X1_135/Y vdd
+ AOI22X1
XAOI22X1_124 OAI22X1_49/A INVX4_11/A BUFX4_263/Y BUFX2_96/A gnd AOI22X1_124/Y vdd
+ AOI22X1
XAOI22X1_113 INVX1_574/Y INVX2_76/A INVX1_502/A INVX2_77/Y gnd AOI22X1_113/Y vdd AOI22X1
XFILL_6_5_1 gnd vdd FILL
XFILL_5_0_0 gnd vdd FILL
XAOI22X1_168 BUFX4_254/Y INVX1_728/A AOI22X1_168/C BUFX4_106/Y gnd AOI22X1_168/Y vdd
+ AOI22X1
XBUFX4_108 BUFX4_107/A gnd BUFX4_108/Y vdd BUFX4
XAOI22X1_157 data_memory_interface_data[21] BUFX4_108/Y BUFX4_172/Y BUFX4_250/Y gnd
+ AOI22X1_157/Y vdd AOI22X1
XBUFX4_119 BUFX4_122/A gnd BUFX4_119/Y vdd BUFX4
XFILL_14_4_1 gnd vdd FILL
XOAI21X1_1009 OAI21X1_1009/A NOR3X1_81/Y NAND3X1_357/Y gnd AOI21X1_265/B vdd OAI21X1
XOAI21X1_291 INVX4_4/Y AOI22X1_60/A OAI21X1_291/C gnd NOR2X1_332/B vdd OAI21X1
XOAI21X1_280 NOR2X1_67/A INVX1_297/A INVX1_300/Y gnd OAI21X1_280/Y vdd OAI21X1
XINVX1_300 INVX1_300/A gnd INVX1_300/Y vdd INVX1
XINVX1_344 INVX2_85/A gnd INVX1_344/Y vdd INVX1
XINVX1_333 MUX2X1_6/B gnd INVX1_333/Y vdd INVX1
XINVX1_322 OR2X2_56/A gnd INVX1_322/Y vdd INVX1
XINVX1_311 INVX1_311/A gnd INVX1_311/Y vdd INVX1
XINVX1_366 INVX1_366/A gnd INVX1_366/Y vdd INVX1
XINVX1_377 INVX1_377/A gnd OR2X2_31/A vdd INVX1
XINVX1_355 INVX1_355/A gnd INVX1_355/Y vdd INVX1
XINVX1_399 INVX1_399/A gnd INVX1_399/Y vdd INVX1
XINVX1_388 INVX1_388/A gnd INVX1_388/Y vdd INVX1
XAND2X2_91 AND2X2_91/A AND2X2_91/B gnd AND2X2_91/Y vdd AND2X2
XAND2X2_80 AND2X2_80/A AND2X2_80/B gnd BUFX4_62/A vdd AND2X2
XNAND2X1_1014 data_memory_interface_data[3] OAI21X1_993/B gnd OAI21X1_993/C vdd NAND2X1
XDFFPOSX1_14 AOI22X1_14/D CLKBUF1_24/Y DFFPOSX1_14/D gnd vdd DFFPOSX1
XNAND2X1_1003 BUFX2_78/A BUFX4_116/Y gnd OAI21X1_968/C vdd NAND2X1
XNAND2X1_1025 INVX1_727/A BUFX4_254/Y gnd NAND3X1_360/B vdd NAND2X1
XDFFPOSX1_25 AOI22X1_25/D CLKBUF1_40/Y DFFPOSX1_25/D gnd vdd DFFPOSX1
XDFFPOSX1_36 AOI22X1_36/D CLKBUF1_43/Y DFFPOSX1_36/D gnd vdd DFFPOSX1
XDFFPOSX1_47 AOI22X1_9/A CLKBUF1_31/Y INVX1_100/A gnd vdd DFFPOSX1
XDFFPOSX1_58 AOI22X1_20/A CLKBUF1_11/Y INVX1_111/A gnd vdd DFFPOSX1
XDFFPOSX1_69 AOI22X1_31/A CLKBUF1_24/Y INVX1_122/A gnd vdd DFFPOSX1
XNAND3X1_319 BUFX4_122/Y NAND3X1_318/Y NAND3X1_319/C gnd NAND2X1_908/B vdd NAND3X1
XNAND3X1_308 INVX1_625/Y BUFX4_99/Y BUFX4_167/Y gnd NAND3X1_308/Y vdd NAND3X1
XDFFPOSX1_429 INVX2_76/A CLKBUF1_20/Y NOR3X1_36/Y gnd vdd DFFPOSX1
XDFFPOSX1_407 INVX1_467/A CLKBUF1_38/Y OAI21X1_64/Y gnd vdd DFFPOSX1
XDFFPOSX1_418 OR2X2_8/A CLKBUF1_59/Y NOR3X1_25/Y gnd vdd DFFPOSX1
XINVX1_130 INVX1_130/A gnd INVX1_130/Y vdd INVX1
XINVX1_141 BUFX2_95/A gnd NOR3X1_4/B vdd INVX1
XINVX1_152 NOR2X1_14/A gnd NOR3X1_13/B vdd INVX1
XINVX1_185 instruction_memory_interface_data[29] gnd INVX1_185/Y vdd INVX1
XINVX1_163 instruction_memory_interface_data[7] gnd INVX1_163/Y vdd INVX1
XINVX1_174 instruction_memory_interface_data[18] gnd INVX1_174/Y vdd INVX1
XINVX1_196 INVX1_196/A gnd INVX1_196/Y vdd INVX1
XFILL_37_3_1 gnd vdd FILL
XAOI21X1_101 NOR2X1_248/Y BUFX4_153/Y OAI22X1_23/Y gnd OAI21X1_521/C vdd AOI21X1
XAOI21X1_112 AOI21X1_79/B NOR2X1_152/Y OAI21X1_548/Y gnd OAI21X1_551/A vdd AOI21X1
XAOI21X1_123 OAI22X1_7/C BUFX4_153/Y OAI22X1_32/Y gnd OAI21X1_578/C vdd AOI21X1
XAOI21X1_134 NAND3X1_93/C AOI21X1_134/B OAI21X1_593/Y gnd OAI21X1_594/C vdd AOI21X1
XAOI21X1_145 AOI22X1_70/Y OAI21X1_606/Y AOI21X1_145/C gnd OAI21X1_608/C vdd AOI21X1
XAOI21X1_156 AND2X2_52/Y AOI21X1_185/B INVX1_405/Y gnd INVX1_406/A vdd AOI21X1
XAOI21X1_167 INVX1_410/A INVX1_408/Y INVX2_69/Y gnd INVX1_417/A vdd AOI21X1
XFILL_20_2_1 gnd vdd FILL
XAOI21X1_178 OAI21X1_696/Y INVX1_415/Y INVX1_407/A gnd AOI21X1_178/Y vdd AOI21X1
XAOI21X1_189 INVX2_62/Y AND2X2_40/Y AOI21X1_189/C gnd AOI21X1_189/Y vdd AOI21X1
XFILL_28_3_1 gnd vdd FILL
XFILL_3_3_1 gnd vdd FILL
XNAND3X1_105 BUFX4_228/Y BUFX4_213/Y INVX2_52/A gnd NOR2X1_239/B vdd NAND3X1
XNAND3X1_138 BUFX4_92/Y NAND3X1_138/B NAND3X1_138/C gnd NAND3X1_138/Y vdd NAND3X1
XNAND3X1_116 OAI21X1_480/Y NAND3X1_116/B NOR2X1_231/Y gnd INVX1_72/A vdd NAND3X1
XNAND3X1_127 OAI21X1_535/Y NAND3X1_127/B NAND3X1_127/C gnd NOR2X1_263/B vdd NAND3X1
XNAND3X1_149 NAND3X1_147/Y NAND3X1_148/Y NAND3X1_149/C gnd INVX1_85/A vdd NAND3X1
XFILL_11_2_1 gnd vdd FILL
XFILL_19_3_1 gnd vdd FILL
XDFFPOSX1_204 INVX1_732/A CLKBUF1_28/Y INVX1_450/A gnd vdd DFFPOSX1
XDFFPOSX1_237 OAI21X1_127/C CLKBUF1_21/Y INVX1_81/A gnd vdd DFFPOSX1
XDFFPOSX1_226 OAI21X1_105/C CLKBUF1_15/Y INVX1_70/A gnd vdd DFFPOSX1
XDFFPOSX1_215 DFFPOSX1_215/Q CLKBUF1_8/Y INVX2_81/A gnd vdd DFFPOSX1
XDFFPOSX1_259 INVX1_242/A CLKBUF1_33/Y NAND3X1_16/A gnd vdd DFFPOSX1
XDFFPOSX1_248 OAI21X1_149/C CLKBUF1_23/Y INVX1_92/A gnd vdd DFFPOSX1
XNAND2X1_307 INVX2_39/A MUX2X1_4/Y gnd AOI22X1_99/C vdd NAND2X1
XNAND2X1_318 INVX1_307/A INVX4_3/Y gnd NAND2X1_318/Y vdd NAND2X1
XNAND2X1_329 INVX8_5/A NAND2X1_400/B gnd NAND2X1_329/Y vdd NAND2X1
XNOR3X1_14 INVX4_1/A INVX1_154/Y BUFX4_45/Y gnd NOR3X1_14/Y vdd NOR3X1
XNOR3X1_25 NOR3X1_35/A INVX1_166/Y NOR3X1_8/C gnd NOR3X1_25/Y vdd NOR3X1
XNOR3X1_58 NOR3X1_58/A NOR3X1_58/B NOR3X1_58/C gnd NOR3X1_58/Y vdd NOR3X1
XNOR3X1_47 INVX1_236/Y NOR2X1_6/B NOR3X1_47/C gnd NOR3X1_47/Y vdd NOR3X1
XNOR3X1_36 NOR3X1_3/A INVX1_177/Y BUFX4_45/Y gnd NOR3X1_36/Y vdd NOR3X1
XNOR3X1_69 INVX2_79/A INVX1_643/A INVX1_642/Y gnd BUFX4_262/A vdd NOR3X1
XNOR2X1_340 BUFX4_53/Y INVX2_66/Y gnd NOR2X1_340/Y vdd NOR2X1
XNOR2X1_351 NOR2X1_76/Y NOR2X1_75/Y gnd INVX1_422/A vdd NOR2X1
XNOR2X1_384 OR2X2_46/Y NOR3X1_65/C gnd INVX1_476/A vdd NOR2X1
XNOR2X1_373 BUFX4_127/Y NOR2X1_373/B gnd NOR2X1_373/Y vdd NOR2X1
XNOR2X1_395 BUFX2_63/A NOR2X1_395/B gnd NOR2X1_395/Y vdd NOR2X1
XNOR2X1_362 INVX2_22/Y NOR2X1_362/B gnd NOR2X1_362/Y vdd NOR2X1
XOAI21X1_824 INVX1_471/A NOR2X1_382/B OAI21X1_824/C gnd OAI21X1_825/A vdd OAI21X1
XOAI21X1_802 BUFX4_181/Y INVX1_455/Y NAND2X1_625/Y gnd OAI21X1_802/Y vdd OAI21X1
XOAI21X1_813 BUFX4_179/Y INVX1_466/Y NAND2X1_636/Y gnd OAI21X1_813/Y vdd OAI21X1
XOAI21X1_846 OAI21X1_846/A INVX1_481/Y INVX1_482/Y gnd OAI21X1_846/Y vdd OAI21X1
XOAI21X1_835 OAI21X1_834/Y OR2X2_45/B OAI21X1_835/C gnd OAI21X1_835/Y vdd OAI21X1
XOAI21X1_857 OAI21X1_857/A NOR2X1_395/Y NAND2X1_684/Y gnd OAI21X1_857/Y vdd OAI21X1
XOAI21X1_868 OAI21X1_867/Y NOR2X1_398/Y OAI21X1_868/C gnd OAI21X1_868/Y vdd OAI21X1
XOAI21X1_879 OAI21X1_877/A INVX1_646/Y OAI21X1_879/C gnd OAI21X1_879/Y vdd OAI21X1
XNAND2X1_830 NAND2X1_828/Y NAND3X1_267/Y gnd NAND2X1_36/B vdd NAND2X1
XNAND2X1_852 OAI21X1_76/Y BUFX4_59/Y gnd NAND2X1_852/Y vdd NAND2X1
XNAND2X1_863 NAND2X1_861/Y NAND2X1_863/B gnd NAND2X1_47/B vdd NAND2X1
XNAND2X1_841 INVX1_590/Y BUFX4_96/Y gnd NAND3X1_275/C vdd NAND2X1
XNAND2X1_896 NAND2X1_896/A NAND2X1_896/B gnd NAND2X1_58/B vdd NAND2X1
XNAND2X1_885 OAI21X1_87/Y BUFX4_63/Y gnd NAND2X1_885/Y vdd NAND2X1
XNAND2X1_874 INVX1_612/Y BUFX4_98/Y gnd NAND2X1_874/Y vdd NAND2X1
XFILL_43_1_1 gnd vdd FILL
XNAND3X1_91 INVX2_47/A INVX1_378/A NAND3X1_91/C gnd NAND3X1_91/Y vdd NAND3X1
XNAND3X1_80 INVX1_243/Y NAND3X1_80/B NAND3X1_80/C gnd NAND3X1_80/Y vdd NAND3X1
XNOR2X1_80 NOR2X1_80/A INVX2_50/A gnd NOR2X1_80/Y vdd NOR2X1
XNOR2X1_91 INVX1_315/A INVX2_27/A gnd NOR2X1_93/A vdd NOR2X1
XFILL_34_1_1 gnd vdd FILL
XOAI21X1_109 BUFX4_269/Y BUFX4_192/Y OAI21X1_109/C gnd OAI21X1_109/Y vdd OAI21X1
XBUFX2_7 BUFX2_7/A gnd data_memory_interface_address[6] vdd BUFX2
XNAND2X1_126 NOR3X1_47/Y NOR3X1_48/Y gnd AOI21X1_8/B vdd NAND2X1
XNAND2X1_115 NOR2X1_14/A NOR2X1_18/A gnd OR2X2_7/B vdd NAND2X1
XNAND2X1_104 NOR2X1_10/B AND2X2_5/Y gnd NOR2X1_8/B vdd NAND2X1
XNAND2X1_148 NAND3X1_83/B NAND2X1_148/B gnd NAND2X1_148/Y vdd NAND2X1
XNAND2X1_159 NOR2X1_50/A OAI21X1_259/Y gnd AOI21X1_27/B vdd NAND2X1
XNAND2X1_137 NAND3X1_82/Y OAI21X1_239/Y gnd AOI21X1_13/C vdd NAND2X1
XNAND2X1_2 BUFX4_23/Y NAND2X1_2/B gnd OAI21X1_2/C vdd NAND2X1
XFILL_25_1_1 gnd vdd FILL
XFILL_0_1_1 gnd vdd FILL
XNOR2X1_170 INVX2_38/A INVX2_39/A gnd NOR2X1_170/Y vdd NOR2X1
XNOR2X1_192 BUFX4_42/Y MUX2X1_5/Y gnd NOR2X1_192/Y vdd NOR2X1
XNOR2X1_181 OR2X2_24/B OR2X2_24/A gnd OAI22X1_43/B vdd NOR2X1
XINVX2_7 INVX2_7/A gnd INVX2_7/Y vdd INVX2
XOAI21X1_621 OAI21X1_621/A BUFX4_216/Y OAI21X1_621/C gnd AND2X2_67/A vdd OAI21X1
XOAI21X1_632 OAI21X1_662/A INVX8_5/A NAND2X1_548/Y gnd INVX1_404/A vdd OAI21X1
XOAI21X1_610 INVX2_67/Y INVX1_401/A BUFX4_91/Y gnd NOR2X1_309/B vdd OAI21X1
XOAI21X1_665 OAI21X1_665/A AND2X2_55/Y NOR3X1_56/Y gnd OAI21X1_665/Y vdd OAI21X1
XOAI21X1_643 AND2X2_51/Y INVX1_406/Y OAI21X1_643/C gnd NAND3X1_151/A vdd OAI21X1
XOAI21X1_654 INVX2_32/A MUX2X1_44/A BUFX4_187/Y gnd NAND3X1_150/C vdd OAI21X1
XAOI21X1_7 AOI21X1_7/A AOI21X1_7/B NOR2X1_28/Y gnd AOI21X1_7/Y vdd AOI21X1
XOAI21X1_687 BUFX4_125/Y INVX1_385/Y OAI21X1_687/C gnd AND2X2_60/B vdd OAI21X1
XOAI21X1_676 INVX2_29/A INVX2_30/A BUFX4_187/Y gnd NAND3X1_153/C vdd OAI21X1
XINVX1_707 INVX1_435/A gnd INVX1_707/Y vdd INVX1
XOAI21X1_698 NOR2X1_81/Y OAI21X1_698/B AOI21X1_181/Y gnd OAI21X1_698/Y vdd OAI21X1
XINVX1_718 BUFX2_77/A gnd INVX1_718/Y vdd INVX1
XINVX1_729 INVX1_729/A gnd INVX1_729/Y vdd INVX1
XXNOR2X1_15 XNOR2X1_15/A AOI21X1_13/C gnd XNOR2X1_15/Y vdd XNOR2X1
XFILL_8_2_1 gnd vdd FILL
XXNOR2X1_26 AOI22X1_47/Y INVX2_8/Y gnd NOR2X1_33/A vdd XNOR2X1
XXNOR2X1_37 XNOR2X1_37/A INVX1_234/A gnd XNOR2X1_37/Y vdd XNOR2X1
XXNOR2X1_48 XNOR2X1_48/A NAND2X1_98/A gnd INVX1_300/A vdd XNOR2X1
XNAND2X1_671 BUFX2_57/A BUFX2_58/A gnd NOR2X1_390/B vdd NAND2X1
XNAND2X1_660 INVX1_477/Y NOR2X1_387/B gnd OAI21X1_834/C vdd NAND2X1
XNAND2X1_682 BUFX2_63/A NOR2X1_395/B gnd XOR2X1_9/A vdd NAND2X1
XINVX1_50 gnd gnd INVX1_50/Y vdd INVX1
XNAND2X1_693 BUFX4_241/Y NOR2X1_67/Y gnd OAI21X1_866/C vdd NAND2X1
XINVX1_83 INVX1_83/A gnd INVX1_83/Y vdd INVX1
XINVX1_72 INVX1_72/A gnd INVX1_72/Y vdd INVX1
XINVX1_61 gnd gnd INVX1_61/Y vdd INVX1
XINVX1_94 INVX1_94/A gnd INVX1_94/Y vdd INVX1
XBUFX2_36 BUFX2_36/A gnd data_memory_interface_frame_mask[2] vdd BUFX2
XBUFX2_14 BUFX2_14/A gnd data_memory_interface_address[13] vdd BUFX2
XBUFX2_25 BUFX2_25/A gnd data_memory_interface_address[24] vdd BUFX2
XBUFX2_47 BUFX2_47/A gnd instruction_memory_interface_address[8] vdd BUFX2
XBUFX2_58 BUFX2_58/A gnd instruction_memory_interface_address[19] vdd BUFX2
XBUFX2_69 BUFX2_69/A gnd instruction_memory_interface_address[30] vdd BUFX2
XDFFPOSX1_2 AND2X2_5/A CLKBUF1_60/Y INVX1_715/A gnd vdd DFFPOSX1
XFILL_16_1_1 gnd vdd FILL
XNOR2X1_5 INVX1_66/A NOR2X1_1/A gnd NOR2X1_5/Y vdd NOR2X1
XAOI21X1_15 MUX2X1_9/B BUFX4_150/Y NOR3X1_53/Y gnd AOI21X1_15/Y vdd AOI21X1
XAOI21X1_26 AOI21X1_26/A AOI21X1_26/B AOI21X1_26/C gnd AOI21X1_26/Y vdd AOI21X1
XAOI21X1_37 NOR2X1_95/Y AOI21X1_37/B NOR2X1_94/Y gnd AOI21X1_37/Y vdd AOI21X1
XAOI21X1_48 AOI21X1_48/A AOI21X1_48/B INVX8_4/A gnd AOI21X1_48/Y vdd AOI21X1
XAOI21X1_59 BUFX4_124/Y AOI21X1_59/B INVX1_357/Y gnd AOI21X1_59/Y vdd AOI21X1
XOAI22X1_12 NOR2X1_149/Y NOR2X1_148/Y NOR2X1_150/Y NOR2X1_151/Y gnd OAI22X1_12/Y vdd
+ OAI22X1
XOAI22X1_23 INVX2_58/Y OAI22X1_43/B INVX8_12/Y NOR2X1_249/Y gnd OAI22X1_23/Y vdd OAI22X1
XOAI22X1_34 OAI22X1_30/A OAI22X1_34/B OAI22X1_34/C OAI22X1_34/D gnd OAI22X1_34/Y vdd
+ OAI22X1
XOAI22X1_56 INVX1_742/Y OAI22X1_58/B OAI22X1_58/C INVX1_743/Y gnd OAI22X1_56/Y vdd
+ OAI22X1
XOAI22X1_45 INVX2_75/Y INVX1_495/A INVX1_501/Y INVX2_73/A gnd OAI22X1_45/Y vdd OAI22X1
XOAI21X1_440 INVX1_361/Y INVX8_5/A OAI21X1_440/C gnd MUX2X1_32/A vdd OAI21X1
XOAI21X1_484 NAND2X1_430/B BUFX4_223/Y NAND2X1_457/Y gnd OAI21X1_485/B vdd OAI21X1
XOAI21X1_451 INVX1_375/Y INVX8_4/A OAI21X1_451/C gnd OAI22X1_14/A vdd OAI21X1
XOAI21X1_473 BUFX4_53/Y NOR2X1_223/Y OAI21X1_473/C gnd INVX1_379/A vdd OAI21X1
XOAI21X1_462 OR2X2_23/A INVX1_376/Y OR2X2_31/A gnd NAND2X1_435/B vdd OAI21X1
XOAI21X1_495 OAI21X1_470/A MUX2X1_40/S NAND2X1_464/Y gnd OAI21X1_543/B vdd OAI21X1
XINVX1_515 INVX1_515/A gnd INVX1_515/Y vdd INVX1
XINVX1_526 INVX1_599/A gnd INVX1_526/Y vdd INVX1
XINVX1_504 INVX1_504/A gnd INVX1_504/Y vdd INVX1
XINVX1_548 INVX1_621/A gnd INVX1_548/Y vdd INVX1
XINVX1_537 INVX1_537/A gnd INVX1_537/Y vdd INVX1
XINVX1_559 INVX1_632/A gnd INVX1_559/Y vdd INVX1
XNAND2X1_490 BUFX4_229/Y OAI21X1_531/Y gnd NAND2X1_490/Y vdd NAND2X1
XFILL_39_0_1 gnd vdd FILL
XAOI22X1_103 INVX1_414/Y BUFX4_155/Y OR2X2_24/Y OR2X2_38/B gnd AOI22X1_103/Y vdd AOI22X1
XAOI22X1_136 OR2X2_67/A NOR2X1_460/Y NAND2X1_993/Y INVX1_713/Y gnd AOI22X1_136/Y vdd
+ AOI22X1
XAOI22X1_125 OAI22X1_49/A INVX4_11/A BUFX4_263/Y BUFX2_97/A gnd AOI22X1_125/Y vdd
+ AOI22X1
XAOI22X1_114 OAI22X1_49/A OAI21X1_887/B NOR2X1_412/Y OAI22X1_6/Y gnd OAI21X1_877/A
+ vdd AOI22X1
XAOI22X1_169 BUFX4_252/Y INVX1_731/A AOI22X1_169/C BUFX4_106/Y gnd AOI22X1_169/Y vdd
+ AOI22X1
XAOI22X1_158 data_memory_interface_data[22] BUFX4_109/Y BUFX4_169/Y BUFX4_253/Y gnd
+ AOI22X1_158/Y vdd AOI22X1
XBUFX4_109 BUFX4_107/A gnd BUFX4_109/Y vdd BUFX4
XAOI22X1_147 data_memory_interface_data[11] BUFX4_107/Y AOI22X1_147/C BUFX4_10/Y gnd
+ AOI22X1_147/Y vdd AOI22X1
XFILL_5_0_1 gnd vdd FILL
XFILL_42_7_0 gnd vdd FILL
XOAI21X1_292 INVX1_318/Y INVX4_4/A NAND2X1_208/Y gnd MUX2X1_46/B vdd OAI21X1
XINVX1_301 OR2X2_1/B gnd NOR2X1_70/B vdd INVX1
XOAI21X1_281 INVX1_302/Y INVX4_4/A NAND2X1_196/Y gnd INVX2_17/A vdd OAI21X1
XOAI21X1_270 XOR2X1_6/A XOR2X1_6/B INVX2_15/Y gnd XNOR2X1_45/A vdd OAI21X1
XINVX1_334 MUX2X1_7/B gnd INVX1_334/Y vdd INVX1
XINVX1_323 MUX2X1_1/B gnd INVX1_323/Y vdd INVX1
XINVX1_312 NOR2X1_89/A gnd NOR2X1_88/A vdd INVX1
XINVX1_378 INVX1_378/A gnd INVX1_378/Y vdd INVX1
XINVX1_345 OR2X2_61/A gnd INVX1_345/Y vdd INVX1
XINVX1_367 INVX1_367/A gnd INVX1_367/Y vdd INVX1
XINVX1_356 INVX1_356/A gnd INVX1_356/Y vdd INVX1
XINVX1_389 INVX1_389/A gnd INVX1_389/Y vdd INVX1
XAND2X2_70 AND2X2_70/A AND2X2_70/B gnd AND2X2_70/Y vdd AND2X2
XAND2X2_81 AND2X2_81/A AND2X2_81/B gnd AND2X2_81/Y vdd AND2X2
XAND2X2_92 AND2X2_92/A AND2X2_92/B gnd AND2X2_92/Y vdd AND2X2
XFILL_33_7_0 gnd vdd FILL
XDFFPOSX1_15 AOI22X1_15/D CLKBUF1_18/Y DFFPOSX1_15/D gnd vdd DFFPOSX1
XNAND2X1_1026 DFFPOSX1_217/Q BUFX4_106/Y gnd NAND3X1_361/A vdd NAND2X1
XNAND2X1_1004 BUFX2_79/A BUFX4_116/Y gnd OAI21X1_969/C vdd NAND2X1
XDFFPOSX1_26 AOI22X1_26/D CLKBUF1_42/Y DFFPOSX1_26/D gnd vdd DFFPOSX1
XNAND2X1_1015 data_memory_interface_data[4] OAI21X1_993/B gnd OAI21X1_997/C vdd NAND2X1
XDFFPOSX1_48 AOI22X1_10/A CLKBUF1_24/Y INVX1_101/A gnd vdd DFFPOSX1
XDFFPOSX1_59 AOI22X1_21/A CLKBUF1_11/Y INVX1_112/A gnd vdd DFFPOSX1
XDFFPOSX1_37 AOI22X1_37/D CLKBUF1_51/Y DFFPOSX1_37/D gnd vdd DFFPOSX1
XFILL_24_7_0 gnd vdd FILL
XNAND3X1_309 BUFX4_123/Y NAND3X1_308/Y NAND3X1_309/C gnd NAND2X1_893/B vdd NAND3X1
XFILL_15_7_0 gnd vdd FILL
XDFFPOSX1_408 INVX1_149/A CLKBUF1_20/Y NAND3X1_70/Y gnd vdd DFFPOSX1
XDFFPOSX1_419 NOR2X1_23/A CLKBUF1_59/Y NOR3X1_26/Y gnd vdd DFFPOSX1
XINVX1_142 BUFX2_96/A gnd NOR3X1_5/B vdd INVX1
XINVX1_131 BUFX2_92/A gnd NOR3X1_1/B vdd INVX1
XINVX1_120 INVX1_120/A gnd INVX1_120/Y vdd INVX1
XINVX1_175 instruction_memory_interface_data[19] gnd INVX1_175/Y vdd INVX1
XINVX1_186 instruction_memory_interface_data[30] gnd INVX1_186/Y vdd INVX1
XINVX1_153 INVX1_228/A gnd INVX1_153/Y vdd INVX1
XINVX1_164 instruction_memory_interface_data[8] gnd INVX1_164/Y vdd INVX1
XINVX1_197 INVX1_197/A gnd INVX1_197/Y vdd INVX1
XAOI21X1_102 AOI22X1_72/Y AOI21X1_92/B OAI21X1_526/Y gnd AOI22X1_92/C vdd AOI21X1
XAOI21X1_113 AOI22X1_71/Y AOI21X1_113/B AOI21X1_113/C gnd AOI21X1_113/Y vdd AOI21X1
XAOI21X1_124 BUFX4_57/Y AOI21X1_124/B AOI21X1_124/C gnd OAI22X1_34/D vdd AOI21X1
XAOI21X1_135 INVX1_399/A AOI21X1_180/B BUFX4_87/Y gnd OAI21X1_595/C vdd AOI21X1
XAOI21X1_146 NOR2X1_108/Y AOI21X1_92/B AOI21X1_146/C gnd NOR2X1_308/B vdd AOI21X1
XAOI21X1_157 AND2X2_51/Y INVX1_406/Y INVX8_11/A gnd OAI21X1_643/C vdd AOI21X1
XAOI21X1_168 INVX2_70/Y AOI21X1_168/B INVX8_11/A gnd OAI21X1_670/C vdd AOI21X1
XAOI21X1_179 NOR2X1_333/Y AOI21X1_38/B NOR2X1_332/Y gnd AND2X2_62/B vdd AOI21X1
XNAND3X1_139 NAND3X1_138/Y OAI21X1_582/Y NAND3X1_139/C gnd INVX1_81/A vdd NAND3X1
XNAND3X1_117 INVX8_11/Y OAI21X1_491/Y NAND3X1_117/C gnd NAND3X1_117/Y vdd NAND3X1
XNAND3X1_106 BUFX4_124/Y NOR2X1_182/Y NOR3X1_56/Y gnd NAND3X1_106/Y vdd NAND3X1
XNAND3X1_128 OAI21X1_528/Y AOI22X1_95/Y NOR2X1_263/Y gnd INVX1_76/A vdd NAND3X1
XFILL_30_5_0 gnd vdd FILL
XDFFPOSX1_227 DFFPOSX1_83/D CLKBUF1_31/Y INVX1_71/A gnd vdd DFFPOSX1
XDFFPOSX1_216 AOI22X1_168/C CLKBUF1_28/Y OR2X2_55/B gnd vdd DFFPOSX1
XDFFPOSX1_205 INVX1_733/A CLKBUF1_8/Y INVX1_451/A gnd vdd DFFPOSX1
XDFFPOSX1_238 OAI21X1_129/C CLKBUF1_15/Y INVX1_82/A gnd vdd DFFPOSX1
XDFFPOSX1_249 OAI21X1_151/C CLKBUF1_57/Y INVX1_93/A gnd vdd DFFPOSX1
XNAND2X1_308 AOI21X1_42/Y NAND2X1_308/B gnd AOI21X1_43/C vdd NAND2X1
XNAND2X1_319 NOR2X1_80/A INVX2_50/Y gnd NAND2X1_319/Y vdd NAND2X1
XNOR3X1_26 INVX4_1/A NOR3X1_26/B NOR3X1_8/C gnd NOR3X1_26/Y vdd NOR3X1
XNOR3X1_15 INVX4_1/A INVX1_155/Y NOR3X1_8/C gnd NOR3X1_15/Y vdd NOR3X1
XFILL_38_6_0 gnd vdd FILL
XNOR3X1_59 NOR3X1_59/A AND2X2_53/Y NOR3X1_59/C gnd NOR3X1_59/Y vdd NOR3X1
XNOR3X1_48 NOR3X1_48/A NOR2X1_1/A NOR3X1_48/C gnd NOR3X1_48/Y vdd NOR3X1
XNOR3X1_37 NOR3X1_35/A INVX1_178/Y BUFX4_48/Y gnd NOR3X1_37/Y vdd NOR3X1
XBUFX4_270 NAND3X1_1/Y gnd BUFX4_270/Y vdd BUFX4
XNOR2X1_330 INVX8_3/A MUX2X1_45/Y gnd NOR2X1_330/Y vdd NOR2X1
XNOR2X1_341 AOI21X1_38/B INVX2_70/A gnd NOR2X1_341/Y vdd NOR2X1
XNOR2X1_352 NOR2X1_352/A NOR2X1_352/B gnd NOR2X1_352/Y vdd NOR2X1
XNOR2X1_385 BUFX2_51/A INVX1_476/A gnd NOR2X1_385/Y vdd NOR2X1
XNOR2X1_374 INVX1_315/A INVX2_27/Y gnd INVX1_434/A vdd NOR2X1
XNOR2X1_363 BUFX4_88/Y NOR2X1_362/Y gnd NOR2X1_363/Y vdd NOR2X1
XNOR2X1_396 NOR3X1_66/B INVX1_491/A gnd INVX1_487/A vdd NOR2X1
XFILL_21_5_0 gnd vdd FILL
XOAI21X1_803 BUFX4_181/Y INVX1_456/Y NAND2X1_626/Y gnd OAI21X1_803/Y vdd OAI21X1
XOAI21X1_814 BUFX4_179/Y INVX1_467/Y NAND2X1_637/Y gnd OAI21X1_814/Y vdd OAI21X1
XOAI21X1_825 OAI21X1_825/A OR2X2_45/B OAI21X1_825/C gnd OAI21X1_168/C vdd OAI21X1
XOAI21X1_836 XNOR2X1_51/Y BUFX4_245/Y OAI21X1_836/C gnd OAI21X1_836/Y vdd OAI21X1
XOAI21X1_847 NAND2X1_673/Y INVX8_13/A OAI21X1_847/C gnd OAI21X1_847/Y vdd OAI21X1
XOAI21X1_858 XOR2X1_9/Y BUFX4_241/Y OAI21X1_858/C gnd OAI21X1_858/Y vdd OAI21X1
XOAI21X1_869 INVX2_74/Y INVX1_502/A INVX1_504/A gnd NOR2X1_401/A vdd OAI21X1
XNAND2X1_831 OAI21X1_69/Y BUFX4_60/Y gnd NAND2X1_831/Y vdd NAND2X1
XNAND2X1_820 NAND2X1_820/A AOI22X1_113/Y gnd NOR2X1_408/B vdd NAND2X1
XNAND2X1_864 OAI21X1_80/Y BUFX4_60/Y gnd NAND2X1_864/Y vdd NAND2X1
XNAND2X1_842 NAND2X1_840/Y NAND2X1_842/B gnd NAND2X1_40/B vdd NAND2X1
XNAND2X1_853 INVX1_598/Y BUFX4_96/Y gnd NAND3X1_283/C vdd NAND2X1
XNAND2X1_897 OAI21X1_91/Y BUFX4_63/Y gnd NAND2X1_897/Y vdd NAND2X1
XNAND2X1_875 NAND2X1_873/Y NAND2X1_875/B gnd NAND2X1_51/B vdd NAND2X1
XNAND2X1_886 INVX1_620/Y BUFX4_97/Y gnd NAND3X1_305/C vdd NAND2X1
XFILL_4_6_0 gnd vdd FILL
XFILL_29_6_0 gnd vdd FILL
XFILL_12_5_0 gnd vdd FILL
XNAND3X1_81 INVX1_245/A NAND3X1_81/B NAND3X1_81/C gnd NAND3X1_81/Y vdd NAND3X1
XNAND3X1_92 NAND3X1_92/A INVX1_352/A INVX1_348/Y gnd AND2X2_21/A vdd NAND3X1
XNAND3X1_70 INVX4_1/Y INVX1_156/Y NAND3X1_7/C gnd NAND3X1_70/Y vdd NAND3X1
XNOR2X1_70 NOR2X1_6/B NOR2X1_70/B gnd NOR2X1_70/Y vdd NOR2X1
XNOR2X1_81 NOR2X1_80/Y INVX2_19/Y gnd NOR2X1_81/Y vdd NOR2X1
XNOR2X1_92 INVX1_315/Y INVX2_27/Y gnd NOR2X1_93/B vdd NOR2X1
XBUFX2_8 BUFX2_8/A gnd data_memory_interface_address[7] vdd BUFX2
XNAND2X1_105 NOR2X1_13/A INVX1_190/Y gnd NOR2X1_9/B vdd NAND2X1
XNAND2X1_116 INVX1_685/A BUFX4_148/Y gnd AOI21X1_5/B vdd NAND2X1
XNAND2X1_149 XNOR2X1_33/Y XNOR2X1_34/Y gnd NOR2X1_39/A vdd NAND2X1
XNAND2X1_138 AOI21X1_13/Y NOR2X1_29/Y gnd AOI21X1_14/C vdd NAND2X1
XNAND2X1_127 NAND3X1_79/Y OAI21X1_232/Y gnd NOR2X1_29/A vdd NAND2X1
XNAND2X1_3 BUFX4_24/Y NAND2X1_3/B gnd OAI21X1_3/C vdd NAND2X1
XNOR2X1_160 INVX8_8/A NOR2X1_160/B gnd NOR2X1_160/Y vdd NOR2X1
XNOR2X1_171 NOR2X1_171/A OR2X2_21/Y gnd NOR2X1_171/Y vdd NOR2X1
XNOR2X1_182 INVX8_3/A NOR2X1_239/B gnd NOR2X1_182/Y vdd NOR2X1
XNOR2X1_193 INVX1_369/Y OAI22X1_43/B gnd NOR2X1_193/Y vdd NOR2X1
XINVX2_8 INVX2_8/A gnd INVX2_8/Y vdd INVX2
XOAI21X1_633 INVX8_4/A INVX1_404/Y NAND2X1_547/Y gnd MUX2X1_50/A vdd OAI21X1
XOAI21X1_600 OAI21X1_694/A NOR2X1_103/Y INVX1_329/A gnd OAI21X1_605/B vdd OAI21X1
XOAI21X1_611 INVX2_67/A OAI21X1_609/Y NOR2X1_309/Y gnd OAI21X1_611/Y vdd OAI21X1
XOAI21X1_622 NOR2X1_315/Y NOR2X1_314/Y BUFX4_125/Y gnd OAI21X1_623/C vdd OAI21X1
XOAI21X1_644 INVX2_34/Y NOR2X1_94/B NOR2X1_319/Y gnd OAI21X1_644/Y vdd OAI21X1
XOAI21X1_666 INVX1_410/Y INVX8_12/Y AOI22X1_102/Y gnd AOI21X1_165/C vdd OAI21X1
XOAI21X1_655 OR2X2_24/A OR2X2_24/B AND2X2_51/Y gnd OAI21X1_655/Y vdd OAI21X1
XAOI21X1_8 AOI21X1_8/A AOI21X1_8/B INVX1_235/Y gnd AOI21X1_8/Y vdd AOI21X1
XOAI21X1_688 NOR2X1_334/Y AND2X2_61/Y BUFX4_125/Y gnd AOI21X1_173/A vdd OAI21X1
XOAI21X1_677 OR2X2_24/A OR2X2_24/B INVX2_70/Y gnd OAI21X1_677/Y vdd OAI21X1
XOAI21X1_699 NOR2X1_332/B BUFX4_38/Y OAI21X1_699/C gnd OAI21X1_725/B vdd OAI21X1
XINVX1_708 INVX1_708/A gnd INVX1_708/Y vdd INVX1
XINVX1_719 INVX1_719/A gnd INVX1_719/Y vdd INVX1
XXNOR2X1_27 NOR2X1_32/B INVX2_10/Y gnd NOR2X1_34/B vdd XNOR2X1
XXNOR2X1_16 XNOR2X1_16/A INVX1_249/A gnd XNOR2X1_16/Y vdd XNOR2X1
XXNOR2X1_38 AOI22X1_45/Y INVX1_243/A gnd XNOR2X1_38/Y vdd XNOR2X1
XXNOR2X1_49 XNOR2X1_49/A INVX2_58/Y gnd AOI22X1_92/B vdd XNOR2X1
XNAND2X1_661 BUFX2_51/A BUFX2_52/A gnd OR2X2_47/A vdd NAND2X1
XNAND2X1_650 INVX8_13/Y XOR2X1_8/A gnd OAI21X1_826/A vdd NAND2X1
XNAND2X1_672 AND2X2_78/A NOR3X1_65/Y gnd OR2X2_48/A vdd NAND2X1
XINVX1_51 gnd gnd INVX1_51/Y vdd INVX1
XINVX1_40 gnd gnd INVX1_40/Y vdd INVX1
XNAND2X1_694 BUFX2_69/A INVX1_490/A gnd INVX1_492/A vdd NAND2X1
XNAND2X1_683 INVX8_13/Y XOR2X1_9/A gnd OAI21X1_857/A vdd NAND2X1
XINVX1_73 INVX1_73/A gnd INVX1_73/Y vdd INVX1
XINVX1_62 gnd gnd INVX1_62/Y vdd INVX1
XINVX1_84 INVX1_84/A gnd INVX1_84/Y vdd INVX1
XBUFX2_15 BUFX2_15/A gnd data_memory_interface_address[14] vdd BUFX2
XBUFX2_26 BUFX2_26/A gnd data_memory_interface_address[25] vdd BUFX2
XINVX1_95 INVX1_95/A gnd INVX1_95/Y vdd INVX1
XBUFX2_37 BUFX2_37/A gnd data_memory_interface_frame_mask[3] vdd BUFX2
XBUFX2_48 XOR2X1_8/B gnd instruction_memory_interface_address[9] vdd BUFX2
XBUFX2_59 BUFX2_59/A gnd instruction_memory_interface_address[20] vdd BUFX2
XDFFPOSX1_3 NOR2X1_10/B CLKBUF1_62/Y OR2X2_69/A gnd vdd DFFPOSX1
XNOR2X1_6 NOR2X1_6/A NOR2X1_6/B gnd NOR2X1_6/Y vdd NOR2X1
XFILL_35_4_0 gnd vdd FILL
XAOI21X1_16 AOI21X1_8/A AOI21X1_8/B INVX1_255/Y gnd AOI21X1_16/Y vdd AOI21X1
XAOI21X1_27 AOI21X1_27/A AOI21X1_27/B INVX1_265/Y gnd XOR2X1_4/A vdd AOI21X1
XAOI21X1_38 AOI21X1_38/A AOI21X1_38/B NOR2X1_99/Y gnd AOI21X1_38/Y vdd AOI21X1
XAOI21X1_49 INVX1_376/A AOI21X1_49/B INVX1_377/A gnd NOR2X1_185/B vdd AOI21X1
XFILL_1_4_0 gnd vdd FILL
XFILL_26_4_0 gnd vdd FILL
XOAI22X1_24 NOR2X1_124/Y OAI22X1_24/B OAI22X1_24/C OAI22X1_24/D gnd NOR2X1_253/A vdd
+ OAI22X1
XOAI22X1_13 INVX1_369/A AOI21X1_56/A AOI21X1_60/Y NOR2X1_193/Y gnd OAI22X1_13/Y vdd
+ OAI22X1
XOAI22X1_35 BUFX4_128/Y INVX1_397/Y AND2X2_45/Y INVX4_5/Y gnd NOR2X1_295/B vdd OAI22X1
XOAI22X1_57 INVX1_745/Y OAI22X1_58/B OAI22X1_58/C INVX1_746/Y gnd OAI22X1_57/Y vdd
+ OAI22X1
XOAI22X1_46 INVX2_73/Y INVX1_501/A INVX1_502/Y INVX2_74/A gnd OAI22X1_46/Y vdd OAI22X1
XOAI21X1_430 INVX8_5/A OAI21X1_393/Y NAND2X1_415/Y gnd MUX2X1_22/B vdd OAI21X1
XOAI21X1_441 NOR2X1_235/B INVX8_5/A INVX8_4/A gnd OAI21X1_441/Y vdd OAI21X1
XOAI21X1_452 BUFX4_39/Y MUX2X1_11/Y OAI21X1_452/C gnd NAND2X1_430/B vdd OAI21X1
XOAI21X1_463 OAI21X1_463/A OAI22X1_20/A AOI22X1_82/Y gnd AOI21X1_75/C vdd OAI21X1
XOAI21X1_474 OAI21X1_474/A INVX8_4/A OAI21X1_474/C gnd AOI21X1_118/B vdd OAI21X1
XINVX1_505 INVX1_578/A gnd INVX1_505/Y vdd INVX1
XOAI21X1_485 INVX8_4/A OAI21X1_485/B OAI21X1_485/C gnd AOI22X1_98/A vdd OAI21X1
XOAI21X1_496 AND2X2_32/A BUFX4_216/Y NAND2X1_465/Y gnd MUX2X1_38/B vdd OAI21X1
XINVX1_516 INVX1_589/A gnd INVX1_516/Y vdd INVX1
XINVX1_527 INVX1_527/A gnd INVX1_527/Y vdd INVX1
XINVX1_549 INVX1_549/A gnd INVX1_549/Y vdd INVX1
XINVX1_538 INVX1_611/A gnd INVX1_538/Y vdd INVX1
XFILL_9_5_0 gnd vdd FILL
XNAND2X1_480 INVX2_44/A MUX2X1_9/Y gnd NAND2X1_481/A vdd NAND2X1
XNAND2X1_491 BUFX4_57/Y NOR2X1_315/A gnd OAI21X1_534/C vdd NAND2X1
XFILL_17_4_0 gnd vdd FILL
XOAI21X1_90 INVX1_91/Y BUFX4_162/Y NAND2X1_92/Y gnd OAI21X1_90/Y vdd OAI21X1
XAOI22X1_137 data_memory_interface_data[0] BUFX4_105/Y OAI21X1_981/Y BUFX4_8/Y gnd
+ OAI21X1_982/C vdd AOI22X1
XAOI22X1_104 NOR2X1_78/Y BUFX4_152/Y OR2X2_24/Y AND2X2_64/B gnd NAND3X1_162/C vdd
+ AOI22X1
XAOI22X1_126 AOI22X1_126/A OR2X2_53/Y NAND2X1_933/Y NAND2X1_932/Y gnd AOI22X1_126/Y
+ vdd AOI22X1
XAOI22X1_115 OAI22X1_49/A INVX4_11/A BUFX4_262/Y BUFX2_87/A gnd OAI21X1_891/C vdd
+ AOI22X1
XAOI22X1_148 data_memory_interface_data[12] BUFX4_107/Y AOI22X1_148/C BUFX4_9/Y gnd
+ AOI22X1_148/Y vdd AOI22X1
XAOI22X1_159 data_memory_interface_data[23] INVX4_14/A BUFX4_169/Y BUFX4_253/Y gnd
+ AOI22X1_159/Y vdd AOI22X1
XFILL_42_7_1 gnd vdd FILL
XFILL_41_2_0 gnd vdd FILL
XOAI21X1_260 INVX1_266/Y INVX1_267/Y NAND3X1_84/C gnd NAND2X1_163/B vdd OAI21X1
XOAI21X1_271 NOR2X1_54/B INVX2_15/Y INVX1_280/Y gnd INVX1_281/A vdd OAI21X1
XOAI21X1_282 INVX1_304/Y INVX4_4/A NAND2X1_197/Y gnd INVX4_2/A vdd OAI21X1
XINVX1_324 MUX2X1_2/B gnd INVX1_324/Y vdd INVX1
XINVX1_335 OR2X2_59/A gnd INVX1_335/Y vdd INVX1
XOAI21X1_293 INVX1_319/Y INVX4_4/A NAND2X1_210/Y gnd INVX2_30/A vdd OAI21X1
XINVX1_313 INVX1_664/A gnd INVX1_313/Y vdd INVX1
XINVX1_302 OR2X2_55/A gnd INVX1_302/Y vdd INVX1
XINVX1_368 INVX1_368/A gnd INVX1_368/Y vdd INVX1
XINVX1_357 AND2X2_31/B gnd INVX1_357/Y vdd INVX1
XINVX1_346 INVX1_66/A gnd INVX1_346/Y vdd INVX1
XAND2X2_60 NOR3X1_56/Y AND2X2_60/B gnd AND2X2_60/Y vdd AND2X2
XINVX1_379 INVX1_379/A gnd INVX1_379/Y vdd INVX1
XAND2X2_71 AND2X2_71/A INVX2_55/A gnd AND2X2_71/Y vdd AND2X2
XAND2X2_82 AND2X2_82/A AND2X2_82/B gnd AND2X2_82/Y vdd AND2X2
XAND2X2_93 AND2X2_93/A AND2X2_93/B gnd AND2X2_93/Y vdd AND2X2
XFILL_32_2_0 gnd vdd FILL
XFILL_33_7_1 gnd vdd FILL
XNAND2X1_1016 data_memory_interface_data[5] OAI21X1_993/B gnd NAND2X1_1016/Y vdd NAND2X1
XDFFPOSX1_16 AOI22X1_16/D CLKBUF1_18/Y DFFPOSX1_16/D gnd vdd DFFPOSX1
XNAND2X1_1027 INVX1_729/A BUFX4_254/Y gnd NAND3X1_361/B vdd NAND2X1
XNAND2X1_1005 BUFX2_80/A BUFX4_117/Y gnd NAND3X1_361/C vdd NAND2X1
XDFFPOSX1_27 AOI22X1_27/D CLKBUF1_42/Y DFFPOSX1_27/D gnd vdd DFFPOSX1
XDFFPOSX1_38 AOI22X1_38/D CLKBUF1_12/Y DFFPOSX1_38/D gnd vdd DFFPOSX1
XDFFPOSX1_49 AOI22X1_11/A CLKBUF1_55/Y INVX1_102/A gnd vdd DFFPOSX1
XFILL_23_2_0 gnd vdd FILL
XFILL_24_7_1 gnd vdd FILL
XFILL_6_3_0 gnd vdd FILL
XFILL_15_7_1 gnd vdd FILL
XFILL_14_2_0 gnd vdd FILL
XDFFPOSX1_409 INVX1_150/A CLKBUF1_20/Y NAND3X1_71/Y gnd vdd DFFPOSX1
XINVX1_110 INVX1_110/A gnd INVX1_110/Y vdd INVX1
XINVX1_143 BUFX2_97/A gnd NOR3X1_6/B vdd INVX1
XINVX1_121 INVX1_121/A gnd INVX1_121/Y vdd INVX1
XINVX1_132 BUFX2_87/A gnd INVX1_132/Y vdd INVX1
XINVX1_176 instruction_memory_interface_data[20] gnd NOR3X1_35/B vdd INVX1
XINVX1_154 INVX1_225/A gnd INVX1_154/Y vdd INVX1
XINVX1_165 instruction_memory_interface_data[9] gnd INVX1_165/Y vdd INVX1
XINVX1_187 instruction_memory_interface_data[31] gnd INVX1_187/Y vdd INVX1
XINVX1_198 INVX1_198/A gnd INVX1_198/Y vdd INVX1
XFILL_34_1 gnd vdd FILL
XAOI21X1_103 INVX2_59/Y NOR2X1_254/Y BUFX4_274/Y gnd AOI21X1_103/Y vdd AOI21X1
XAOI21X1_114 AOI22X1_96/Y NOR2X1_254/A OAI21X1_553/Y gnd AOI21X1_114/Y vdd AOI21X1
XAOI21X1_147 OAI21X1_391/Y INVX4_7/A OAI21X1_617/Y gnd AOI21X1_147/Y vdd AOI21X1
XAOI21X1_136 INVX8_3/A NOR2X1_238/B INVX8_7/A gnd AOI21X1_136/Y vdd AOI21X1
XAOI21X1_158 NOR2X1_104/Y AOI21X1_180/B OAI21X1_646/Y gnd NOR2X1_325/B vdd AOI21X1
XAOI21X1_125 INVX2_64/Y NOR2X1_294/Y BUFX4_274/Y gnd AOI21X1_125/Y vdd AOI21X1
XAOI21X1_169 BUFX4_38/Y INVX2_30/A NOR2X1_201/B gnd OAI21X1_700/A vdd AOI21X1
XNAND3X1_129 INVX1_393/Y OAI22X1_25/C INVX1_392/A gnd NAND3X1_129/Y vdd NAND3X1
XNAND3X1_118 BUFX4_79/Y INVX2_54/A INVX1_382/Y gnd NAND3X1_119/A vdd NAND3X1
XNAND3X1_107 AND2X2_27/Y NAND3X1_106/Y AOI21X1_56/Y gnd AOI21X1_57/C vdd NAND3X1
XFILL_30_5_1 gnd vdd FILL
XDFFPOSX1_217 DFFPOSX1_217/Q CLKBUF1_28/Y OR2X2_54/B gnd vdd DFFPOSX1
XDFFPOSX1_228 OAI21X1_109/C CLKBUF1_23/Y INVX1_72/A gnd vdd DFFPOSX1
XDFFPOSX1_206 DFFPOSX1_206/Q CLKBUF1_16/Y INVX1_452/A gnd vdd DFFPOSX1
XDFFPOSX1_239 DFFPOSX1_95/D CLKBUF1_3/Y INVX1_83/A gnd vdd DFFPOSX1
XNAND2X1_309 NOR2X1_89/A INVX2_25/Y gnd NAND3X1_92/A vdd NAND2X1
XNOR3X1_16 NOR3X1_16/A NOR3X1_16/B XOR2X1_1/Y gnd AOI22X1_7/A vdd NOR3X1
XNOR3X1_49 INVX1_239/Y AOI21X1_4/C NOR3X1_49/C gnd NOR3X1_49/Y vdd NOR3X1
XNOR3X1_27 NOR3X1_9/A INVX1_168/Y NOR3X1_9/C gnd NOR3X1_27/Y vdd NOR3X1
XNOR3X1_38 NOR3X1_35/A NOR3X1_38/B BUFX4_48/Y gnd NOR3X1_38/Y vdd NOR3X1
XFILL_37_1_0 gnd vdd FILL
XFILL_38_6_1 gnd vdd FILL
XBUFX4_260 BUFX4_262/A gnd BUFX4_260/Y vdd BUFX4
XBUFX4_271 NAND3X1_1/Y gnd OR2X2_2/A vdd BUFX4
XNOR2X1_320 NOR2X1_319/Y AND2X2_48/Y gnd NOR2X1_320/Y vdd NOR2X1
XNOR2X1_342 NOR2X1_342/A NOR2X1_342/B gnd NOR2X1_342/Y vdd NOR2X1
XNOR2X1_331 INVX8_10/A AND2X2_58/Y gnd NOR2X1_331/Y vdd NOR2X1
XNOR2X1_386 OR2X2_46/A OR2X2_46/B gnd NOR2X1_386/Y vdd NOR2X1
XNOR2X1_353 BUFX4_55/Y MUX2X1_50/A gnd MUX2X1_52/B vdd NOR2X1
XNOR2X1_364 NOR2X1_86/Y NOR2X1_87/Y gnd INVX2_71/A vdd NOR2X1
XNOR2X1_375 NOR2X1_375/A INVX1_436/Y gnd BUFX4_264/A vdd NOR2X1
XNOR2X1_397 INVX1_488/Y INVX1_489/Y gnd INVX1_490/A vdd NOR2X1
XFILL_20_0_0 gnd vdd FILL
XOAI21X1_815 INVX1_468/Y NOR3X1_4/A OAI21X1_815/C gnd OAI21X1_161/C vdd OAI21X1
XOAI21X1_804 BUFX4_180/Y INVX1_457/Y NAND2X1_627/Y gnd OAI21X1_804/Y vdd OAI21X1
XFILL_21_5_1 gnd vdd FILL
XOAI21X1_837 INVX1_476/Y OR2X2_47/Y INVX8_13/Y gnd OAI21X1_837/Y vdd OAI21X1
XOAI21X1_826 OAI21X1_826/A NOR2X1_383/Y OAI21X1_826/C gnd OAI21X1_169/C vdd OAI21X1
XOAI21X1_848 OR2X2_48/A INVX1_483/Y INVX8_13/Y gnd OAI21X1_848/Y vdd OAI21X1
XOAI21X1_859 XNOR2X1_52/Y BUFX4_241/Y OAI21X1_859/C gnd OAI21X1_859/Y vdd OAI21X1
XNAND2X1_821 NAND2X1_812/Y NAND2X1_821/B gnd NAND2X1_33/A vdd NAND2X1
XNAND2X1_810 INVX2_76/A INVX1_570/Y gnd NAND3X1_257/A vdd NAND2X1
XNAND2X1_843 OAI21X1_73/Y BUFX4_61/Y gnd NAND2X1_843/Y vdd NAND2X1
XNAND2X1_854 NAND2X1_852/Y NAND2X1_854/B gnd NAND2X1_44/B vdd NAND2X1
XNAND2X1_832 INVX1_584/Y BUFX4_95/Y gnd NAND3X1_269/C vdd NAND2X1
XNAND2X1_876 OAI21X1_84/Y BUFX4_63/Y gnd NAND2X1_876/Y vdd NAND2X1
XNAND2X1_887 NAND2X1_885/Y NAND2X1_887/B gnd NAND2X1_55/B vdd NAND2X1
XNAND2X1_865 INVX1_606/Y BUFX4_95/Y gnd NAND3X1_291/C vdd NAND2X1
XNAND2X1_898 INVX1_628/Y BUFX4_97/Y gnd NAND3X1_313/C vdd NAND2X1
XFILL_4_6_1 gnd vdd FILL
XFILL_28_1_0 gnd vdd FILL
XFILL_29_6_1 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XFILL_12_5_1 gnd vdd FILL
XFILL_11_0_0 gnd vdd FILL
XNAND3X1_93 AOI22X1_71/Y AOI22X1_72/Y NAND3X1_93/C gnd NAND3X1_93/Y vdd NAND3X1
XNAND3X1_82 INVX1_249/Y NAND3X1_82/B NAND3X1_82/C gnd NAND3X1_82/Y vdd NAND3X1
XNAND3X1_60 NAND3X1_60/A AND2X2_2/B AND2X2_2/A gnd NAND3X1_61/B vdd NAND3X1
XNAND3X1_71 INVX4_1/Y INVX1_157/Y NAND3X1_7/C gnd NAND3X1_71/Y vdd NAND3X1
XFILL_19_1_0 gnd vdd FILL
XNOR2X1_71 NOR2X1_71/A NOR2X1_71/B gnd OR2X2_44/B vdd NOR2X1
XNOR2X1_60 NOR2X1_61/B NOR2X1_59/Y gnd NOR2X1_60/Y vdd NOR2X1
XNOR2X1_82 NOR2X1_81/Y AND2X2_64/B gnd NOR2X1_82/Y vdd NOR2X1
XNOR2X1_93 NOR2X1_93/A NOR2X1_93/B gnd INVX2_28/A vdd NOR2X1
XBUFX2_9 BUFX2_9/A gnd data_memory_interface_address[8] vdd BUFX2
XNAND2X1_106 NOR2X1_11/A INVX1_189/A gnd NOR2X1_13/B vdd NAND2X1
XNAND2X1_117 NOR2X1_24/Y AND2X2_9/Y gnd AOI21X1_4/A vdd NAND2X1
XNAND2X1_139 INVX1_248/A XNOR2X1_16/Y gnd NOR2X1_42/A vdd NAND2X1
XNAND2X1_128 INVX2_85/A BUFX4_147/Y gnd NAND3X1_80/C vdd NAND2X1
XNAND2X1_4 BUFX4_18/Y NAND2X1_4/B gnd OAI21X1_4/C vdd NAND2X1
XNOR2X1_150 BUFX4_126/Y AND2X2_34/A gnd NOR2X1_150/Y vdd NOR2X1
XNOR2X1_161 BUFX4_44/Y INVX1_321/Y gnd NOR2X1_201/B vdd NOR2X1
XNOR2X1_194 INVX8_6/A OR2X2_29/B gnd NOR2X1_194/Y vdd NOR2X1
XNOR2X1_183 INVX2_56/A INVX1_348/A gnd BUFX4_188/A vdd NOR2X1
XNOR2X1_172 NOR2X1_135/A INVX1_355/Y gnd AND2X2_23/A vdd NOR2X1
XINVX2_9 INVX2_9/A gnd INVX2_9/Y vdd INVX2
XOAI21X1_601 NOR2X1_302/B OAI21X1_601/B OAI21X1_601/C gnd AOI21X1_144/B vdd OAI21X1
XOAI21X1_612 OAI21X1_612/A MUX2X1_40/S NAND2X1_537/Y gnd NAND2X1_556/B vdd OAI21X1
XOAI21X1_623 BUFX4_126/Y INVX1_372/A OAI21X1_623/C gnd AND2X2_49/A vdd OAI21X1
XOAI21X1_634 INVX8_3/A MUX2X1_50/A OAI21X1_634/C gnd NAND2X1_549/B vdd OAI21X1
XOAI21X1_645 INVX2_34/A MUX2X1_1/Y OAI21X1_644/Y gnd INVX1_407/A vdd OAI21X1
XOAI21X1_656 OAI21X1_457/A OR2X2_40/A AOI21X1_162/Y gnd NOR3X1_59/C vdd OAI21X1
XOAI21X1_667 AND2X2_54/Y OAI21X1_667/B OAI21X1_667/C gnd INVX1_87/A vdd OAI21X1
XOAI21X1_678 OR2X2_40/A OAI22X1_19/B OAI21X1_678/C gnd NOR3X1_60/C vdd OAI21X1
XAOI21X1_9 AOI21X1_8/A AOI21X1_8/B AOI21X1_9/C gnd AOI21X1_9/Y vdd AOI21X1
XOAI21X1_689 INVX1_317/A MUX2X1_46/B BUFX4_187/Y gnd OAI21X1_689/Y vdd OAI21X1
XINVX1_709 INVX1_443/A gnd INVX1_709/Y vdd INVX1
XXNOR2X1_17 AOI22X1_47/Y INVX2_8/A gnd XNOR2X1_17/Y vdd XNOR2X1
XXNOR2X1_28 XNOR2X1_28/A INVX2_11/A gnd NAND3X1_83/C vdd XNOR2X1
XXNOR2X1_39 AOI21X1_27/B OR2X2_11/B gnd XNOR2X1_39/Y vdd XNOR2X1
XNAND2X1_651 BUFX4_245/Y XNOR2X1_18/Y gnd OAI21X1_826/C vdd NAND2X1
XNAND2X1_662 OR2X2_45/B XNOR2X1_30/Y gnd OAI21X1_835/C vdd NAND2X1
XNAND2X1_673 OR2X2_48/A OAI21X1_846/Y gnd NAND2X1_673/Y vdd NAND2X1
XNAND2X1_640 NOR3X1_9/A XNOR2X1_5/Y gnd OAI21X1_816/C vdd NAND2X1
XINVX1_30 gnd gnd INVX1_30/Y vdd INVX1
XINVX1_41 gnd gnd INVX1_41/Y vdd INVX1
XNAND2X1_695 INVX8_13/Y NOR2X1_398/B gnd NAND2X1_695/Y vdd NAND2X1
XNAND2X1_684 BUFX4_241/Y XOR2X1_6/Y gnd NAND2X1_684/Y vdd NAND2X1
XINVX1_74 INVX1_74/A gnd INVX1_74/Y vdd INVX1
XINVX1_63 gnd gnd INVX1_63/Y vdd INVX1
XINVX1_85 INVX1_85/A gnd INVX1_85/Y vdd INVX1
XINVX1_52 gnd gnd INVX1_52/Y vdd INVX1
XBUFX2_16 BUFX2_16/A gnd data_memory_interface_address[15] vdd BUFX2
XBUFX2_27 BUFX2_27/A gnd data_memory_interface_address[26] vdd BUFX2
XINVX1_96 INVX1_96/A gnd INVX1_96/Y vdd INVX1
XBUFX2_38 BUFX2_38/A gnd data_memory_interface_state vdd BUFX2
XBUFX2_49 BUFX2_49/A gnd instruction_memory_interface_address[10] vdd BUFX2
XDFFPOSX1_4 NOR2X1_8/A CLKBUF1_60/Y OR2X2_69/B gnd vdd DFFPOSX1
XNOR2X1_7 NOR2X1_7/A NOR2X1_7/B gnd NOR2X1_7/Y vdd NOR2X1
XFILL_35_4_1 gnd vdd FILL
XAOI21X1_17 AOI21X1_17/A AOI21X1_17/B NOR2X1_31/Y gnd XNOR2X1_25/A vdd AOI21X1
XNAND3X1_290 INVX1_607/Y BUFX4_102/Y BUFX4_168/Y gnd NAND3X1_290/Y vdd NAND3X1
XAOI21X1_39 AOI21X1_39/A INVX2_33/Y AOI21X1_39/C gnd AOI21X1_39/Y vdd AOI21X1
XAOI21X1_28 NOR2X1_45/Y INVX1_272/A AOI21X1_28/C gnd XOR2X1_5/A vdd AOI21X1
XFILL_1_4_1 gnd vdd FILL
XFILL_26_4_1 gnd vdd FILL
XOAI22X1_14 OAI22X1_14/A INVX2_55/Y OAI22X1_14/C BUFX4_57/Y gnd AND2X2_33/A vdd OAI22X1
XOAI22X1_25 AOI22X1_93/Y OAI22X1_9/D OAI22X1_25/C AOI22X1_94/Y gnd OAI22X1_25/Y vdd
+ OAI22X1
XOAI22X1_58 INVX1_748/Y OAI22X1_58/B OAI22X1_58/C INVX1_749/Y gnd OAI22X1_58/Y vdd
+ OAI22X1
XOAI22X1_36 OAI22X1_20/A OAI22X1_36/B INVX2_64/Y OAI22X1_43/B gnd OAI22X1_36/Y vdd
+ OAI22X1
XOAI22X1_47 INVX2_78/Y BUFX2_87/A INVX1_574/Y INVX2_76/A gnd OAI22X1_47/Y vdd OAI22X1
XOAI21X1_431 INVX1_367/Y BUFX4_227/Y NAND2X1_416/Y gnd MUX2X1_33/B vdd OAI21X1
XOAI21X1_420 BUFX4_58/Y AND2X2_29/Y NOR2X1_204/Y gnd OAI21X1_421/C vdd OAI21X1
XOAI21X1_453 BUFX4_228/Y MUX2X1_21/Y NAND2X1_430/Y gnd OAI21X1_506/B vdd OAI21X1
XOAI21X1_464 OAI22X1_21/A AOI22X1_81/D AOI22X1_81/A gnd AOI21X1_77/C vdd OAI21X1
XOAI21X1_475 INVX8_3/A MUX2X1_27/Y OAI21X1_475/C gnd NAND2X1_444/A vdd OAI21X1
XOAI21X1_442 MUX2X1_32/A INVX8_4/A OAI21X1_441/Y gnd OR2X2_41/A vdd OAI21X1
XINVX1_506 INVX1_579/A gnd INVX1_506/Y vdd INVX1
XOAI21X1_486 AOI21X1_77/Y OAI22X1_12/Y AOI21X1_88/Y gnd NOR2X1_228/B vdd OAI21X1
XOAI21X1_497 MUX2X1_32/Y INVX8_3/A OAI21X1_497/C gnd AOI22X1_87/B vdd OAI21X1
XINVX1_517 INVX1_517/A gnd INVX1_517/Y vdd INVX1
XINVX1_528 INVX1_601/A gnd INVX1_528/Y vdd INVX1
XINVX1_539 INVX1_539/A gnd INVX1_539/Y vdd INVX1
XFILL_9_5_1 gnd vdd FILL
XFILL_8_0_0 gnd vdd FILL
XNAND2X1_481 NAND2X1_481/A NAND2X1_297/Y gnd INVX2_58/A vdd NAND2X1
XNAND2X1_470 BUFX4_77/Y MUX2X1_30/A gnd AOI22X1_88/A vdd NAND2X1
XNAND2X1_492 NOR2X1_256/Y NOR3X1_56/Y gnd NAND3X1_127/C vdd NAND2X1
XFILL_17_4_1 gnd vdd FILL
XOAI21X1_80 INVX1_81/Y BUFX4_159/Y OAI21X1_80/C gnd OAI21X1_80/Y vdd OAI21X1
XOAI21X1_91 INVX1_92/Y BUFX4_160/Y OAI21X1_91/C gnd OAI21X1_91/Y vdd OAI21X1
XAOI22X1_105 NOR2X1_75/Y BUFX4_152/Y OR2X2_24/Y INVX1_422/A gnd OAI21X1_739/C vdd
+ AOI22X1
XAOI22X1_127 OR2X2_54/Y NAND2X1_934/Y AOI22X1_127/C OR2X2_55/Y gnd AOI22X1_127/Y vdd
+ AOI22X1
XAOI22X1_116 OAI22X1_49/A INVX4_11/A BUFX4_262/Y INVX2_76/A gnd OAI21X1_892/C vdd
+ AOI22X1
XAOI22X1_149 data_memory_interface_data[13] BUFX4_105/Y AOI22X1_149/C BUFX4_8/Y gnd
+ AOI22X1_149/Y vdd AOI22X1
XAOI22X1_138 data_memory_interface_data[1] BUFX4_105/Y AOI22X1_138/C BUFX4_8/Y gnd
+ AOI22X1_138/Y vdd AOI22X1
XFILL_41_2_1 gnd vdd FILL
XOAI21X1_250 AOI21X1_19/Y NOR3X1_54/Y INVX1_258/A gnd NAND3X1_83/A vdd OAI21X1
XOAI21X1_261 OR2X2_11/A OR2X2_10/Y NAND2X1_163/Y gnd INVX1_269/A vdd OAI21X1
XOAI21X1_283 NOR2X1_75/Y NOR2X1_76/Y INVX2_18/Y gnd INVX1_305/A vdd OAI21X1
XOAI21X1_272 XOR2X1_6/A INVX1_282/Y INVX1_281/Y gnd XNOR2X1_46/A vdd OAI21X1
XINVX1_325 INVX1_325/A gnd INVX1_325/Y vdd INVX1
XOAI21X1_294 INVX1_320/Y INVX4_4/A OAI21X1_294/C gnd MUX2X1_44/B vdd OAI21X1
XINVX1_303 NOR2X1_76/A gnd INVX1_303/Y vdd INVX1
XINVX1_314 INVX1_667/A gnd INVX1_314/Y vdd INVX1
XINVX1_336 MUX2X1_9/B gnd INVX1_336/Y vdd INVX1
XINVX1_369 INVX1_369/A gnd INVX1_369/Y vdd INVX1
XAND2X2_50 OR2X2_42/A INVX4_7/Y gnd AND2X2_50/Y vdd AND2X2
XINVX1_358 INVX1_358/A gnd INVX1_358/Y vdd INVX1
XINVX1_347 OR2X2_22/B gnd INVX1_347/Y vdd INVX1
XAND2X2_72 INVX4_9/A MUX2X1_56/B gnd AND2X2_72/Y vdd AND2X2
XAND2X2_61 INVX2_55/A MUX2X1_56/B gnd AND2X2_61/Y vdd AND2X2
XAND2X2_83 AND2X2_83/A AND2X2_83/B gnd AND2X2_83/Y vdd AND2X2
XAND2X2_94 INVX1_686/Y OR2X2_62/B gnd AND2X2_94/Y vdd AND2X2
XFILL_32_2_1 gnd vdd FILL
XNAND2X1_1017 data_memory_interface_data[6] OAI21X1_993/B gnd NAND2X1_1017/Y vdd NAND2X1
XDFFPOSX1_17 AOI22X1_17/D CLKBUF1_2/Y DFFPOSX1_17/D gnd vdd DFFPOSX1
XNAND2X1_1006 BUFX2_81/A BUFX4_115/Y gnd OAI21X1_971/C vdd NAND2X1
XDFFPOSX1_39 AOI22X1_39/D CLKBUF1_31/Y DFFPOSX1_39/D gnd vdd DFFPOSX1
XNAND2X1_1028 DFFPOSX1_218/Q BUFX4_106/Y gnd NAND3X1_362/A vdd NAND2X1
XDFFPOSX1_28 AOI22X1_28/D CLKBUF1_19/Y DFFPOSX1_28/D gnd vdd DFFPOSX1
XFILL_23_2_1 gnd vdd FILL
XFILL_6_3_1 gnd vdd FILL
XFILL_14_2_1 gnd vdd FILL
XINVX1_100 INVX1_100/A gnd INVX1_100/Y vdd INVX1
XINVX1_111 INVX1_111/A gnd INVX1_111/Y vdd INVX1
XINVX1_122 INVX1_122/A gnd INVX1_122/Y vdd INVX1
XINVX1_133 OR2X2_52/B gnd AOI22X1_2/D vdd INVX1
XINVX1_144 INVX8_14/A gnd NOR3X1_7/B vdd INVX1
XINVX1_177 instruction_memory_interface_data[21] gnd INVX1_177/Y vdd INVX1
XINVX1_155 INVX2_4/A gnd INVX1_155/Y vdd INVX1
XINVX1_166 instruction_memory_interface_data[10] gnd INVX1_166/Y vdd INVX1
XINVX1_188 INVX1_188/A gnd INVX1_188/Y vdd INVX1
XINVX1_199 INVX1_199/A gnd INVX1_199/Y vdd INVX1
XFILL_34_2 gnd vdd FILL
XAOI21X1_104 NAND2X1_481/A OAI22X1_24/D OAI22X1_24/B gnd OAI21X1_529/C vdd AOI21X1
XAOI21X1_115 INVX2_62/Y OAI22X1_28/Y OAI21X1_560/Y gnd AOI21X1_115/Y vdd AOI21X1
XAOI21X1_137 AOI21X1_137/A NAND2X1_533/Y OAI22X1_30/C gnd NOR2X1_300/A vdd AOI21X1
XAOI21X1_126 BUFX4_51/Y INVX1_384/Y AOI21X1_126/C gnd NOR2X1_295/A vdd AOI21X1
XAOI21X1_148 INVX1_401/Y INVX2_67/A NOR2X1_96/Y gnd OAI21X1_646/A vdd AOI21X1
XAOI21X1_159 AND2X2_51/Y NOR2X1_325/B INVX8_10/A gnd OAI21X1_647/C vdd AOI21X1
XNAND3X1_119 NAND3X1_119/A AOI22X1_87/Y AOI21X1_89/Y gnd AOI21X1_90/C vdd NAND3X1
XNAND3X1_108 AOI22X1_76/Y AOI22X1_77/Y OAI22X1_13/Y gnd NOR2X1_200/A vdd NAND3X1
XDFFPOSX1_218 DFFPOSX1_218/Q CLKBUF1_22/Y OR2X2_53/B gnd vdd DFFPOSX1
XDFFPOSX1_207 INVX1_719/A CLKBUF1_22/Y INVX2_83/A gnd vdd DFFPOSX1
XDFFPOSX1_229 OAI21X1_111/C CLKBUF1_2/Y INVX1_73/A gnd vdd DFFPOSX1
XNOR3X1_17 NOR3X1_17/A NOR3X1_17/B XOR2X1_2/Y gnd NOR3X1_17/Y vdd NOR3X1
XNOR3X1_28 NOR3X1_4/A INVX1_169/Y NOR3X1_4/C gnd NOR3X1_28/Y vdd NOR3X1
XNOR3X1_39 NOR3X1_3/A INVX1_180/Y BUFX4_49/Y gnd NOR3X1_39/Y vdd NOR3X1
XNOR2X1_310 NOR2X1_310/A OAI22X1_30/C gnd NOR3X1_57/A vdd NOR2X1
XBUFX4_261 BUFX4_262/A gnd BUFX4_261/Y vdd BUFX4
XBUFX4_272 NAND3X1_1/Y gnd BUFX4_272/Y vdd BUFX4
XBUFX4_250 BUFX4_253/A gnd BUFX4_250/Y vdd BUFX4
XFILL_37_1_1 gnd vdd FILL
XNOR2X1_321 AOI21X1_37/B INVX1_403/A gnd AND2X2_52/B vdd NOR2X1
XNOR2X1_332 INVX1_317/A NOR2X1_332/B gnd NOR2X1_332/Y vdd NOR2X1
XNOR2X1_343 NOR2X1_80/A INVX2_50/Y gnd INVX1_419/A vdd NOR2X1
XNOR2X1_365 NOR2X1_85/B INVX2_71/A gnd NOR2X1_365/Y vdd NOR2X1
XNOR2X1_354 INVX2_16/A INVX2_17/Y gnd NOR2X1_354/Y vdd NOR2X1
XNOR2X1_376 OR2X2_63/B BUFX4_177/Y gnd NOR2X1_378/B vdd NOR2X1
XNOR2X1_387 INVX1_477/Y NOR2X1_387/B gnd XNOR2X1_51/A vdd NOR2X1
XNOR2X1_398 INVX1_493/Y NOR2X1_398/B gnd NOR2X1_398/Y vdd NOR2X1
XOAI21X1_805 BUFX4_180/Y INVX1_458/Y NAND2X1_628/Y gnd OAI21X1_805/Y vdd OAI21X1
XOAI21X1_838 AOI21X1_216/Y OAI21X1_837/Y OAI21X1_838/C gnd OAI21X1_838/Y vdd OAI21X1
XOAI21X1_827 XOR2X1_8/Y BUFX4_245/Y OAI21X1_827/C gnd OAI21X1_827/Y vdd OAI21X1
XOAI21X1_849 OAI21X1_848/Y AOI21X1_218/Y OAI21X1_849/C gnd OAI21X1_849/Y vdd OAI21X1
XOAI21X1_816 INVX1_469/Y NOR3X1_4/A OAI21X1_816/C gnd OAI21X1_816/Y vdd OAI21X1
XFILL_20_0_1 gnd vdd FILL
XNAND2X1_822 OAI21X1_66/Y BUFX4_61/Y gnd NAND2X1_822/Y vdd NAND2X1
XNAND2X1_800 INVX1_563/Y BUFX4_205/Y gnd NAND3X1_251/C vdd NAND2X1
XNAND2X1_811 XOR2X1_2/A INVX2_77/Y gnd NAND3X1_257/B vdd NAND2X1
XNAND2X1_855 OAI21X1_77/Y BUFX4_59/Y gnd NAND2X1_855/Y vdd NAND2X1
XNAND2X1_833 NAND2X1_831/Y NAND2X1_833/B gnd NAND2X1_37/B vdd NAND2X1
XNAND2X1_844 INVX1_592/Y BUFX4_95/Y gnd NAND3X1_277/C vdd NAND2X1
XNAND2X1_888 OAI21X1_88/Y BUFX4_63/Y gnd NAND2X1_890/A vdd NAND2X1
XNAND2X1_866 NAND2X1_864/Y NAND2X1_866/B gnd NAND2X1_48/B vdd NAND2X1
XNAND2X1_877 INVX1_614/Y BUFX4_97/Y gnd NAND3X1_299/C vdd NAND2X1
XNAND2X1_899 NAND2X1_897/Y NAND2X1_899/B gnd NAND2X1_59/B vdd NAND2X1
XFILL_3_1_1 gnd vdd FILL
XFILL_28_1_1 gnd vdd FILL
XFILL_11_0_1 gnd vdd FILL
XNAND3X1_50 NAND3X1_50/A BUFX4_114/Y BUFX4_137/Y gnd NAND3X1_51/B vdd NAND3X1
XNAND3X1_83 NAND3X1_83/A NAND3X1_83/B NAND3X1_83/C gnd NOR2X1_39/B vdd NAND3X1
XNAND3X1_61 BUFX4_76/Y NAND3X1_61/B NAND3X1_61/C gnd NAND3X1_61/Y vdd NAND3X1
XNAND3X1_72 INVX4_1/Y INVX1_160/Y NAND3X1_7/C gnd NAND3X1_72/Y vdd NAND3X1
XNAND3X1_94 NAND3X1_94/A NOR2X1_153/Y NAND3X1_94/C gnd NAND3X1_94/Y vdd NAND3X1
XFILL_19_1_1 gnd vdd FILL
XNOR2X1_50 NOR2X1_50/A OR2X2_11/Y gnd NOR2X1_50/Y vdd NOR2X1
XNOR2X1_72 INVX2_16/Y INVX2_17/Y gnd NOR2X1_72/Y vdd NOR2X1
XNOR2X1_61 NOR2X1_58/Y NOR2X1_61/B gnd NOR2X1_61/Y vdd NOR2X1
XNOR2X1_94 INVX2_34/Y NOR2X1_94/B gnd NOR2X1_94/Y vdd NOR2X1
XNOR2X1_83 INVX2_20/A INVX2_21/A gnd NOR2X1_85/A vdd NOR2X1
XNAND2X1_107 AOI22X1_40/Y NAND3X1_73/Y gnd OR2X2_4/B vdd NAND2X1
XNAND2X1_129 INVX1_242/A BUFX4_232/Y gnd NAND3X1_80/B vdd NAND2X1
XNAND2X1_118 AND2X2_9/Y AND2X2_10/Y gnd AOI21X1_4/B vdd NAND2X1
XNAND2X1_5 BUFX4_21/Y NAND2X1_5/B gnd OAI21X1_5/C vdd NAND2X1
XNOR2X1_140 BUFX4_54/Y MUX2X1_11/Y gnd AOI22X1_80/A vdd NOR2X1
XNOR2X1_151 INVX8_7/A NOR2X1_151/B gnd NOR2X1_151/Y vdd NOR2X1
XNOR2X1_173 NOR2X1_203/B OR2X2_36/B gnd AND2X2_31/B vdd NOR2X1
XNOR2X1_184 BUFX4_44/Y MUX2X1_13/Y gnd AOI21X1_56/A vdd NOR2X1
XNOR2X1_162 NOR2X1_89/A INVX1_315/A gnd NOR2X1_162/Y vdd NOR2X1
XNOR2X1_195 NOR2X1_195/A INVX1_369/Y gnd NOR2X1_195/Y vdd NOR2X1
XOAI21X1_613 BUFX4_214/Y MUX2X1_36/Y NAND2X1_538/Y gnd OAI21X1_719/A vdd OAI21X1
XOAI21X1_602 NOR2X1_304/B OAI21X1_602/B AOI21X1_143/Y gnd OAI21X1_602/Y vdd OAI21X1
XOAI21X1_624 AND2X2_67/A INVX8_3/A AOI21X1_149/Y gnd AOI21X1_150/A vdd OAI21X1
XOAI21X1_635 BUFX4_125/Y INVX1_374/A OAI21X1_635/C gnd AOI21X1_154/B vdd OAI21X1
XOAI21X1_646 OAI21X1_646/A OR2X2_39/B INVX1_407/Y gnd OAI21X1_646/Y vdd OAI21X1
XOAI21X1_657 INVX1_406/A NAND3X1_89/B INVX1_408/A gnd AND2X2_54/A vdd OAI21X1
XOAI21X1_679 NOR2X1_101/Y INVX1_409/A INVX1_411/A gnd INVX1_413/A vdd OAI21X1
XOAI21X1_668 INVX1_411/Y NOR2X1_101/Y AND2X2_51/Y gnd NOR2X1_336/A vdd OAI21X1
XXNOR2X1_18 NOR2X1_35/B XNOR2X1_17/Y gnd XNOR2X1_18/Y vdd XNOR2X1
XXNOR2X1_29 NOR2X1_36/Y NAND3X1_83/C gnd XNOR2X1_29/Y vdd XNOR2X1
XNAND2X1_630 INVX1_278/A BUFX4_266/Y gnd NAND2X1_630/Y vdd NAND2X1
XNAND2X1_663 BUFX4_245/Y XNOR2X1_32/Y gnd OAI21X1_836/C vdd NAND2X1
XNAND2X1_652 BUFX4_245/Y XNOR2X1_19/Y gnd OAI21X1_827/C vdd NAND2X1
XNAND2X1_641 INVX8_13/A XNOR2X1_7/Y gnd OAI21X1_817/C vdd NAND2X1
XINVX1_20 gnd gnd INVX1_20/Y vdd INVX1
XINVX1_31 gnd gnd INVX1_31/Y vdd INVX1
XINVX1_42 gnd gnd INVX1_42/Y vdd INVX1
XNAND2X1_674 INVX8_13/A XOR2X1_4/Y gnd OAI21X1_847/C vdd NAND2X1
XNAND2X1_696 BUFX4_241/Y NAND2X1_192/Y gnd OAI21X1_868/C vdd NAND2X1
XNAND2X1_685 NOR3X1_9/A XNOR2X1_45/Y gnd OAI21X1_858/C vdd NAND2X1
XINVX1_75 INVX1_75/A gnd INVX1_75/Y vdd INVX1
XINVX1_64 gnd gnd INVX1_64/Y vdd INVX1
XINVX1_53 gnd gnd INVX1_53/Y vdd INVX1
XBUFX2_17 BUFX2_17/A gnd data_memory_interface_address[16] vdd BUFX2
XINVX1_97 INVX1_97/A gnd INVX1_97/Y vdd INVX1
XINVX1_86 INVX1_86/A gnd INVX1_86/Y vdd INVX1
XBUFX2_39 BUFX2_39/A gnd instruction_memory_interface_address[0] vdd BUFX2
XBUFX2_28 BUFX2_28/A gnd data_memory_interface_address[27] vdd BUFX2
XDFFPOSX1_5 NOR2X1_13/A CLKBUF1_60/Y NOR2X1_3/B gnd vdd DFFPOSX1
XNOR2X1_8 NOR2X1_8/A NOR2X1_8/B gnd AND2X2_6/A vdd NOR2X1
XNAND3X1_291 BUFX4_120/Y NAND3X1_290/Y NAND3X1_291/C gnd NAND2X1_866/B vdd NAND3X1
XNAND3X1_280 INVX1_597/Y BUFX4_101/Y BUFX4_166/Y gnd NAND3X1_280/Y vdd NAND3X1
XAOI21X1_18 NOR2X1_31/Y XNOR2X1_24/Y NOR2X1_32/Y gnd AOI21X1_18/Y vdd AOI21X1
XAOI21X1_29 AOI21X1_29/A AOI21X1_29/B AOI21X1_29/C gnd NOR2X1_51/B vdd AOI21X1
XOAI22X1_15 OAI22X1_20/A OAI22X1_15/B INVX2_47/A OAI22X1_43/B gnd AOI21X1_82/C vdd
+ OAI22X1
XOAI22X1_26 INVX1_393/Y OAI22X1_43/B INVX8_12/Y OAI22X1_9/A gnd OAI22X1_26/Y vdd OAI22X1
XOAI22X1_37 OAI22X1_37/A OAI22X1_37/B NOR2X1_301/Y NOR2X1_269/A gnd NOR2X1_302/B vdd
+ OAI22X1
XOAI22X1_48 INVX2_76/Y INVX1_501/A INVX1_575/Y BUFX2_90/A gnd OAI22X1_48/Y vdd OAI22X1
XOAI22X1_59 INVX1_751/Y OAI22X1_58/B OAI22X1_58/C INVX1_752/Y gnd OAI22X1_59/Y vdd
+ OAI22X1
XOAI21X1_432 NOR2X1_191/Y NOR2X1_192/Y BUFX4_229/Y gnd OAI21X1_433/C vdd OAI21X1
XOAI21X1_421 NAND2X1_399/Y INVX2_54/Y OAI21X1_421/C gnd NAND2X1_406/B vdd OAI21X1
XOAI21X1_410 OAI21X1_410/A INVX8_5/A OAI21X1_410/C gnd MUX2X1_28/B vdd OAI21X1
XOAI21X1_443 INVX8_3/A NOR2X1_271/B OAI21X1_443/C gnd AOI21X1_68/B vdd OAI21X1
XOAI21X1_454 INVX2_52/Y INVX8_5/A INVX8_4/A gnd OAI21X1_454/Y vdd OAI21X1
XOAI21X1_465 AND2X2_34/Y OAI22X1_17/D AOI21X1_77/Y gnd AOI22X1_83/C vdd OAI21X1
XOAI21X1_498 INVX8_4/A INVX1_383/Y OAI21X1_498/C gnd INVX1_384/A vdd OAI21X1
XOAI21X1_487 NOR2X1_232/A NOR2X1_147/Y NOR2X1_228/B gnd NAND2X1_460/A vdd OAI21X1
XOAI21X1_476 INVX8_7/A INVX4_5/A OR2X2_42/A gnd AOI21X1_89/A vdd OAI21X1
XINVX1_507 INVX1_507/A gnd INVX1_507/Y vdd INVX1
XINVX1_518 INVX1_591/A gnd INVX1_518/Y vdd INVX1
XINVX1_529 INVX1_529/A gnd INVX1_529/Y vdd INVX1
XDFFPOSX1_390 INVX1_450/A CLKBUF1_37/Y OAI21X1_47/Y gnd vdd DFFPOSX1
XFILL_8_0_1 gnd vdd FILL
XNAND2X1_460 NAND2X1_460/A BUFX4_91/Y gnd NAND2X1_460/Y vdd NAND2X1
XNAND2X1_471 BUFX4_227/Y AOI21X1_93/Y gnd OAI21X1_505/C vdd NAND2X1
XNAND2X1_482 BUFX4_54/Y NAND2X1_482/B gnd NAND2X1_482/Y vdd NAND2X1
XNAND2X1_493 INVX8_7/A AND2X2_43/A gnd OAI21X1_537/A vdd NAND2X1
XFILL_36_7_0 gnd vdd FILL
XOAI21X1_81 INVX1_82/Y BUFX4_157/Y NAND2X1_83/Y gnd OAI21X1_81/Y vdd OAI21X1
XOAI21X1_70 INVX1_71/Y BUFX4_158/Y OAI21X1_70/C gnd OAI21X1_70/Y vdd OAI21X1
XOAI21X1_92 INVX1_93/Y BUFX4_159/Y NAND2X1_94/Y gnd OAI21X1_92/Y vdd OAI21X1
XAOI22X1_106 MUX2X1_54/A INVX2_55/A INVX1_425/Y INVX8_3/A gnd MUX2X1_53/B vdd AOI22X1
XAOI22X1_128 AOI22X1_128/A OR2X2_56/Y NAND2X1_941/Y NAND2X1_940/Y gnd AND2X2_83/B
+ vdd AOI22X1
XAOI22X1_117 OAI22X1_49/A INVX4_11/A BUFX4_262/Y OR2X2_52/B gnd OAI21X1_893/C vdd
+ AOI22X1
XAOI22X1_139 data_memory_interface_data[2] BUFX4_107/Y OAI21X1_989/Y BUFX4_9/Y gnd
+ OAI21X1_990/C vdd AOI22X1
XFILL_2_7_0 gnd vdd FILL
XFILL_27_7_0 gnd vdd FILL
XOAI21X1_240 AOI21X1_13/C OAI21X1_237/Y OAI21X1_239/Y gnd INVX1_252/A vdd OAI21X1
XFILL_10_6_0 gnd vdd FILL
XOAI21X1_251 INVX2_11/Y XNOR2X1_28/A NAND3X1_83/A gnd NAND2X1_148/B vdd OAI21X1
XOAI21X1_262 OR2X2_11/Y NOR2X1_50/A INVX1_269/Y gnd INVX1_270/A vdd OAI21X1
XOAI21X1_273 NOR2X1_51/B NOR2X1_51/A INVX1_287/Y gnd AOI21X1_32/B vdd OAI21X1
XINVX1_326 NOR2X1_96/Y gnd INVX1_326/Y vdd INVX1
XOAI21X1_295 INVX1_322/Y INVX4_4/A OAI21X1_295/C gnd MUX2X1_44/A vdd OAI21X1
XOAI21X1_284 INVX1_306/Y INVX4_4/A NAND2X1_198/Y gnd INVX4_3/A vdd OAI21X1
XINVX1_304 OR2X2_54/A gnd INVX1_304/Y vdd INVX1
XINVX1_315 INVX1_315/A gnd INVX1_315/Y vdd INVX1
XINVX1_337 INVX1_681/A gnd INVX1_337/Y vdd INVX1
XAND2X2_40 AND2X2_40/A BUFX4_84/Y gnd AND2X2_40/Y vdd AND2X2
XINVX1_348 INVX1_348/A gnd INVX1_348/Y vdd INVX1
XINVX1_359 INVX1_685/A gnd INVX1_359/Y vdd INVX1
XAND2X2_62 AND2X2_62/A AND2X2_62/B gnd AND2X2_62/Y vdd AND2X2
XAND2X2_51 AND2X2_51/A INVX1_408/A gnd AND2X2_51/Y vdd AND2X2
XAND2X2_73 OR2X2_25/B AND2X2_70/B gnd AND2X2_73/Y vdd AND2X2
XAND2X2_95 AND2X2_95/A AND2X2_95/B gnd AND2X2_95/Y vdd AND2X2
XAND2X2_84 MUX2X1_1/B INVX2_86/A gnd AND2X2_84/Y vdd AND2X2
XNAND2X1_290 AOI22X1_82/A OAI21X1_463/A gnd INVX1_378/A vdd NAND2X1
XFILL_18_7_0 gnd vdd FILL
XNAND2X1_1018 data_memory_interface_data[23] OAI21X1_981/B gnd NAND2X1_1018/Y vdd
+ NAND2X1
XDFFPOSX1_18 AOI22X1_18/D CLKBUF1_2/Y DFFPOSX1_18/D gnd vdd DFFPOSX1
XNAND2X1_1007 BUFX2_82/A BUFX4_115/Y gnd OAI21X1_972/C vdd NAND2X1
XNAND2X1_1029 INVX1_730/A BUFX4_254/Y gnd NAND3X1_362/B vdd NAND2X1
XDFFPOSX1_29 AOI22X1_29/D CLKBUF1_40/Y DFFPOSX1_29/D gnd vdd DFFPOSX1
XCLKBUF1_60 BUFX4_2/Y gnd CLKBUF1_60/Y vdd CLKBUF1
XFILL_42_5_0 gnd vdd FILL
XINVX1_101 INVX1_101/A gnd INVX1_101/Y vdd INVX1
XINVX1_123 INVX1_123/A gnd INVX1_123/Y vdd INVX1
XINVX1_112 INVX1_112/A gnd INVX1_112/Y vdd INVX1
XINVX1_134 BUFX2_91/A gnd AOI22X1_3/D vdd INVX1
XINVX1_156 instruction_memory_interface_data[0] gnd INVX1_156/Y vdd INVX1
XINVX1_145 INVX1_145/A gnd NOR3X1_8/B vdd INVX1
XINVX1_167 instruction_memory_interface_data[11] gnd NOR3X1_26/B vdd INVX1
XINVX1_189 INVX1_189/A gnd NOR2X1_9/A vdd INVX1
XINVX1_178 instruction_memory_interface_data[22] gnd INVX1_178/Y vdd INVX1
XFILL_34_3 gnd vdd FILL
XFILL_33_5_0 gnd vdd FILL
XAOI21X1_105 INVX8_7/A INVX1_391/Y OR2X2_31/Y gnd AOI21X1_106/B vdd AOI21X1
XAOI21X1_116 BUFX4_79/Y OAI22X1_27/Y AOI21X1_116/C gnd NAND3X1_135/C vdd AOI21X1
XAOI21X1_138 BUFX4_54/Y INVX2_66/Y BUFX4_176/Y gnd AOI21X1_139/B vdd AOI21X1
XAOI21X1_127 AOI22X1_70/B BUFX4_189/Y OAI22X1_36/Y gnd AOI21X1_127/Y vdd AOI21X1
XAOI21X1_149 INVX8_3/A NOR2X1_315/A INVX8_7/A gnd AOI21X1_149/Y vdd AOI21X1
XINVX1_690 INVX1_690/A gnd INVX1_690/Y vdd INVX1
XNAND3X1_109 NAND2X1_391/Y NAND2X1_363/Y NOR2X1_200/Y gnd INVX1_67/A vdd NAND3X1
XFILL_24_5_0 gnd vdd FILL
XFILL_7_6_0 gnd vdd FILL
XFILL_15_5_0 gnd vdd FILL
XDFFPOSX1_208 INVX1_720/A CLKBUF1_22/Y INVX1_454/A gnd vdd DFFPOSX1
XDFFPOSX1_219 AOI22X1_169/C CLKBUF1_8/Y INVX2_80/A gnd vdd DFFPOSX1
XNOR3X1_29 NOR3X1_3/A INVX1_170/Y BUFX4_49/Y gnd NOR3X1_29/Y vdd NOR3X1
XNOR3X1_18 INVX4_1/A INVX1_158/Y BUFX4_45/Y gnd NOR3X1_18/Y vdd NOR3X1
XBUFX4_240 AND2X2_8/Y gnd OR2X2_3/B vdd BUFX4
XNOR2X1_300 NOR2X1_300/A NOR2X1_300/B gnd NOR2X1_300/Y vdd NOR2X1
XBUFX4_262 BUFX4_262/A gnd BUFX4_262/Y vdd BUFX4
XBUFX4_273 NAND3X1_1/Y gnd BUFX4_273/Y vdd BUFX4
XBUFX4_251 BUFX4_253/A gnd BUFX4_251/Y vdd BUFX4
XNOR2X1_311 OR2X2_40/A NOR2X1_311/B gnd NOR3X1_57/B vdd NOR2X1
XNOR2X1_322 INVX8_3/A INVX1_425/A gnd NOR2X1_322/Y vdd NOR2X1
XNOR2X1_333 INVX2_29/A INVX2_30/Y gnd NOR2X1_333/Y vdd NOR2X1
XNOR2X1_344 INVX8_7/A NOR2X1_344/B gnd NOR2X1_344/Y vdd NOR2X1
XNOR2X1_355 NOR2X1_354/Y NOR2X1_355/B gnd NOR2X1_355/Y vdd NOR2X1
XNOR2X1_377 INVX2_6/A INVX1_437/Y gnd NOR2X1_377/Y vdd NOR2X1
XNOR2X1_366 INVX2_22/A NOR2X1_366/B gnd NOR2X1_366/Y vdd NOR2X1
XNOR2X1_388 BUFX2_55/A NOR3X1_65/Y gnd NOR2X1_388/Y vdd NOR2X1
XNOR2X1_399 XOR2X1_10/Y XOR2X1_11/Y gnd AND2X2_79/B vdd NOR2X1
XOAI21X1_806 BUFX4_177/Y INVX1_459/Y NAND2X1_629/Y gnd OAI21X1_806/Y vdd OAI21X1
XOAI21X1_817 INVX8_13/A BUFX2_41/A OAI21X1_817/C gnd OAI21X1_163/C vdd OAI21X1
XOAI21X1_839 NOR3X1_66/C INVX1_478/Y INVX8_13/Y gnd OAI21X1_839/Y vdd OAI21X1
XOAI21X1_828 NAND2X1_654/Y INVX1_474/Y INVX8_13/Y gnd OAI21X1_829/A vdd OAI21X1
XNAND2X1_801 NAND2X1_799/Y NAND2X1_801/B gnd NAND2X1_31/B vdd NAND2X1
XNAND2X1_812 OAI21X1_65/Y BUFX4_59/Y gnd NAND2X1_812/Y vdd NAND2X1
XNAND2X1_823 INVX1_578/Y BUFX4_98/Y gnd NAND3X1_263/C vdd NAND2X1
XNAND2X1_834 OAI21X1_70/Y BUFX4_63/Y gnd NAND2X1_834/Y vdd NAND2X1
XNAND2X1_845 NAND2X1_843/Y NAND2X1_845/B gnd NAND2X1_41/B vdd NAND2X1
XNAND2X1_867 OAI21X1_81/Y BUFX4_60/Y gnd NAND2X1_867/Y vdd NAND2X1
XNAND2X1_878 NAND2X1_876/Y NAND2X1_878/B gnd NAND2X1_52/B vdd NAND2X1
XNAND2X1_889 INVX1_622/Y BUFX4_95/Y gnd NAND3X1_307/C vdd NAND2X1
XNAND2X1_856 INVX1_600/Y BUFX4_96/Y gnd NAND3X1_285/C vdd NAND2X1
XNAND3X1_40 NAND3X1_40/A BUFX4_110/Y BUFX4_138/Y gnd NAND3X1_41/B vdd NAND3X1
XNAND3X1_73 NOR2X1_13/A NOR2X1_11/Y AND2X2_6/A gnd NAND3X1_73/Y vdd NAND3X1
XNAND3X1_51 BUFX4_73/Y NAND3X1_51/B NAND3X1_51/C gnd NAND3X1_51/Y vdd NAND3X1
XNAND3X1_84 INVX1_268/Y NAND3X1_84/B NAND3X1_84/C gnd NAND3X1_84/Y vdd NAND3X1
XNAND3X1_62 NAND3X1_62/A AND2X2_2/B AND2X2_2/A gnd NAND3X1_63/B vdd NAND3X1
XNAND3X1_95 INVX2_23/Y INVX2_20/Y NOR2X1_162/Y gnd NOR2X1_165/A vdd NAND3X1
XNOR2X1_40 INVX2_13/Y NOR2X1_40/B gnd NOR2X1_40/Y vdd NOR2X1
XNOR2X1_51 NOR2X1_51/A NOR2X1_51/B gnd XOR2X1_6/A vdd NOR2X1
XNOR2X1_62 NOR2X1_62/A INVX1_291/Y gnd NOR2X1_62/Y vdd NOR2X1
XNOR2X1_73 INVX2_16/A INVX2_17/A gnd NOR2X1_73/Y vdd NOR2X1
XNOR2X1_95 INVX2_35/Y MUX2X1_42/B gnd NOR2X1_95/Y vdd NOR2X1
XNOR2X1_84 INVX2_20/Y INVX2_21/Y gnd NOR2X1_85/B vdd NOR2X1
XFILL_30_3_0 gnd vdd FILL
XNAND2X1_108 INVX1_150/A INVX1_149/A gnd OR2X2_5/B vdd NAND2X1
XNAND2X1_119 MUX2X1_13/A BUFX4_233/Y gnd AOI21X1_5/A vdd NAND2X1
XNAND2X1_6 BUFX4_19/Y NAND2X1_6/B gnd OAI21X1_6/C vdd NAND2X1
XFILL_38_4_0 gnd vdd FILL
XNOR2X1_141 BUFX4_213/Y MUX2X1_12/Y gnd AOI22X1_79/D vdd NOR2X1
XNOR2X1_152 NOR2X1_152/A OAI22X1_12/Y gnd NOR2X1_152/Y vdd NOR2X1
XNOR2X1_130 INVX2_51/A INVX1_358/A gnd AND2X2_26/A vdd NOR2X1
XNOR2X1_185 INVX2_56/A NOR2X1_185/B gnd BUFX4_152/A vdd NOR2X1
XNOR2X1_174 AND2X2_93/B INVX2_49/A gnd AND2X2_25/A vdd NOR2X1
XNOR2X1_163 INVX1_307/A NOR2X1_80/A gnd NOR2X1_163/Y vdd NOR2X1
XNOR2X1_196 NAND3X1_94/A NOR2X1_195/Y gnd NOR2X1_196/Y vdd NOR2X1
XOAI21X1_614 OAI21X1_520/A BUFX4_51/Y OAI21X1_614/C gnd NAND2X1_540/B vdd OAI21X1
XOAI21X1_603 NOR2X1_253/B OAI21X1_603/B AOI21X1_144/Y gnd AOI21X1_185/B vdd OAI21X1
XFILL_21_3_0 gnd vdd FILL
XOAI21X1_636 MUX2X1_50/A INVX2_55/Y BUFX4_125/Y gnd AOI21X1_152/C vdd OAI21X1
XOAI21X1_625 INVX2_35/A MUX2X1_42/B BUFX4_190/Y gnd OAI21X1_625/Y vdd OAI21X1
XOAI21X1_647 AND2X2_51/Y NOR2X1_325/B OAI21X1_647/C gnd OAI21X1_647/Y vdd OAI21X1
XOAI21X1_658 AND2X2_54/A INVX4_10/Y INVX8_11/Y gnd OAI21X1_667/B vdd OAI21X1
XOAI21X1_669 INVX1_406/A NOR2X1_336/A INVX1_417/A gnd AOI21X1_168/B vdd OAI21X1
XXNOR2X1_19 XNOR2X1_19/A NOR2X1_33/B gnd XNOR2X1_19/Y vdd XNOR2X1
XNAND2X1_620 INVX2_12/A BUFX4_265/Y gnd NAND2X1_620/Y vdd NAND2X1
XNAND2X1_642 BUFX4_245/Y XNOR2X1_10/Y gnd OAI21X1_818/C vdd NAND2X1
XNAND2X1_664 BUFX4_245/Y XNOR2X1_35/Y gnd OAI21X1_838/C vdd NAND2X1
XNAND2X1_653 BUFX2_47/A XOR2X1_8/B gnd OR2X2_46/A vdd NAND2X1
XINVX1_21 gnd gnd INVX1_21/Y vdd INVX1
XINVX1_10 gnd gnd INVX1_10/Y vdd INVX1
XNAND2X1_631 INVX1_279/A BUFX4_266/Y gnd NAND2X1_631/Y vdd NAND2X1
XINVX1_32 gnd gnd INVX1_32/Y vdd INVX1
XNAND2X1_675 INVX8_13/A XNOR2X1_40/Y gnd OAI21X1_849/C vdd NAND2X1
XNAND2X1_686 BUFX2_63/A BUFX2_64/A gnd NOR3X1_66/B vdd NAND2X1
XINVX1_76 INVX1_76/A gnd INVX1_76/Y vdd INVX1
XINVX1_65 INVX1_65/A gnd INVX1_65/Y vdd INVX1
XINVX1_43 gnd gnd INVX1_43/Y vdd INVX1
XINVX1_54 gnd gnd INVX1_54/Y vdd INVX1
XNAND2X1_697 INVX2_1/A INVX1_495/Y gnd NAND3X1_186/A vdd NAND2X1
XBUFX2_18 BUFX2_18/A gnd data_memory_interface_address[17] vdd BUFX2
XFILL_4_4_0 gnd vdd FILL
XFILL_29_4_0 gnd vdd FILL
XINVX1_98 INVX1_98/A gnd INVX1_98/Y vdd INVX1
XINVX1_87 INVX1_87/A gnd INVX1_87/Y vdd INVX1
XBUFX2_29 BUFX2_29/A gnd data_memory_interface_address[28] vdd BUFX2
XDFFPOSX1_6 INVX1_189/A CLKBUF1_60/Y NOR2X1_3/A gnd vdd DFFPOSX1
XFILL_12_3_0 gnd vdd FILL
XNOR2X1_9 NOR2X1_9/A NOR2X1_9/B gnd AND2X2_6/B vdd NOR2X1
XNAND3X1_281 BUFX4_121/Y NAND3X1_280/Y NAND3X1_281/C gnd NAND2X1_851/B vdd NAND3X1
XNAND3X1_270 INVX1_587/Y BUFX4_99/Y BUFX4_167/Y gnd NAND3X1_271/B vdd NAND3X1
XNAND3X1_292 INVX1_609/Y BUFX4_103/Y BUFX4_164/Y gnd NAND3X1_293/B vdd NAND3X1
XAOI21X1_19 AOI21X1_8/A AOI21X1_8/B INVX1_256/Y gnd AOI21X1_19/Y vdd AOI21X1
XOAI22X1_38 OAI22X1_38/A OAI22X1_38/B NOR2X1_303/Y NOR2X1_293/A gnd NOR2X1_304/B vdd
+ OAI22X1
XOAI22X1_16 OR2X2_29/B NOR2X1_327/B INVX1_379/A OAI22X1_27/A gnd AOI22X1_84/C vdd
+ OAI22X1
XOAI22X1_27 OAI22X1_27/A OR2X2_42/B OR2X2_33/Y OR2X2_29/B gnd OAI22X1_27/Y vdd OAI22X1
XOAI22X1_49 OAI22X1_49/A OAI22X1_49/B OAI22X1_49/C INVX1_641/Y gnd OAI22X1_49/Y vdd
+ OAI22X1
XOAI21X1_400 BUFX4_42/Y MUX2X1_8/Y NAND2X1_385/Y gnd INVX1_367/A vdd OAI21X1
XOAI21X1_411 INVX8_5/A OAI21X1_411/B OAI21X1_411/C gnd OAI21X1_412/A vdd OAI21X1
XOAI21X1_422 NOR2X1_206/Y NOR2X1_205/Y BUFX4_124/Y gnd NAND2X1_407/A vdd OAI21X1
XOAI21X1_444 AOI21X1_68/B BUFX4_176/Y INVX8_7/A gnd AND2X2_31/A vdd OAI21X1
XOAI21X1_466 OAI22X1_10/Y AOI21X1_63/Y AOI21X1_78/Y gnd AOI21X1_79/B vdd OAI21X1
XOAI21X1_455 OAI21X1_506/B INVX8_4/A OAI21X1_454/Y gnd OR2X2_26/A vdd OAI21X1
XOAI21X1_433 INVX1_368/Y BUFX4_229/Y OAI21X1_433/C gnd MUX2X1_33/A vdd OAI21X1
XOAI21X1_499 INVX8_3/A MUX2X1_33/Y OAI21X1_499/C gnd AOI21X1_89/B vdd OAI21X1
XOAI21X1_477 AOI21X1_77/Y AND2X2_34/Y AOI22X1_88/D gnd OR2X2_28/A vdd OAI21X1
XOAI21X1_488 AOI21X1_124/B BUFX4_57/Y INVX4_7/A gnd OAI21X1_489/B vdd OAI21X1
XINVX1_508 INVX1_581/A gnd INVX1_508/Y vdd INVX1
XINVX1_519 INVX1_592/A gnd INVX1_519/Y vdd INVX1
XDFFPOSX1_380 OR2X2_61/B CLKBUF1_37/Y OAI21X1_37/Y gnd vdd DFFPOSX1
XDFFPOSX1_391 INVX1_451/A CLKBUF1_29/Y OAI21X1_48/Y gnd vdd DFFPOSX1
XNAND2X1_461 AOI22X1_87/A MUX2X1_29/Y gnd NAND2X1_462/A vdd NAND2X1
XNAND2X1_472 BUFX4_215/Y NAND2X1_472/B gnd NAND2X1_472/Y vdd NAND2X1
XNAND2X1_450 INVX4_4/Y INVX1_344/Y gnd AOI21X1_85/B vdd NAND2X1
XNAND2X1_483 INVX8_7/A AND2X2_40/A gnd OAI21X1_523/C vdd NAND2X1
XNAND2X1_494 INVX1_360/Y NOR2X1_265/Y gnd NAND2X1_494/Y vdd NAND2X1
XFILL_36_7_1 gnd vdd FILL
XFILL_35_2_0 gnd vdd FILL
XOAI21X1_60 INVX1_60/Y BUFX4_26/Y OAI21X1_60/C gnd OAI21X1_60/Y vdd OAI21X1
XOAI21X1_71 INVX1_72/Y BUFX4_159/Y NAND2X1_73/Y gnd OAI21X1_71/Y vdd OAI21X1
XOAI21X1_82 INVX1_83/Y BUFX4_161/Y NAND2X1_84/Y gnd OAI21X1_82/Y vdd OAI21X1
XOAI21X1_93 INVX1_94/Y BUFX4_156/Y NAND2X1_95/Y gnd OAI21X1_93/Y vdd OAI21X1
XAOI22X1_107 INVX2_55/A OAI22X1_42/Y NOR2X1_328/Y INVX8_3/A gnd MUX2X1_55/B vdd AOI22X1
XAOI22X1_118 OAI22X1_49/A INVX4_11/A BUFX4_262/Y BUFX2_90/A gnd OAI21X1_894/C vdd
+ AOI22X1
XAOI22X1_129 AOI22X1_129/A OR2X2_57/Y NAND2X1_948/Y NAND2X1_947/Y gnd NAND3X1_341/B
+ vdd AOI22X1
XFILL_2_7_1 gnd vdd FILL
XFILL_27_7_1 gnd vdd FILL
XFILL_1_2_0 gnd vdd FILL
XFILL_26_2_0 gnd vdd FILL
XOAI21X1_241 NOR2X1_42/A INVX1_244/A INVX1_252/Y gnd NOR2X1_30/A vdd OAI21X1
XFILL_10_6_1 gnd vdd FILL
XOAI21X1_230 AND2X2_13/Y OAI21X1_230/B OR2X2_9/Y gnd NAND3X1_78/C vdd OAI21X1
XOAI21X1_252 NOR2X1_36/Y NOR2X1_39/B NAND2X1_148/Y gnd XNOR2X1_32/A vdd OAI21X1
XOAI21X1_263 AOI21X1_26/Y OAI21X1_276/B AND2X2_14/Y gnd OAI21X1_263/Y vdd OAI21X1
XOAI21X1_274 XOR2X1_7/B INVX1_284/Y INVX1_286/Y gnd AOI21X1_31/C vdd OAI21X1
XOAI21X1_296 INVX4_4/Y AOI22X1_57/A OAI21X1_296/C gnd NOR2X1_160/B vdd OAI21X1
XINVX1_316 OR2X2_15/Y gnd INVX1_316/Y vdd INVX1
XOAI21X1_285 INVX1_308/Y INVX4_4/A NAND2X1_199/Y gnd INVX2_50/A vdd OAI21X1
XINVX1_305 INVX1_305/A gnd INVX1_305/Y vdd INVX1
XINVX1_327 INVX1_327/A gnd INVX1_327/Y vdd INVX1
XINVX1_338 OR2X2_62/A gnd INVX1_338/Y vdd INVX1
XAND2X2_41 AND2X2_41/A INVX2_59/Y gnd AND2X2_41/Y vdd AND2X2
XAND2X2_30 MUX2X1_14/Y MUX2X1_47/S gnd AND2X2_30/Y vdd AND2X2
XINVX1_349 INVX1_349/A gnd INVX1_349/Y vdd INVX1
XAND2X2_52 AND2X2_52/A AND2X2_52/B gnd AND2X2_52/Y vdd AND2X2
XAND2X2_63 AND2X2_63/A NOR3X1_56/Y gnd AND2X2_63/Y vdd AND2X2
XAND2X2_74 AND2X2_74/A INVX2_55/A gnd AND2X2_74/Y vdd AND2X2
XFILL_9_3_0 gnd vdd FILL
XAND2X2_85 MUX2X1_2/B INVX1_454/A gnd AND2X2_85/Y vdd AND2X2
XAND2X2_96 MUX2X1_7/B OR2X2_58/B gnd AND2X2_96/Y vdd AND2X2
XNAND2X1_280 INVX4_4/A INVX1_247/A gnd OAI21X1_321/C vdd NAND2X1
XNAND2X1_291 INVX1_342/A MUX2X1_15/Y gnd AOI22X1_89/B vdd NAND2X1
XFILL_18_7_1 gnd vdd FILL
XFILL_17_2_0 gnd vdd FILL
XNAND2X1_1008 BUFX2_83/A BUFX4_115/Y gnd OAI21X1_973/C vdd NAND2X1
XDFFPOSX1_19 AOI22X1_19/D CLKBUF1_61/Y DFFPOSX1_19/D gnd vdd DFFPOSX1
XNAND2X1_1019 INVX2_88/A INVX2_90/A gnd OAI22X1_60/D vdd NAND2X1
XCLKBUF1_50 BUFX4_7/Y gnd CLKBUF1_50/Y vdd CLKBUF1
XCLKBUF1_61 BUFX4_4/Y gnd CLKBUF1_61/Y vdd CLKBUF1
XFILL_42_5_1 gnd vdd FILL
XFILL_41_0_0 gnd vdd FILL
XINVX1_124 INVX1_124/A gnd INVX1_124/Y vdd INVX1
XINVX1_113 INVX1_113/A gnd INVX1_113/Y vdd INVX1
XINVX1_102 INVX1_102/A gnd INVX1_102/Y vdd INVX1
XINVX1_168 instruction_memory_interface_data[12] gnd INVX1_168/Y vdd INVX1
XINVX1_146 BUFX2_84/A gnd NOR3X1_9/B vdd INVX1
XINVX1_157 instruction_memory_interface_data[1] gnd INVX1_157/Y vdd INVX1
XINVX1_135 OR2X2_50/B gnd AOI22X1_4/D vdd INVX1
XINVX1_179 instruction_memory_interface_data[23] gnd NOR3X1_38/B vdd INVX1
XFILL_33_5_1 gnd vdd FILL
XAOI21X1_106 OAI21X1_536/Y AOI21X1_106/B OAI22X1_25/Y gnd NAND3X1_127/B vdd AOI21X1
XFILL_32_0_0 gnd vdd FILL
XAOI21X1_139 AOI21X1_136/Y AOI21X1_139/B NOR2X1_299/Y gnd OAI21X1_599/B vdd AOI21X1
XAOI21X1_128 INVX4_6/Y MUX2X1_38/Y OR2X2_35/Y gnd NAND3X1_139/C vdd AOI21X1
XAOI21X1_117 NOR2X1_281/A OAI21X1_565/B BUFX4_274/Y gnd AOI21X1_117/Y vdd AOI21X1
XINVX1_680 INVX1_449/A gnd INVX1_680/Y vdd INVX1
XINVX1_691 INVX1_691/A gnd INVX1_691/Y vdd INVX1
XFILL_24_5_1 gnd vdd FILL
XFILL_23_0_0 gnd vdd FILL
XINVX4_10 INVX4_10/A gnd INVX4_10/Y vdd INVX4
XFILL_7_6_1 gnd vdd FILL
XFILL_6_1_0 gnd vdd FILL
XFILL_15_5_1 gnd vdd FILL
XFILL_14_0_0 gnd vdd FILL
XDFFPOSX1_209 INVX1_721/A CLKBUF1_38/Y INVX2_86/A gnd vdd DFFPOSX1
XBUFX4_230 INVX8_5/Y gnd MUX2X1_47/S vdd BUFX4
XNOR3X1_19 NOR3X1_3/A INVX1_159/Y BUFX4_45/Y gnd NOR3X1_19/Y vdd NOR3X1
XNOR2X1_301 INVX2_43/Y NOR2X1_123/B gnd NOR2X1_301/Y vdd NOR2X1
XBUFX4_241 BUFX4_242/A gnd BUFX4_241/Y vdd BUFX4
XBUFX4_263 BUFX4_262/A gnd BUFX4_263/Y vdd BUFX4
XBUFX4_252 BUFX4_253/A gnd BUFX4_252/Y vdd BUFX4
XBUFX4_274 BUFX4_276/A gnd BUFX4_274/Y vdd BUFX4
XNOR2X1_312 INVX2_37/A MUX2X1_42/A gnd NOR2X1_312/Y vdd NOR2X1
XNOR2X1_334 INVX4_9/Y MUX2X1_38/A gnd NOR2X1_334/Y vdd NOR2X1
XNOR2X1_323 INVX4_9/Y NOR2X1_323/B gnd NOR2X1_323/Y vdd NOR2X1
XNOR2X1_345 AND2X2_56/B OR2X2_30/A gnd NOR2X1_345/Y vdd NOR2X1
XNOR2X1_356 NOR2X1_356/A NOR2X1_356/B gnd INVX1_423/A vdd NOR2X1
XNOR2X1_367 INVX2_20/A INVX2_21/Y gnd NOR2X1_367/Y vdd NOR2X1
XFILL_32_1 gnd vdd FILL
XNOR2X1_389 OR2X2_47/A OR2X2_47/B gnd NOR2X1_389/Y vdd NOR2X1
XNOR2X1_378 NOR2X1_377/Y NOR2X1_378/B gnd NOR2X1_378/Y vdd NOR2X1
XOAI21X1_818 OR2X2_45/Y NOR2X1_380/Y OAI21X1_818/C gnd OAI21X1_164/C vdd OAI21X1
XOAI21X1_829 OAI21X1_829/A AOI21X1_215/Y OAI21X1_829/C gnd OAI21X1_829/Y vdd OAI21X1
XOAI21X1_807 BUFX4_178/Y INVX1_460/Y NAND2X1_630/Y gnd OAI21X1_807/Y vdd OAI21X1
XNAND2X1_802 OAI21X1_96/Y BUFX4_131/Y gnd NAND2X1_802/Y vdd NAND2X1
XNAND2X1_813 AND2X2_80/B AND2X2_80/A gnd BUFX4_122/A vdd NAND2X1
XNAND2X1_824 NAND2X1_822/Y NAND2X1_824/B gnd NAND2X1_34/B vdd NAND2X1
XNAND2X1_846 OAI21X1_74/Y BUFX4_62/Y gnd NAND2X1_846/Y vdd NAND2X1
XNAND2X1_835 INVX1_586/Y BUFX4_97/Y gnd NAND3X1_271/C vdd NAND2X1
XNAND2X1_857 NAND2X1_855/Y NAND2X1_857/B gnd NAND2X1_45/B vdd NAND2X1
XNAND2X1_879 OAI21X1_85/Y BUFX4_62/Y gnd NAND2X1_879/Y vdd NAND2X1
XNAND2X1_868 INVX1_608/Y BUFX4_98/Y gnd NAND3X1_293/C vdd NAND2X1
XNAND3X1_41 BUFX4_72/Y NAND3X1_41/B NAND3X1_41/C gnd NAND3X1_41/Y vdd NAND3X1
XNAND3X1_30 NAND3X1_30/A BUFX4_110/Y BUFX4_138/Y gnd NAND3X1_30/Y vdd NAND3X1
XNAND3X1_52 NAND3X1_52/A BUFX4_114/Y BUFX4_136/Y gnd NAND3X1_53/B vdd NAND3X1
XNAND3X1_63 BUFX4_76/Y NAND3X1_63/B NAND3X1_63/C gnd NAND3X1_63/Y vdd NAND3X1
XNAND3X1_74 NOR2X1_20/Y NAND3X1_74/B NOR2X1_21/Y gnd NAND3X1_74/Y vdd NAND3X1
XNOR2X1_30 NOR2X1_30/A NOR2X1_30/B gnd NOR2X1_35/B vdd NOR2X1
XNAND3X1_85 NAND3X1_85/A AND2X2_16/Y NAND3X1_85/C gnd NOR2X1_51/A vdd NAND3X1
XNAND3X1_96 INVX1_303/Y INVX2_16/Y NOR2X1_163/Y gnd OR2X2_20/A vdd NAND3X1
XNOR2X1_41 INVX2_14/Y NOR2X1_41/B gnd NOR2X1_41/Y vdd NOR2X1
XNOR2X1_63 NOR2X1_62/Y INVX1_292/Y gnd INVX1_294/A vdd NOR2X1
XNOR2X1_52 INVX1_278/Y NOR2X1_52/B gnd INVX2_15/A vdd NOR2X1
XNOR2X1_96 INVX2_37/A NOR2X1_96/B gnd NOR2X1_96/Y vdd NOR2X1
XNOR2X1_74 NOR2X1_73/Y NOR2X1_72/Y gnd INVX2_18/A vdd NOR2X1
XNOR2X1_85 NOR2X1_85/A NOR2X1_85/B gnd INVX2_22/A vdd NOR2X1
XFILL_30_3_1 gnd vdd FILL
XNAND2X1_109 NOR2X1_14/Y NOR2X1_15/Y gnd NAND2X1_109/Y vdd NAND2X1
XNAND2X1_7 BUFX4_17/Y NAND2X1_7/B gnd OAI21X1_7/C vdd NAND2X1
XFILL_38_4_1 gnd vdd FILL
XNOR2X1_120 INVX2_42/Y MUX2X1_7/Y gnd OAI22X1_9/B vdd NOR2X1
XNOR2X1_142 AND2X2_22/Y INVX1_369/A gnd NAND3X1_94/A vdd NOR2X1
XNOR2X1_131 NOR2X1_131/A OR2X2_16/Y gnd OR2X2_44/A vdd NOR2X1
XNOR2X1_153 NOR2X1_153/A NAND3X1_93/Y gnd NOR2X1_153/Y vdd NOR2X1
XNOR2X1_164 INVX1_317/A INVX2_29/A gnd NAND3X1_97/C vdd NOR2X1
XNOR2X1_175 INVX2_48/A NOR2X1_175/B gnd NOR2X1_175/Y vdd NOR2X1
XNOR2X1_197 MUX2X1_47/S MUX2X1_14/Y gnd AOI21X1_69/C vdd NOR2X1
XNOR2X1_186 OR2X2_23/B OR2X2_23/A gnd NOR2X1_186/Y vdd NOR2X1
XOAI21X1_604 INVX2_67/A INVX1_329/A OAI21X1_604/C gnd NOR2X1_316/B vdd OAI21X1
XOAI21X1_615 BUFX4_126/Y NOR2X1_188/Y INVX1_400/A gnd NOR2X1_310/A vdd OAI21X1
XFILL_21_3_1 gnd vdd FILL
XOAI21X1_637 AOI22X1_80/D BUFX4_125/Y INVX2_65/A gnd NOR2X1_318/B vdd OAI21X1
XOAI21X1_648 NOR2X1_160/B INVX8_8/A OAI21X1_648/C gnd NAND2X1_564/B vdd OAI21X1
XOAI21X1_626 OR2X2_24/A OR2X2_24/B INVX1_403/Y gnd NAND3X1_143/A vdd OAI21X1
XOAI21X1_659 NOR2X1_325/B AND2X2_51/Y NOR2X1_324/Y gnd OAI21X1_659/Y vdd OAI21X1
XNAND2X1_610 INVX1_234/A BUFX4_264/Y gnd NAND2X1_610/Y vdd NAND2X1
XNAND2X1_621 INVX2_13/A BUFX4_267/Y gnd NAND2X1_621/Y vdd NAND2X1
XNAND2X1_643 INVX8_13/Y INVX1_471/A gnd NAND2X1_643/Y vdd NAND2X1
XNAND2X1_654 INVX1_473/Y NOR2X1_382/Y gnd NAND2X1_654/Y vdd NAND2X1
XINVX1_22 gnd gnd INVX1_22/Y vdd INVX1
XNAND2X1_632 INVX1_283/A BUFX4_266/Y gnd NAND2X1_632/Y vdd NAND2X1
XINVX1_11 gnd gnd INVX1_11/Y vdd INVX1
XINVX1_33 gnd gnd INVX1_33/Y vdd INVX1
XNAND2X1_665 BUFX2_53/A BUFX2_54/A gnd OR2X2_47/B vdd NAND2X1
XNAND2X1_676 BUFX2_59/A BUFX2_60/A gnd OR2X2_48/B vdd NAND2X1
XNAND2X1_687 BUFX4_241/Y XNOR2X1_46/Y gnd OAI21X1_859/C vdd NAND2X1
XINVX1_66 INVX1_66/A gnd INVX1_66/Y vdd INVX1
XINVX1_44 gnd gnd INVX1_44/Y vdd INVX1
XINVX1_55 gnd gnd INVX1_55/Y vdd INVX1
XFILL_4_4_1 gnd vdd FILL
XINVX1_88 INVX1_88/A gnd INVX1_88/Y vdd INVX1
XINVX1_77 INVX1_77/A gnd INVX1_77/Y vdd INVX1
XFILL_29_4_1 gnd vdd FILL
XINVX1_99 INVX2_89/A gnd INVX1_99/Y vdd INVX1
XNAND2X1_698 XOR2X1_1/A INVX2_73/Y gnd NAND3X1_186/B vdd NAND2X1
XBUFX2_19 BUFX2_19/A gnd data_memory_interface_address[18] vdd BUFX2
XDFFPOSX1_7 NOR2X1_11/A CLKBUF1_60/Y INVX2_89/A gnd vdd DFFPOSX1
XFILL_12_3_1 gnd vdd FILL
XNAND3X1_260 INVX1_576/Y BUFX4_102/Y BUFX4_168/Y gnd NAND3X1_260/Y vdd NAND3X1
XNAND3X1_271 BUFX4_123/Y NAND3X1_271/B NAND3X1_271/C gnd NAND2X1_836/B vdd NAND3X1
XNAND3X1_282 INVX1_599/Y BUFX4_101/Y BUFX4_166/Y gnd NAND3X1_283/B vdd NAND3X1
XNAND3X1_293 BUFX4_122/Y NAND3X1_293/B NAND3X1_293/C gnd NAND2X1_869/B vdd NAND3X1
XOAI22X1_39 OAI22X1_20/A OAI22X1_39/B AOI21X1_37/B OAI22X1_43/B gnd OAI22X1_39/Y vdd
+ OAI22X1
XOAI22X1_17 AOI21X1_88/C OAI22X1_17/B AND2X2_34/Y OAI22X1_17/D gnd NOR2X1_246/A vdd
+ OAI22X1
XOAI22X1_28 MUX2X1_26/Y INVX4_9/Y OAI22X1_14/C INVX8_3/A gnd OAI22X1_28/Y vdd OAI22X1
XOAI21X1_423 MUX2X1_21/Y INVX8_5/A NAND2X1_408/Y gnd NAND2X1_409/B vdd OAI21X1
XOAI21X1_401 INVX1_367/Y INVX8_5/A OAI21X1_399/Y gnd MUX2X1_27/A vdd OAI21X1
XOAI21X1_412 OAI21X1_412/A INVX8_4/A OAI21X1_412/C gnd AND2X2_44/A vdd OAI21X1
XOAI21X1_445 AND2X2_31/Y AOI21X1_68/Y OAI21X1_435/Y gnd NAND3X1_111/A vdd OAI21X1
XOAI21X1_434 BUFX4_215/Y INVX1_383/A NAND2X1_417/Y gnd NOR2X1_270/B vdd OAI21X1
XOAI21X1_456 MUX2X1_26/Y INVX8_3/A OAI21X1_456/C gnd AOI22X1_83/A vdd OAI21X1
XOAI21X1_478 AOI21X1_74/Y NOR2X1_246/A AOI21X1_86/Y gnd OAI21X1_480/B vdd OAI21X1
XOAI21X1_467 AOI21X1_74/Y NOR2X1_151/Y OAI21X1_463/A gnd AOI21X1_81/B vdd OAI21X1
XOAI21X1_489 NOR2X1_225/Y OAI21X1_489/B OAI21X1_489/C gnd NOR2X1_230/B vdd OAI21X1
XINVX1_509 INVX1_509/A gnd INVX1_509/Y vdd INVX1
XDFFPOSX1_370 OR2X2_55/A CLKBUF1_53/Y OAI21X1_27/Y gnd vdd DFFPOSX1
XDFFPOSX1_392 INVX1_452/A CLKBUF1_37/Y OAI21X1_49/Y gnd vdd DFFPOSX1
XDFFPOSX1_381 OR2X2_60/B CLKBUF1_22/Y OAI21X1_38/Y gnd vdd DFFPOSX1
XNAND2X1_462 NAND2X1_462/A AOI22X1_85/Y gnd NOR2X1_230/A vdd NAND2X1
XNAND2X1_451 INVX4_4/A INVX1_380/Y gnd AOI21X1_85/A vdd NAND2X1
XNAND2X1_440 BUFX4_53/Y OAI21X1_472/Y gnd OAI21X1_473/C vdd NAND2X1
XNAND2X1_473 BUFX4_54/Y AOI21X1_52/B gnd NAND2X1_473/Y vdd NAND2X1
XNAND2X1_484 INVX2_54/A AND2X2_40/Y gnd OAI21X1_524/C vdd NAND2X1
XNAND2X1_495 BUFX4_85/Y INVX1_391/A gnd OR2X2_40/B vdd NAND2X1
XOAI21X1_990 AOI21X1_260/Y OAI21X1_994/B OAI21X1_990/C gnd OAI21X1_990/Y vdd OAI21X1
XFILL_35_2_1 gnd vdd FILL
XOAI21X1_72 INVX1_73/Y BUFX4_157/Y NAND2X1_74/Y gnd OAI21X1_72/Y vdd OAI21X1
XOAI21X1_50 INVX1_50/Y BUFX4_26/Y OAI21X1_50/C gnd OAI21X1_50/Y vdd OAI21X1
XOAI21X1_61 INVX1_61/Y BUFX4_25/Y OAI21X1_61/C gnd OAI21X1_61/Y vdd OAI21X1
XOAI21X1_94 INVX1_95/Y BUFX4_156/Y OAI21X1_94/C gnd OAI21X1_94/Y vdd OAI21X1
XOAI21X1_83 INVX1_84/Y BUFX4_158/Y NAND2X1_85/Y gnd OAI21X1_83/Y vdd OAI21X1
XAOI22X1_108 INVX1_431/Y INVX8_12/A OR2X2_24/Y INVX2_28/A gnd AOI22X1_108/Y vdd AOI22X1
XAOI22X1_119 OAI22X1_49/A INVX4_11/A BUFX4_261/Y BUFX2_91/A gnd AOI22X1_119/Y vdd
+ AOI22X1
XFILL_1_2_1 gnd vdd FILL
XFILL_26_2_1 gnd vdd FILL
XOAI21X1_231 AND2X2_10/Y NOR2X1_24/Y AND2X2_9/Y gnd NOR3X1_49/C vdd OAI21X1
XOAI21X1_220 BUFX4_145/Y INVX1_218/Y AOI22X1_35/Y gnd OAI21X1_220/Y vdd OAI21X1
XOAI21X1_242 NOR2X1_30/B NOR2X1_30/A XNOR2X1_17/Y gnd OAI21X1_242/Y vdd OAI21X1
XOAI21X1_253 NOR2X1_39/A NAND2X1_148/Y AOI21X1_22/Y gnd INVX1_263/A vdd OAI21X1
XOAI21X1_264 INVX1_272/Y NOR2X1_45/A OR2X2_12/Y gnd XNOR2X1_41/A vdd OAI21X1
XOAI21X1_297 INVX1_323/Y INVX4_4/A NAND2X1_222/Y gnd NOR2X1_94/B vdd OAI21X1
XINVX1_317 INVX1_317/A gnd NOR2X1_99/A vdd INVX1
XOAI21X1_275 XOR2X1_6/A INVX1_287/A INVX1_293/A gnd NOR2X1_59/B vdd OAI21X1
XINVX1_306 INVX1_306/A gnd INVX1_306/Y vdd INVX1
XOAI21X1_286 INVX1_309/Y INVX4_4/A NAND2X1_202/Y gnd INVX2_21/A vdd OAI21X1
XAND2X2_31 AND2X2_31/A AND2X2_31/B gnd AND2X2_31/Y vdd AND2X2
XINVX1_339 OR2X2_63/A gnd INVX1_339/Y vdd INVX1
XINVX1_328 INVX1_328/A gnd INVX1_328/Y vdd INVX1
XAND2X2_20 AND2X2_1/A AND2X2_1/B gnd AND2X2_20/Y vdd AND2X2
XAND2X2_53 NOR3X1_56/Y AND2X2_53/B gnd AND2X2_53/Y vdd AND2X2
XAND2X2_42 AND2X2_42/A AND2X2_42/B gnd AND2X2_42/Y vdd AND2X2
XAND2X2_64 AND2X2_64/A AND2X2_64/B gnd AND2X2_64/Y vdd AND2X2
XFILL_9_3_1 gnd vdd FILL
XAND2X2_75 BUFX2_41/A BUFX2_42/A gnd OR2X2_45/A vdd AND2X2
XAND2X2_86 AND2X2_86/A AND2X2_86/B gnd AND2X2_86/Y vdd AND2X2
XAND2X2_97 OR2X2_59/A OR2X2_59/B gnd AND2X2_97/Y vdd AND2X2
XNAND2X1_270 INVX8_4/A MUX2X1_21/B gnd AOI22X1_73/D vdd NAND2X1
XNAND2X1_281 INVX2_46/A MUX2X1_30/B gnd AOI22X1_74/C vdd NAND2X1
XNAND2X1_292 INVX2_46/A MUX2X1_16/Y gnd AOI22X1_89/C vdd NAND2X1
XFILL_17_2_1 gnd vdd FILL
XNAND2X1_1009 OAI21X1_966/C BUFX4_115/Y gnd OAI21X1_974/C vdd NAND2X1
XCLKBUF1_40 BUFX4_1/Y gnd CLKBUF1_40/Y vdd CLKBUF1
XCLKBUF1_51 BUFX4_4/Y gnd CLKBUF1_51/Y vdd CLKBUF1
XCLKBUF1_62 BUFX4_2/Y gnd CLKBUF1_62/Y vdd CLKBUF1
XFILL_41_0_1 gnd vdd FILL
XINVX1_114 INVX1_114/A gnd INVX1_114/Y vdd INVX1
XINVX1_103 INVX1_103/A gnd INVX1_103/Y vdd INVX1
XINVX1_125 INVX1_125/A gnd INVX1_125/Y vdd INVX1
XINVX1_147 BUFX2_85/A gnd INVX1_147/Y vdd INVX1
XINVX1_158 instruction_memory_interface_data[2] gnd INVX1_158/Y vdd INVX1
XINVX1_136 INVX1_495/A gnd INVX1_136/Y vdd INVX1
XINVX1_169 instruction_memory_interface_data[13] gnd INVX1_169/Y vdd INVX1
XFILL_32_0_1 gnd vdd FILL
XAOI21X1_107 INVX1_393/A NOR2X1_269/Y BUFX4_86/Y gnd OAI21X1_541/C vdd AOI21X1
XAOI21X1_118 BUFX4_52/Y AOI21X1_118/B AOI21X1_118/C gnd AOI21X1_118/Y vdd AOI21X1
XAOI21X1_129 AOI22X1_99/Y OAI21X1_588/Y OAI21X1_589/Y gnd AOI21X1_129/Y vdd AOI21X1
XINVX1_681 INVX1_681/A gnd INVX1_681/Y vdd INVX1
XINVX1_670 INVX1_460/A gnd INVX1_670/Y vdd INVX1
XINVX1_692 OR2X2_58/B gnd INVX1_692/Y vdd INVX1
XFILL_23_0_1 gnd vdd FILL
XINVX4_11 INVX4_11/A gnd INVX4_11/Y vdd INVX4
XFILL_6_1_1 gnd vdd FILL
XFILL_14_0_1 gnd vdd FILL
XBUFX4_220 BUFX4_222/A gnd BUFX4_220/Y vdd BUFX4
XBUFX4_231 BUFX4_233/A gnd BUFX4_231/Y vdd BUFX4
XBUFX4_264 BUFX4_264/A gnd BUFX4_264/Y vdd BUFX4
XBUFX4_242 BUFX4_242/A gnd INVX4_1/A vdd BUFX4
XBUFX4_253 BUFX4_253/A gnd BUFX4_253/Y vdd BUFX4
XNOR2X1_313 BUFX4_87/Y AND2X2_48/Y gnd NOR2X1_313/Y vdd NOR2X1
XBUFX4_275 BUFX4_276/A gnd BUFX4_275/Y vdd BUFX4
XNOR2X1_302 NOR2X1_253/A NOR2X1_302/B gnd NOR2X1_302/Y vdd NOR2X1
XNOR2X1_324 INVX1_409/Y INVX4_10/A gnd NOR2X1_324/Y vdd NOR2X1
XNOR2X1_357 INVX2_22/Y NOR2X1_357/B gnd NOR2X1_357/Y vdd NOR2X1
XNOR2X1_368 BUFX4_127/Y NOR2X1_368/B gnd NOR2X1_368/Y vdd NOR2X1
XNOR2X1_335 NOR2X1_333/Y AND2X2_58/Y gnd NOR2X1_335/Y vdd NOR2X1
XNOR2X1_346 NOR2X1_73/Y INVX8_12/Y gnd NOR2X1_347/A vdd NOR2X1
XFILL_32_2 gnd vdd FILL
XNOR2X1_379 NOR2X1_71/A NOR2X1_71/B gnd NOR2X1_379/Y vdd NOR2X1
XFILL_25_1 gnd vdd FILL
XOAI21X1_819 NOR2X1_381/Y NAND2X1_643/Y OAI21X1_819/C gnd OAI21X1_819/Y vdd OAI21X1
XOAI21X1_808 BUFX4_178/Y INVX1_461/Y NAND2X1_631/Y gnd OAI21X1_808/Y vdd OAI21X1
XNAND2X1_803 INVX1_565/Y BUFX4_204/Y gnd NAND3X1_253/C vdd NAND2X1
XNAND2X1_814 OR2X2_49/A BUFX2_91/A gnd NAND2X1_814/Y vdd NAND2X1
XNAND2X1_825 OAI21X1_67/Y BUFX4_60/Y gnd NAND2X1_825/Y vdd NAND2X1
XNAND2X1_836 NAND2X1_834/Y NAND2X1_836/B gnd NAND2X1_38/B vdd NAND2X1
XNAND2X1_858 OAI21X1_78/Y BUFX4_61/Y gnd NAND2X1_858/Y vdd NAND2X1
XNAND2X1_869 NAND2X1_867/Y NAND2X1_869/B gnd NAND2X1_49/B vdd NAND2X1
XNAND2X1_847 INVX1_594/Y BUFX4_94/Y gnd NAND3X1_279/C vdd NAND2X1
XNAND3X1_20 NAND3X1_20/A BUFX4_110/Y BUFX4_138/Y gnd NAND3X1_21/B vdd NAND3X1
XNAND3X1_31 BUFX4_75/Y NAND3X1_30/Y NAND3X1_31/C gnd NAND3X1_31/Y vdd NAND3X1
XNAND3X1_42 NAND3X1_42/A INVX8_2/A BUFX4_137/Y gnd NAND3X1_43/B vdd NAND3X1
XNAND3X1_53 BUFX4_73/Y NAND3X1_53/B NAND3X1_53/C gnd NAND3X1_53/Y vdd NAND3X1
XNAND3X1_64 NAND3X1_64/A BUFX4_114/Y BUFX4_136/Y gnd NAND3X1_64/Y vdd NAND3X1
XNAND3X1_75 NOR2X1_6/A OR2X2_1/B INVX1_231/Y gnd AOI21X1_4/C vdd NAND3X1
XNAND3X1_97 INVX2_31/Y INVX2_32/Y NAND3X1_97/C gnd OR2X2_20/B vdd NAND3X1
XNAND3X1_86 AND2X2_16/B NAND3X1_85/A AND2X2_16/A gnd AOI21X1_33/C vdd NAND3X1
XNOR2X1_20 OR2X2_6/B NOR2X1_20/B gnd NOR2X1_20/Y vdd NOR2X1
XNOR2X1_31 INVX2_9/Y NOR2X1_31/B gnd NOR2X1_31/Y vdd NOR2X1
XNOR2X1_42 NOR2X1_42/A NOR2X1_42/B gnd NOR2X1_42/Y vdd NOR2X1
XNOR2X1_64 NOR2X1_64/A INVX1_294/Y gnd NOR2X1_64/Y vdd NOR2X1
XNOR2X1_53 INVX1_279/Y NOR2X1_53/B gnd INVX1_280/A vdd NOR2X1
XNOR2X1_97 INVX2_36/Y INVX2_53/A gnd NOR2X1_97/Y vdd NOR2X1
XNOR2X1_75 INVX1_303/Y INVX4_2/Y gnd NOR2X1_75/Y vdd NOR2X1
XNOR2X1_86 INVX2_23/A INVX2_24/A gnd NOR2X1_86/Y vdd NOR2X1
XNAND2X1_8 BUFX4_17/Y NAND2X1_8/B gnd OAI21X1_8/C vdd NAND2X1
XNOR2X1_110 INVX8_3/A MUX2X1_11/Y gnd NOR2X1_110/Y vdd NOR2X1
XNOR2X1_121 INVX2_42/A MUX2X1_35/A gnd OAI22X1_9/A vdd NOR2X1
XNOR2X1_132 INVX2_51/A NOR2X1_132/B gnd AND2X2_42/A vdd NOR2X1
XNOR2X1_143 NOR2X1_143/A OR2X2_15/Y gnd NAND3X1_94/C vdd NOR2X1
XNOR2X1_176 OR2X2_23/B NOR2X1_176/B gnd NOR2X1_176/Y vdd NOR2X1
XNOR2X1_165 NOR2X1_165/A OR2X2_20/Y gnd NOR2X1_165/Y vdd NOR2X1
XNOR2X1_154 INVX2_51/Y INVX1_358/A gnd INVX1_377/A vdd NOR2X1
XNOR2X1_198 BUFX4_126/Y INVX4_5/A gnd AOI22X1_87/A vdd NOR2X1
XNOR2X1_187 INVX8_5/A MUX2X1_25/A gnd NOR2X1_187/Y vdd NOR2X1
XOAI21X1_605 INVX2_67/Y OAI21X1_605/B NOR2X1_307/Y gnd OAI21X1_605/Y vdd OAI21X1
XOAI21X1_638 AND2X2_50/Y AOI21X1_68/B AOI21X1_153/Y gnd OR2X2_37/A vdd OAI21X1
XOAI21X1_616 INVX1_370/Y BUFX4_126/Y NOR2X1_186/Y gnd OR2X2_36/A vdd OAI21X1
XOAI21X1_627 NAND2X1_399/Y OR2X2_40/A AOI21X1_151/Y gnd NOR3X1_58/A vdd OAI21X1
XOAI21X1_649 NAND2X1_564/B INVX8_5/A NAND2X1_550/Y gnd NAND2X1_572/B vdd OAI21X1
XNAND2X1_611 INVX1_243/A BUFX4_264/Y gnd NAND2X1_611/Y vdd NAND2X1
XNAND2X1_600 INVX1_429/Y OAI21X1_744/B gnd AOI21X1_208/B vdd NAND2X1
XNAND2X1_644 BUFX4_245/Y XNOR2X1_12/Y gnd OAI21X1_819/C vdd NAND2X1
XNAND2X1_655 OR2X2_45/B XNOR2X1_22/Y gnd OAI21X1_829/C vdd NAND2X1
XINVX1_23 gnd gnd INVX1_23/Y vdd INVX1
XNAND2X1_622 INVX2_14/A BUFX4_265/Y gnd NAND2X1_622/Y vdd NAND2X1
XNAND2X1_633 INVX1_285/A BUFX4_266/Y gnd NAND2X1_633/Y vdd NAND2X1
XINVX1_12 gnd gnd INVX1_12/Y vdd INVX1
XNAND2X1_666 OR2X2_45/B XNOR2X1_36/Y gnd OAI21X1_840/C vdd NAND2X1
XNAND2X1_677 INVX8_13/A XNOR2X1_41/Y gnd OAI21X1_852/C vdd NAND2X1
XNAND2X1_688 BUFX4_241/Y XOR2X1_7/Y gnd OAI21X1_861/C vdd NAND2X1
XINVX1_45 gnd gnd INVX1_45/Y vdd INVX1
XINVX1_34 gnd gnd INVX1_34/Y vdd INVX1
XINVX1_67 INVX1_67/A gnd INVX1_67/Y vdd INVX1
XINVX1_56 gnd gnd INVX1_56/Y vdd INVX1
XINVX1_78 INVX1_78/A gnd INVX1_78/Y vdd INVX1
XINVX1_89 INVX1_89/A gnd INVX1_89/Y vdd INVX1
XNAND2X1_699 INVX1_495/A INVX1_496/Y gnd NAND3X1_186/C vdd NAND2X1
XDFFPOSX1_8 AOI22X1_8/D CLKBUF1_18/Y DFFPOSX1_8/D gnd vdd DFFPOSX1
XFILL_40_6_0 gnd vdd FILL
XFILL_31_6_0 gnd vdd FILL
XNAND3X1_250 INVX1_564/Y BUFX4_206/Y BUFX4_33/Y gnd NAND3X1_250/Y vdd NAND3X1
XNAND3X1_261 BUFX4_121/Y NAND3X1_260/Y NAND3X1_261/C gnd NAND2X1_821/B vdd NAND3X1
XNAND3X1_283 BUFX4_119/Y NAND3X1_283/B NAND3X1_283/C gnd NAND2X1_854/B vdd NAND3X1
XNAND3X1_272 INVX1_589/Y BUFX4_101/Y BUFX4_166/Y gnd NAND3X1_272/Y vdd NAND3X1
XNAND3X1_294 INVX1_611/Y BUFX4_102/Y BUFX4_168/Y gnd NAND3X1_294/Y vdd NAND3X1
XFILL_39_7_0 gnd vdd FILL
XOAI22X1_18 OAI22X1_43/B INVX2_57/Y AOI21X1_87/Y BUFX4_275/Y gnd OAI22X1_18/Y vdd
+ OAI22X1
XOAI22X1_29 OAI22X1_29/A OAI22X1_43/B INVX8_12/Y OAI22X1_8/D gnd OAI22X1_29/Y vdd
+ OAI22X1
XFILL_22_6_0 gnd vdd FILL
XOAI21X1_402 INVX2_53/Y BUFX4_43/Y OAI21X1_583/C gnd MUX2X1_23/A vdd OAI21X1
XOAI21X1_413 BUFX4_58/Y MUX2X1_20/Y NAND2X1_398/Y gnd NOR2X1_207/B vdd OAI21X1
XOAI21X1_446 AOI21X1_63/Y AOI21X1_62/Y AOI22X1_81/D gnd NOR2X1_214/A vdd OAI21X1
XOAI21X1_435 INVX8_3/A MUX2X1_22/Y AOI21X1_67/Y gnd OAI21X1_435/Y vdd OAI21X1
XOAI21X1_457 OAI21X1_457/A INVX2_54/Y OAI21X1_457/C gnd OAI21X1_458/A vdd OAI21X1
XOAI21X1_424 AND2X2_30/Y OAI21X1_424/B OAI21X1_424/C gnd NOR2X1_210/B vdd OAI21X1
XOAI21X1_468 INVX2_47/Y AOI21X1_81/B AOI21X1_81/Y gnd OAI21X1_468/Y vdd OAI21X1
XOAI21X1_479 AOI21X1_88/C OAI22X1_17/B AOI21X1_81/B gnd AOI21X1_87/B vdd OAI21X1
XDFFPOSX1_360 INVX1_327/A CLKBUF1_4/Y OAI21X1_17/Y gnd vdd DFFPOSX1
XDFFPOSX1_371 OR2X2_54/A CLKBUF1_57/Y OAI21X1_28/Y gnd vdd DFFPOSX1
XDFFPOSX1_382 INVX1_442/A CLKBUF1_38/Y OAI21X1_39/Y gnd vdd DFFPOSX1
XDFFPOSX1_393 INVX2_83/A CLKBUF1_37/Y OAI21X1_50/Y gnd vdd DFFPOSX1
XNAND2X1_441 AOI22X1_87/A INVX1_379/Y gnd NAND3X1_114/C vdd NAND2X1
XNAND2X1_430 BUFX4_223/Y NAND2X1_430/B gnd NAND2X1_430/Y vdd NAND2X1
XNAND2X1_463 NOR2X1_229/Y NOR2X1_194/Y gnd OAI21X1_489/C vdd NAND2X1
XNAND2X1_452 MUX2X1_20/S AND2X2_28/Y gnd MUX2X1_29/B vdd NAND2X1
XFILL_5_7_0 gnd vdd FILL
XNAND2X1_485 INVX2_45/Y NOR2X1_125/B gnd OAI21X1_526/B vdd NAND2X1
XNAND2X1_496 INVX8_5/A NAND2X1_496/B gnd NAND2X1_496/Y vdd NAND2X1
XNAND2X1_474 AOI22X1_88/Y AOI21X1_96/A gnd NAND2X1_474/Y vdd NAND2X1
XFILL_13_6_0 gnd vdd FILL
XOAI21X1_980 NOR2X1_481/Y INVX4_12/A data_memory_interface_data[16] gnd OAI21X1_980/Y
+ vdd OAI21X1
XOAI21X1_991 INVX4_13/Y INVX8_16/Y data_memory_interface_data[27] gnd OAI21X1_991/Y
+ vdd OAI21X1
XOAI21X1_62 INVX1_62/Y BUFX4_29/Y OAI21X1_62/C gnd OAI21X1_62/Y vdd OAI21X1
XOAI21X1_51 INVX1_51/Y BUFX4_31/Y NAND2X1_51/Y gnd OAI21X1_51/Y vdd OAI21X1
XOAI21X1_40 INVX1_40/Y BUFX4_27/Y NAND2X1_40/Y gnd OAI21X1_40/Y vdd OAI21X1
XOAI21X1_95 INVX1_96/Y BUFX4_162/Y NAND2X1_97/Y gnd OAI21X1_95/Y vdd OAI21X1
XOAI21X1_73 INVX1_74/Y BUFX4_162/Y NAND2X1_75/Y gnd OAI21X1_73/Y vdd OAI21X1
XOAI21X1_84 INVX1_85/Y BUFX4_158/Y NAND2X1_86/Y gnd OAI21X1_84/Y vdd OAI21X1
XAOI22X1_109 INVX1_433/Y INVX8_12/A OR2X2_24/Y INVX2_26/A gnd AOI22X1_109/Y vdd AOI22X1
XOAI21X1_210 BUFX4_142/Y INVX1_208/Y AOI22X1_25/Y gnd OAI21X1_210/Y vdd OAI21X1
XOAI21X1_221 OR2X2_4/A INVX1_219/Y AOI22X1_36/Y gnd OAI21X1_221/Y vdd OAI21X1
XOAI21X1_254 NOR2X1_35/B AOI21X1_26/C AOI21X1_29/A gnd XNOR2X1_36/A vdd OAI21X1
XOAI21X1_243 INVX2_8/Y AOI22X1_47/Y OAI21X1_242/Y gnd XNOR2X1_19/A vdd OAI21X1
XOAI21X1_265 NOR2X1_45/B OR2X2_12/Y OR2X2_13/Y gnd AOI21X1_28/C vdd OAI21X1
XOAI21X1_232 AOI21X1_8/Y NOR3X1_49/Y INVX1_234/A gnd OAI21X1_232/Y vdd OAI21X1
XOAI21X1_298 INVX1_324/Y INVX4_4/A NAND2X1_223/Y gnd MUX2X1_42/B vdd OAI21X1
XOAI21X1_276 AOI21X1_26/Y OAI21X1_276/B AND2X2_18/Y gnd AOI21X1_34/B vdd OAI21X1
XINVX1_307 INVX1_307/A gnd NOR2X1_78/A vdd INVX1
XOAI21X1_287 INVX1_310/Y INVX4_4/A NAND2X1_203/Y gnd INVX2_24/A vdd OAI21X1
XAND2X2_32 AND2X2_32/A BUFX4_216/Y gnd MUX2X1_34/B vdd AND2X2
XINVX1_329 INVX1_329/A gnd INVX1_329/Y vdd INVX1
XINVX1_318 INVX2_82/A gnd INVX1_318/Y vdd INVX1
XAND2X2_10 INVX1_66/A NOR2X1_1/A gnd AND2X2_10/Y vdd AND2X2
XAND2X2_21 AND2X2_21/A INVX2_26/A gnd AND2X2_21/Y vdd AND2X2
XAND2X2_54 AND2X2_54/A INVX4_10/Y gnd AND2X2_54/Y vdd AND2X2
XAND2X2_43 AND2X2_43/A BUFX4_78/Y gnd AND2X2_43/Y vdd AND2X2
XAND2X2_65 AND2X2_64/B AND2X2_65/B gnd AND2X2_65/Y vdd AND2X2
XAND2X2_76 BUFX2_43/A BUFX2_44/A gnd AND2X2_76/Y vdd AND2X2
XAND2X2_87 AND2X2_87/A AND2X2_87/B gnd AND2X2_87/Y vdd AND2X2
XDFFPOSX1_190 BUFX2_77/A CLKBUF1_16/Y INVX1_435/A gnd vdd DFFPOSX1
XAND2X2_98 NAND3X1_1/B NOR2X1_3/A gnd AND2X2_98/Y vdd AND2X2
XNAND2X1_260 INVX2_44/Y MUX2X1_9/Y gnd AOI22X1_72/B vdd NAND2X1
XNAND2X1_271 INVX8_5/A MUX2X1_14/Y gnd AOI21X1_63/A vdd NAND2X1
XNAND2X1_282 INVX2_46/Y MUX2X1_16/Y gnd AOI22X1_85/B vdd NAND2X1
XNAND2X1_293 INVX1_342/Y MUX2X1_31/B gnd AOI22X1_89/A vdd NAND2X1
XFILL_36_5_0 gnd vdd FILL
XCLKBUF1_41 BUFX4_3/Y gnd CLKBUF1_41/Y vdd CLKBUF1
XCLKBUF1_30 BUFX4_4/Y gnd CLKBUF1_30/Y vdd CLKBUF1
XCLKBUF1_52 BUFX4_5/Y gnd CLKBUF1_52/Y vdd CLKBUF1
XCLKBUF1_63 BUFX4_7/Y gnd CLKBUF1_63/Y vdd CLKBUF1
XFILL_2_5_0 gnd vdd FILL
XFILL_27_5_0 gnd vdd FILL
XFILL_10_4_0 gnd vdd FILL
XINVX1_104 INVX1_104/A gnd INVX1_104/Y vdd INVX1
XINVX1_115 INVX1_115/A gnd INVX1_115/Y vdd INVX1
XINVX1_148 BUFX2_86/A gnd INVX1_148/Y vdd INVX1
XINVX1_159 instruction_memory_interface_data[3] gnd INVX1_159/Y vdd INVX1
XINVX1_126 INVX1_126/A gnd INVX1_126/Y vdd INVX1
XINVX1_137 OR2X2_49/B gnd AOI22X1_6/D vdd INVX1
XFILL_18_5_0 gnd vdd FILL
XAOI21X1_108 INVX8_8/A NOR2X1_123/B NOR2X1_191/Y gnd MUX2X1_36/B vdd AOI21X1
XAOI21X1_119 OAI22X1_8/C BUFX4_153/Y OAI22X1_29/Y gnd AOI21X1_119/Y vdd AOI21X1
XINVX1_671 INVX1_458/A gnd INVX1_671/Y vdd INVX1
XINVX1_660 INVX2_74/A gnd INVX1_660/Y vdd INVX1
XINVX1_693 OR2X2_59/A gnd INVX1_693/Y vdd INVX1
XINVX1_682 INVX1_444/A gnd INVX1_682/Y vdd INVX1
XINVX4_12 INVX4_12/A gnd INVX4_12/Y vdd INVX4
XFILL_42_3_0 gnd vdd FILL
XBUFX4_210 BUFX4_210/A gnd BUFX4_210/Y vdd BUFX4
XBUFX4_221 BUFX4_222/A gnd BUFX4_221/Y vdd BUFX4
XBUFX4_243 BUFX4_242/A gnd OR2X2_45/B vdd BUFX4
XBUFX4_254 BUFX4_253/A gnd BUFX4_254/Y vdd BUFX4
XBUFX4_232 BUFX4_233/A gnd BUFX4_232/Y vdd BUFX4
XNOR2X1_303 INVX2_39/Y MUX2X1_37/B gnd NOR2X1_303/Y vdd NOR2X1
XNOR2X1_325 NOR2X1_325/A NOR2X1_325/B gnd NOR2X1_326/B vdd NOR2X1
XNOR2X1_314 INVX8_3/A NOR2X1_314/B gnd NOR2X1_314/Y vdd NOR2X1
XBUFX4_276 BUFX4_276/A gnd BUFX4_276/Y vdd BUFX4
XBUFX4_265 BUFX4_264/A gnd BUFX4_265/Y vdd BUFX4
XNOR2X1_336 NOR2X1_336/A NOR2X1_336/B gnd NOR2X1_336/Y vdd NOR2X1
XNOR2X1_347 NOR2X1_347/A NOR2X1_347/B gnd NOR2X1_347/Y vdd NOR2X1
XNOR2X1_358 BUFX4_276/Y NOR2X1_357/Y gnd NOR2X1_358/Y vdd NOR2X1
XNOR2X1_369 NOR2X1_369/A OR2X2_42/A gnd NOR3X1_64/A vdd NOR2X1
XFILL_33_3_0 gnd vdd FILL
XFILL_18_1 gnd vdd FILL
XOAI21X1_809 BUFX4_178/Y INVX1_462/Y NAND2X1_632/Y gnd OAI21X1_809/Y vdd OAI21X1
XNAND2X1_804 NAND2X1_802/Y NAND2X1_804/B gnd NAND2X1_32/B vdd NAND2X1
XNAND2X1_815 OR2X2_50/A OR2X2_52/B gnd AOI22X1_112/C vdd NAND2X1
XINVX1_490 INVX1_490/A gnd INVX1_490/Y vdd INVX1
XNAND2X1_837 OAI21X1_71/Y BUFX4_61/Y gnd NAND2X1_837/Y vdd NAND2X1
XNAND2X1_826 INVX1_580/Y BUFX4_95/Y gnd NAND3X1_265/C vdd NAND2X1
XNAND2X1_859 INVX1_602/Y BUFX4_94/Y gnd NAND3X1_287/C vdd NAND2X1
XNAND2X1_848 NAND2X1_846/Y NAND2X1_848/B gnd NAND2X1_42/B vdd NAND2X1
XFILL_24_3_0 gnd vdd FILL
XNAND3X1_10 NAND3X1_10/A INVX8_2/A BUFX4_137/Y gnd NAND3X1_11/B vdd NAND3X1
XFILL_7_4_0 gnd vdd FILL
XNAND3X1_21 BUFX4_75/Y NAND3X1_21/B NAND3X1_21/C gnd NAND3X1_21/Y vdd NAND3X1
XNAND3X1_32 NAND3X1_32/A BUFX4_111/Y BUFX4_139/Y gnd NAND3X1_32/Y vdd NAND3X1
XNAND3X1_43 BUFX4_72/Y NAND3X1_43/B NAND3X1_43/C gnd NAND3X1_43/Y vdd NAND3X1
XNAND3X1_54 NAND3X1_54/A BUFX4_114/Y BUFX4_136/Y gnd NAND3X1_55/B vdd NAND3X1
XNAND3X1_65 BUFX4_76/Y NAND3X1_64/Y NAND3X1_65/C gnd NAND3X1_65/Y vdd NAND3X1
XNAND3X1_98 NOR2X1_166/Y NAND3X1_98/B NAND3X1_98/C gnd NOR2X1_171/A vdd NAND3X1
XNAND3X1_76 INVX1_66/A INVX1_232/Y AND2X2_9/Y gnd NAND3X1_76/Y vdd NAND3X1
XNAND3X1_87 INVX1_297/Y INVX1_300/A NAND3X1_87/C gnd NAND3X1_87/Y vdd NAND3X1
XNOR2X1_21 INVX1_228/A OR2X2_5/B gnd NOR2X1_21/Y vdd NOR2X1
XNOR2X1_10 NOR2X1_8/A NOR2X1_10/B gnd AND2X2_7/B vdd NOR2X1
XNOR2X1_43 XOR2X1_3/B NOR2X1_43/B gnd NOR2X1_43/Y vdd NOR2X1
XNOR2X1_32 INVX2_10/Y NOR2X1_32/B gnd NOR2X1_32/Y vdd NOR2X1
XNOR2X1_54 XOR2X1_6/B NOR2X1_54/B gnd INVX1_282/A vdd NOR2X1
XNOR2X1_65 INVX1_296/Y NOR2X1_65/B gnd INVX1_297/A vdd NOR2X1
XNOR2X1_76 NOR2X1_76/A INVX4_2/A gnd NOR2X1_76/Y vdd NOR2X1
XNOR2X1_87 INVX2_23/Y INVX2_24/Y gnd NOR2X1_87/Y vdd NOR2X1
XNOR2X1_98 INVX2_37/Y MUX2X1_42/A gnd NOR2X1_98/Y vdd NOR2X1
XFILL_15_3_0 gnd vdd FILL
XNAND2X1_9 BUFX4_17/Y NAND2X1_9/B gnd OAI21X1_9/C vdd NAND2X1
XNOR2X1_100 INVX2_29/Y INVX2_30/A gnd AOI21X1_38/A vdd NOR2X1
XNOR2X1_122 INVX2_43/Y MUX2X1_8/Y gnd OAI22X1_9/C vdd NOR2X1
XNOR2X1_111 INVX2_38/Y MUX2X1_3/Y gnd OAI22X1_7/B vdd NOR2X1
XMUX2X1_50 MUX2X1_50/A MUX2X1_50/B INVX8_3/A gnd MUX2X1_50/Y vdd MUX2X1
XNOR2X1_133 NOR2X1_133/A OR2X2_17/Y gnd INVX1_355/A vdd NOR2X1
XNOR2X1_144 INVX1_342/Y MUX2X1_15/Y gnd AOI22X1_86/A vdd NOR2X1
XNOR2X1_166 INVX1_342/A INVX2_46/A gnd NOR2X1_166/Y vdd NOR2X1
XNOR2X1_155 INVX2_51/Y NOR2X1_132/B gnd AOI21X1_49/B vdd NOR2X1
XNOR2X1_188 INVX8_3/A NOR2X1_188/B gnd NOR2X1_188/Y vdd NOR2X1
XNOR2X1_199 INVX8_7/A INVX4_5/A gnd INVX4_7/A vdd NOR2X1
XNOR2X1_177 NOR2X1_1/A INVX1_346/Y gnd NOR2X1_177/Y vdd NOR2X1
XOAI21X1_606 OAI22X1_31/C NAND2X1_500/B OAI21X1_606/C gnd OAI21X1_606/Y vdd OAI21X1
XOAI21X1_639 AND2X2_48/Y NOR2X1_319/Y AOI21X1_37/B gnd OAI21X1_639/Y vdd OAI21X1
XOAI21X1_628 NOR2X1_316/B INVX2_68/Y INVX1_403/Y gnd NAND3X1_146/C vdd OAI21X1
XOAI21X1_617 NOR2X1_312/Y INVX8_12/Y AOI22X1_101/Y gnd OAI21X1_617/Y vdd OAI21X1
XNAND2X1_601 BUFX4_55/Y AND2X2_71/A gnd OAI21X1_769/C vdd NAND2X1
XNAND2X1_612 INVX1_245/A BUFX4_265/Y gnd OAI21X1_789/C vdd NAND2X1
XNAND2X1_645 OR2X2_45/A AND2X2_76/Y gnd INVX1_470/A vdd NAND2X1
XINVX1_24 gnd gnd INVX1_24/Y vdd INVX1
XNAND2X1_623 INVX1_261/A BUFX4_265/Y gnd NAND2X1_623/Y vdd NAND2X1
XINVX1_13 gnd gnd INVX1_13/Y vdd INVX1
XNAND2X1_634 INVX1_288/A BUFX4_266/Y gnd NAND2X1_634/Y vdd NAND2X1
XNAND2X1_667 BUFX2_55/A BUFX2_56/A gnd INVX1_480/A vdd NAND2X1
XNAND2X1_656 BUFX2_49/A BUFX2_50/A gnd OR2X2_46/B vdd NAND2X1
XNAND2X1_678 BUFX4_241/Y XOR2X1_5/Y gnd OAI21X1_854/C vdd NAND2X1
XINVX1_35 gnd gnd INVX1_35/Y vdd INVX1
XINVX1_46 gnd gnd INVX1_46/Y vdd INVX1
XINVX1_57 gnd gnd INVX1_57/Y vdd INVX1
XNAND2X1_689 INVX1_486/Y NOR2X1_395/B gnd NAND2X1_689/Y vdd NAND2X1
XINVX1_79 INVX1_79/A gnd INVX1_79/Y vdd INVX1
XINVX1_68 INVX1_68/A gnd INVX1_68/Y vdd INVX1
XDFFPOSX1_9 AOI22X1_9/D CLKBUF1_31/Y DFFPOSX1_9/D gnd vdd DFFPOSX1
XFILL_40_6_1 gnd vdd FILL
XFILL_31_6_1 gnd vdd FILL
XNAND3X1_240 INVX1_554/Y BUFX4_206/Y BUFX4_33/Y gnd NAND3X1_240/Y vdd NAND3X1
XNAND3X1_251 BUFX4_220/Y NAND3X1_250/Y NAND3X1_251/C gnd NAND2X1_801/B vdd NAND3X1
XNAND3X1_262 INVX1_579/Y BUFX4_103/Y BUFX4_164/Y gnd NAND3X1_262/Y vdd NAND3X1
XFILL_30_1_0 gnd vdd FILL
XNAND3X1_284 INVX1_601/Y BUFX4_101/Y BUFX4_166/Y gnd NAND3X1_284/Y vdd NAND3X1
XNAND3X1_273 BUFX4_119/Y NAND3X1_272/Y NAND3X1_273/C gnd NAND2X1_839/B vdd NAND3X1
XNAND3X1_295 BUFX4_120/Y NAND3X1_294/Y NAND2X1_871/Y gnd NAND2X1_872/B vdd NAND3X1
XFILL_39_7_1 gnd vdd FILL
XFILL_38_2_0 gnd vdd FILL
XOAI22X1_19 INVX2_54/Y OAI22X1_19/B OAI22X1_19/C NOR2X1_225/Y gnd OAI22X1_19/Y vdd
+ OAI22X1
XFILL_22_6_1 gnd vdd FILL
XOAI21X1_403 BUFX4_43/Y MUX2X1_4/Y OAI21X1_403/C gnd INVX1_368/A vdd OAI21X1
XOAI21X1_414 INVX1_354/Y BUFX4_227/Y NAND2X1_400/Y gnd NAND2X1_455/B vdd OAI21X1
XFILL_21_1_0 gnd vdd FILL
XOAI21X1_447 AOI21X1_69/Y AOI21X1_48/Y AOI22X1_73/D gnd INVX1_373/A vdd OAI21X1
XOAI21X1_425 AOI21X1_62/Y AOI21X1_78/B NOR2X1_210/B gnd AOI22X1_78/B vdd OAI21X1
XOAI21X1_436 INVX1_363/Y INVX8_5/A OAI21X1_436/C gnd MUX2X1_32/B vdd OAI21X1
XOAI21X1_469 BUFX4_41/Y AND2X2_34/A OAI21X1_469/C gnd OAI21X1_470/A vdd OAI21X1
XOAI21X1_458 OAI21X1_458/A AND2X2_33/Y BUFX4_80/Y gnd NAND3X1_112/A vdd OAI21X1
XDFFPOSX1_350 INVX1_690/A CLKBUF1_58/Y OAI21X1_7/Y gnd vdd DFFPOSX1
XDFFPOSX1_361 INVX1_325/A CLKBUF1_4/Y OAI21X1_18/Y gnd vdd DFFPOSX1
XDFFPOSX1_372 OR2X2_53/A CLKBUF1_57/Y OAI21X1_29/Y gnd vdd DFFPOSX1
XDFFPOSX1_383 INVX1_443/A CLKBUF1_29/Y OAI21X1_40/Y gnd vdd DFFPOSX1
XNAND2X1_420 BUFX4_228/Y INVX1_362/Y gnd NAND2X1_420/Y vdd NAND2X1
XDFFPOSX1_394 INVX1_454/A CLKBUF1_37/Y OAI21X1_51/Y gnd vdd DFFPOSX1
XNAND2X1_442 INVX8_4/A OAI21X1_390/B gnd OAI21X1_474/C vdd NAND2X1
XNAND2X1_453 BUFX4_83/Y MUX2X1_29/Y gnd OAI22X1_19/B vdd NAND2X1
XNAND2X1_431 NOR2X1_217/Y INVX1_360/Y gnd OAI21X1_457/C vdd NAND2X1
XNAND2X1_486 INVX4_8/Y AOI21X1_92/B gnd NAND3X1_123/C vdd NAND2X1
XFILL_5_7_1 gnd vdd FILL
XNAND2X1_497 BUFX4_214/Y NAND2X1_497/B gnd NAND2X1_497/Y vdd NAND2X1
XNAND2X1_464 BUFX4_229/Y MUX2X1_31/Y gnd NAND2X1_464/Y vdd NAND2X1
XNAND2X1_475 INVX2_54/A AND2X2_39/Y gnd NAND3X1_121/C vdd NAND2X1
XFILL_4_2_0 gnd vdd FILL
XFILL_29_2_0 gnd vdd FILL
XFILL_13_6_1 gnd vdd FILL
XFILL_12_1_0 gnd vdd FILL
XOAI21X1_970 INVX1_728/Y BUFX4_117/Y NAND3X1_361/C gnd OAI21X1_970/Y vdd OAI21X1
XOAI21X1_981 INVX1_735/Y OAI21X1_981/B OAI21X1_980/Y gnd OAI21X1_981/Y vdd OAI21X1
XOAI21X1_992 INVX1_741/Y OAI21X1_992/B OAI21X1_991/Y gnd AOI21X1_261/B vdd OAI21X1
XOAI21X1_30 INVX1_30/Y BUFX4_20/Y OAI21X1_30/C gnd OAI21X1_30/Y vdd OAI21X1
XOAI21X1_63 INVX1_63/Y BUFX4_30/Y OAI21X1_63/C gnd OAI21X1_63/Y vdd OAI21X1
XOAI21X1_52 INVX1_52/Y BUFX4_31/Y OAI21X1_52/C gnd OAI21X1_52/Y vdd OAI21X1
XOAI21X1_41 INVX1_41/Y BUFX4_32/Y NAND2X1_41/Y gnd OAI21X1_41/Y vdd OAI21X1
XOAI21X1_74 INVX1_75/Y BUFX4_163/Y NAND2X1_76/Y gnd OAI21X1_74/Y vdd OAI21X1
XOAI21X1_96 INVX1_97/Y BUFX4_156/Y NAND2X1_98/Y gnd OAI21X1_96/Y vdd OAI21X1
XOAI21X1_85 INVX1_86/Y BUFX4_158/Y NAND2X1_87/Y gnd OAI21X1_85/Y vdd OAI21X1
XOAI21X1_200 BUFX4_144/Y INVX1_198/Y AOI22X1_15/Y gnd OAI21X1_200/Y vdd OAI21X1
XOAI21X1_211 BUFX4_142/Y INVX1_209/Y AOI22X1_26/Y gnd OAI21X1_211/Y vdd OAI21X1
XOAI21X1_222 OR2X2_4/A INVX1_220/Y AOI22X1_37/Y gnd OAI21X1_222/Y vdd OAI21X1
XOAI21X1_255 INVX2_14/Y NOR2X1_41/B NAND2X1_153/Y gnd OAI21X1_255/Y vdd OAI21X1
XOAI21X1_244 AOI21X1_16/Y NOR3X1_53/Y INVX1_253/A gnd OAI21X1_244/Y vdd OAI21X1
XOAI21X1_233 INVX1_240/Y NOR2X1_29/A OAI21X1_232/Y gnd XNOR2X1_13/A vdd OAI21X1
XOAI21X1_299 INVX4_4/Y AOI22X1_54/A OAI21X1_299/C gnd NOR2X1_96/B vdd OAI21X1
XOAI21X1_266 XOR2X1_5/A XOR2X1_5/B OR2X2_14/Y gnd XNOR2X1_42/A vdd OAI21X1
XOAI21X1_277 AOI21X1_34/Y INVX1_293/Y NOR2X1_64/Y gnd AOI21X1_35/B vdd OAI21X1
XINVX1_308 INVX1_669/A gnd INVX1_308/Y vdd INVX1
XOAI21X1_288 NOR2X1_86/Y NOR2X1_87/Y INVX2_22/Y gnd INVX1_311/A vdd OAI21X1
XAND2X2_22 MUX2X1_13/Y INVX8_8/A gnd AND2X2_22/Y vdd AND2X2
XINVX1_319 INVX1_700/A gnd INVX1_319/Y vdd INVX1
XAND2X2_11 AND2X2_11/A INVX1_685/A gnd AND2X2_11/Y vdd AND2X2
XAND2X2_55 AND2X2_55/A INVX8_7/A gnd AND2X2_55/Y vdd AND2X2
XAND2X2_33 AND2X2_33/A INVX1_371/A gnd AND2X2_33/Y vdd AND2X2
XAND2X2_44 AND2X2_44/A BUFX4_85/Y gnd AND2X2_44/Y vdd AND2X2
XAND2X2_77 INVX2_72/A BUFX2_46/A gnd AND2X2_77/Y vdd AND2X2
XDFFPOSX1_180 BUFX2_23/A CLKBUF1_6/Y XOR2X1_5/Y gnd vdd DFFPOSX1
XAND2X2_66 AND2X2_66/A BUFX4_56/Y gnd AND2X2_66/Y vdd AND2X2
XAND2X2_88 AND2X2_88/A AND2X2_88/B gnd AND2X2_88/Y vdd AND2X2
XDFFPOSX1_191 BUFX2_78/A CLKBUF1_8/Y OR2X2_64/B gnd vdd DFFPOSX1
XAND2X2_99 INVX8_15/Y AND2X2_99/B gnd BUFX4_9/A vdd AND2X2
XNAND2X1_261 INVX4_4/A MUX2X1_10/A gnd NAND2X1_261/Y vdd NAND2X1
XNAND2X1_250 INVX2_41/Y MUX2X1_6/Y gnd AOI21X1_122/A vdd NAND2X1
XNAND2X1_283 INVX4_4/A INVX1_242/A gnd OAI21X1_322/C vdd NAND2X1
XNAND2X1_294 AOI22X1_89/B AOI22X1_89/A gnd AND2X2_35/B vdd NAND2X1
XNAND2X1_272 INVX4_4/A MUX2X1_14/A gnd NAND2X1_272/Y vdd NAND2X1
XFILL_6_1 gnd vdd FILL
XFILL_36_5_1 gnd vdd FILL
XFILL_35_0_0 gnd vdd FILL
XCLKBUF1_31 BUFX4_4/Y gnd CLKBUF1_31/Y vdd CLKBUF1
XCLKBUF1_20 BUFX4_1/Y gnd CLKBUF1_20/Y vdd CLKBUF1
XCLKBUF1_42 BUFX4_4/Y gnd CLKBUF1_42/Y vdd CLKBUF1
XCLKBUF1_53 BUFX4_7/Y gnd CLKBUF1_53/Y vdd CLKBUF1
XFILL_2_5_1 gnd vdd FILL
XFILL_27_5_1 gnd vdd FILL
XFILL_1_0_0 gnd vdd FILL
XFILL_26_0_0 gnd vdd FILL
XFILL_10_4_1 gnd vdd FILL
XINVX1_105 INVX1_105/A gnd INVX1_105/Y vdd INVX1
XINVX1_116 INVX1_116/A gnd INVX1_116/Y vdd INVX1
XINVX1_149 INVX1_149/A gnd INVX1_149/Y vdd INVX1
XINVX1_138 OR2X2_1/B gnd INVX1_138/Y vdd INVX1
XINVX1_127 INVX1_127/A gnd INVX1_127/Y vdd INVX1
XFILL_9_1_0 gnd vdd FILL
XFILL_18_5_1 gnd vdd FILL
XFILL_17_0_0 gnd vdd FILL
XAOI21X1_109 OAI22X1_9/B BUFX4_153/Y OAI22X1_26/Y gnd AOI21X1_109/Y vdd AOI21X1
XINVX1_672 INVX1_672/A gnd INVX1_672/Y vdd INVX1
XINVX1_650 BUFX2_94/A gnd INVX1_650/Y vdd INVX1
XINVX1_661 OR2X2_49/B gnd INVX1_661/Y vdd INVX1
XINVX1_683 OR2X2_64/B gnd INVX1_683/Y vdd INVX1
XINVX1_694 OR2X2_57/A gnd INVX1_694/Y vdd INVX1
XINVX4_13 INVX4_13/A gnd INVX4_13/Y vdd INVX4
XFILL_42_3_1 gnd vdd FILL
XBUFX4_200 INVX8_2/Y gnd BUFX4_200/Y vdd BUFX4
XBUFX4_211 INVX8_4/Y gnd MUX2X1_20/S vdd BUFX4
XBUFX4_233 BUFX4_233/A gnd BUFX4_233/Y vdd BUFX4
XBUFX4_244 BUFX4_242/A gnd NOR3X1_35/A vdd BUFX4
XBUFX4_255 AND2X2_6/Y gnd OR2X2_3/A vdd BUFX4
XBUFX4_222 BUFX4_222/A gnd BUFX4_222/Y vdd BUFX4
XNOR2X1_304 NOR2X1_304/A NOR2X1_304/B gnd NOR2X1_304/Y vdd NOR2X1
XNOR2X1_315 NOR2X1_315/A INVX4_9/Y gnd NOR2X1_315/Y vdd NOR2X1
XBUFX4_277 BUFX4_276/A gnd INVX8_11/A vdd BUFX4
XBUFX4_266 BUFX4_264/A gnd BUFX4_266/Y vdd BUFX4
XNOR2X1_337 INVX2_33/A OR2X2_39/Y gnd NOR2X1_337/Y vdd NOR2X1
XNOR2X1_326 NOR2X1_326/A NOR2X1_326/B gnd NOR2X1_326/Y vdd NOR2X1
XNOR2X1_359 INVX8_7/A MUX2X1_54/Y gnd NOR2X1_359/Y vdd NOR2X1
XNOR2X1_348 NOR2X1_348/A NOR2X1_348/B gnd NOR3X1_63/B vdd NOR2X1
XFILL_33_3_1 gnd vdd FILL
XINVX1_480 INVX1_480/A gnd INVX1_480/Y vdd INVX1
XNAND2X1_805 DFFPOSX1_41/Q INVX2_73/Y gnd NAND2X1_805/Y vdd NAND2X1
XINVX1_491 INVX1_491/A gnd INVX1_491/Y vdd INVX1
XNAND2X1_827 NAND2X1_825/Y NAND2X1_827/B gnd NAND2X1_35/B vdd NAND2X1
XNAND2X1_816 INVX1_573/Y BUFX4_94/Y gnd NAND3X1_261/C vdd NAND2X1
XNAND2X1_849 OAI21X1_75/Y BUFX4_61/Y gnd NAND2X1_849/Y vdd NAND2X1
XNAND2X1_838 INVX1_588/Y BUFX4_96/Y gnd NAND3X1_273/C vdd NAND2X1
XFILL_24_3_1 gnd vdd FILL
XNAND3X1_11 BUFX4_72/Y NAND3X1_11/B NAND3X1_11/C gnd NAND3X1_11/Y vdd NAND3X1
XFILL_7_4_1 gnd vdd FILL
XNAND3X1_22 NAND3X1_22/A BUFX4_110/Y BUFX4_138/Y gnd NAND3X1_23/B vdd NAND3X1
XNAND3X1_33 BUFX4_74/Y NAND3X1_32/Y NAND3X1_33/C gnd NAND3X1_33/Y vdd NAND3X1
XNAND3X1_44 NAND3X1_44/A INVX8_2/A BUFX4_137/Y gnd NAND3X1_45/B vdd NAND3X1
XNAND3X1_66 NAND3X1_66/A BUFX4_114/Y BUFX4_136/Y gnd NAND3X1_67/B vdd NAND3X1
XNAND3X1_55 BUFX4_73/Y NAND3X1_55/B NAND3X1_55/C gnd NAND3X1_55/Y vdd NAND3X1
XNOR2X1_11 NOR2X1_11/A INVX1_189/A gnd NOR2X1_11/Y vdd NOR2X1
XNAND3X1_99 INVX2_37/Y INVX2_36/Y NAND3X1_99/C gnd OR2X2_21/A vdd NAND3X1
XNAND3X1_77 NOR2X1_24/Y NOR2X1_25/Y AND2X2_9/Y gnd AOI21X1_8/A vdd NAND3X1
XNAND3X1_88 INVX2_26/Y INVX2_28/Y INVX1_311/Y gnd OR2X2_15/A vdd NAND3X1
XNOR2X1_33 NOR2X1_33/A NOR2X1_33/B gnd NOR2X1_33/Y vdd NOR2X1
XNOR2X1_44 OR2X2_11/B OR2X2_11/A gnd AND2X2_14/B vdd NOR2X1
XNOR2X1_55 INVX1_283/Y NOR2X1_55/B gnd NOR2X1_55/Y vdd NOR2X1
XNOR2X1_22 NOR2X1_22/A NOR2X1_22/B gnd NOR2X1_22/Y vdd NOR2X1
XNOR2X1_66 AND2X2_19/Y NOR2X1_66/B gnd NOR2X1_67/B vdd NOR2X1
XNOR2X1_77 INVX1_307/A INVX4_3/A gnd NOR2X1_77/Y vdd NOR2X1
XNOR2X1_88 NOR2X1_88/A INVX2_25/Y gnd INVX1_432/A vdd NOR2X1
XFILL_15_3_1 gnd vdd FILL
XNOR2X1_99 NOR2X1_99/A MUX2X1_46/B gnd NOR2X1_99/Y vdd NOR2X1
XNOR2X1_123 INVX2_43/A NOR2X1_123/B gnd OAI22X1_9/D vdd NOR2X1
XMUX2X1_40 MUX2X1_43/B MUX2X1_37/Y MUX2X1_40/S gnd MUX2X1_40/Y vdd MUX2X1
XNOR2X1_112 INVX2_38/A MUX2X1_39/A gnd OAI22X1_7/A vdd NOR2X1
XNOR2X1_101 INVX2_31/Y MUX2X1_44/B gnd NOR2X1_101/Y vdd NOR2X1
XMUX2X1_51 INVX2_60/Y MUX2X1_50/Y INVX8_7/A gnd MUX2X1_51/Y vdd MUX2X1
XNOR2X1_167 INVX2_42/A INVX2_43/A gnd NAND3X1_98/B vdd NOR2X1
XNOR2X1_156 BUFX4_41/Y MUX2X1_15/Y gnd AOI21X1_93/C vdd NOR2X1
XNOR2X1_145 INVX1_342/A MUX2X1_31/B gnd OAI22X1_11/A vdd NOR2X1
XNOR2X1_134 NOR2X1_134/A NOR2X1_134/B gnd INVX1_390/A vdd NOR2X1
XFILL_30_1 gnd vdd FILL
XNOR2X1_178 NOR2X1_178/A NOR2X1_176/Y gnd BUFX4_276/A vdd NOR2X1
XNOR2X1_189 INVX8_8/A INVX2_24/Y gnd OR2X2_25/A vdd NOR2X1
XOAI21X1_629 INVX2_35/Y MUX2X1_2/Y NAND3X1_146/C gnd OAI21X1_630/C vdd OAI21X1
XOAI21X1_607 OAI22X1_38/A AOI22X1_99/D AOI22X1_99/A gnd AOI21X1_145/C vdd OAI21X1
XOAI21X1_618 INVX1_400/Y OR2X2_36/Y AOI21X1_147/Y gnd NOR3X1_57/C vdd OAI21X1
XNAND2X1_602 INVX2_28/Y OR2X2_43/A gnd NAND2X1_602/Y vdd NAND2X1
XNAND2X1_646 BUFX4_245/Y XNOR2X1_13/Y gnd OAI21X1_821/C vdd NAND2X1
XNAND2X1_624 INVX1_264/A BUFX4_265/Y gnd OAI21X1_801/C vdd NAND2X1
XNAND2X1_613 INVX1_249/A BUFX4_265/Y gnd NAND2X1_613/Y vdd NAND2X1
XNAND2X1_635 NOR2X1_62/A BUFX4_266/Y gnd NAND2X1_635/Y vdd NAND2X1
XINVX1_14 gnd gnd INVX1_14/Y vdd INVX1
XNAND2X1_668 BUFX4_245/Y XOR2X1_3/Y gnd OAI21X1_843/C vdd NAND2X1
XNAND2X1_657 OR2X2_45/B XNOR2X1_25/Y gnd OAI21X1_832/C vdd NAND2X1
XNAND2X1_679 BUFX4_241/Y XNOR2X1_42/Y gnd OAI21X1_856/C vdd NAND2X1
XINVX1_25 gnd gnd INVX1_25/Y vdd INVX1
XINVX1_47 gnd gnd INVX1_47/Y vdd INVX1
XINVX1_58 gnd gnd INVX1_58/Y vdd INVX1
XINVX1_36 gnd gnd INVX1_36/Y vdd INVX1
XINVX1_69 INVX1_69/A gnd INVX1_69/Y vdd INVX1
XAOI21X1_270 AOI21X1_271/A AOI21X1_271/B AOI21X1_270/C gnd AOI21X1_270/Y vdd AOI21X1
XNAND3X1_230 INVX1_544/Y BUFX4_208/Y BUFX4_36/Y gnd NAND3X1_231/B vdd NAND3X1
XNAND3X1_241 BUFX4_218/Y NAND3X1_240/Y NAND3X1_241/C gnd NAND2X1_786/B vdd NAND3X1
XNAND3X1_263 BUFX4_122/Y NAND3X1_262/Y NAND3X1_263/C gnd NAND2X1_824/B vdd NAND3X1
XNAND3X1_252 INVX1_566/Y BUFX4_210/Y BUFX4_37/Y gnd NAND3X1_252/Y vdd NAND3X1
XFILL_30_1_1 gnd vdd FILL
XNAND3X1_274 INVX1_591/Y BUFX4_101/Y BUFX4_166/Y gnd NAND3X1_274/Y vdd NAND3X1
XNAND3X1_285 BUFX4_119/Y NAND3X1_284/Y NAND3X1_285/C gnd NAND2X1_857/B vdd NAND3X1
XNAND3X1_296 INVX1_613/Y BUFX4_103/Y BUFX4_164/Y gnd NAND3X1_296/Y vdd NAND3X1
XFILL_38_2_1 gnd vdd FILL
XOAI21X1_404 MUX2X1_40/S MUX2X1_23/A NAND2X1_388/Y gnd OAI21X1_474/A vdd OAI21X1
XFILL_21_1_1 gnd vdd FILL
XOAI21X1_437 BUFX4_228/Y NAND2X1_373/B NAND2X1_420/Y gnd OAI21X1_438/A vdd OAI21X1
XOAI21X1_448 AOI21X1_71/Y BUFX4_190/Y AOI21X1_97/A gnd OAI21X1_448/Y vdd OAI21X1
XOAI21X1_415 INVX8_5/A OAI21X1_350/Y NAND2X1_402/Y gnd OAI21X1_416/A vdd OAI21X1
XOAI21X1_426 NOR2X1_212/Y AND2X2_22/Y NAND2X1_273/Y gnd AOI21X1_77/B vdd OAI21X1
XOAI21X1_459 OAI22X1_10/A AOI22X1_73/D AOI22X1_73/A gnd AOI21X1_74/C vdd OAI21X1
XDFFPOSX1_340 INVX2_2/A CLKBUF1_59/Y OR2X2_8/B gnd vdd DFFPOSX1
XDFFPOSX1_351 INVX1_689/A CLKBUF1_53/Y OAI21X1_8/Y gnd vdd DFFPOSX1
XDFFPOSX1_362 MUX2X1_2/B CLKBUF1_21/Y OAI21X1_19/Y gnd vdd DFFPOSX1
XDFFPOSX1_373 INVX1_668/A CLKBUF1_57/Y OAI21X1_30/Y gnd vdd DFFPOSX1
XNAND2X1_410 BUFX4_213/Y MUX2X1_21/B gnd AOI22X1_81/D vdd NAND2X1
XDFFPOSX1_395 INVX2_86/A CLKBUF1_29/Y OAI21X1_52/Y gnd vdd DFFPOSX1
XDFFPOSX1_384 INVX1_444/A CLKBUF1_29/Y OAI21X1_41/Y gnd vdd DFFPOSX1
XNAND2X1_443 INVX8_3/A AOI21X1_118/B gnd OAI21X1_475/C vdd NAND2X1
XNAND2X1_454 BUFX4_215/Y NAND2X1_454/B gnd NAND2X1_454/Y vdd NAND2X1
XNAND2X1_432 INVX8_3/A NOR2X1_218/Y gnd OAI21X1_456/C vdd NAND2X1
XNAND2X1_421 BUFX4_40/Y INVX2_25/A gnd NOR2X1_235/B vdd NAND2X1
XNAND2X1_487 INVX2_43/Y NOR2X1_123/B gnd AOI22X1_96/D vdd NAND2X1
XNAND2X1_465 BUFX4_216/Y OAI21X1_543/B gnd NAND2X1_465/Y vdd NAND2X1
XNAND2X1_476 NOR2X1_241/B INVX1_388/A gnd NAND3X1_121/A vdd NAND2X1
XNAND2X1_498 OAI21X1_546/Y OAI21X1_545/Y gnd NAND2X1_498/Y vdd NAND2X1
XFILL_4_2_1 gnd vdd FILL
XFILL_29_2_1 gnd vdd FILL
XFILL_12_1_1 gnd vdd FILL
XOAI21X1_960 INVX8_17/Y INVX8_15/Y BUFX2_81/A gnd OAI21X1_960/Y vdd OAI21X1
XOAI21X1_993 INVX1_741/Y OAI21X1_993/B OAI21X1_993/C gnd AOI22X1_140/C vdd OAI21X1
XOAI21X1_982 OAI21X1_982/A OAI21X1_994/B OAI21X1_982/C gnd OAI21X1_982/Y vdd OAI21X1
XOAI21X1_971 INVX1_729/Y BUFX4_117/Y OAI21X1_971/C gnd OAI21X1_971/Y vdd OAI21X1
XINVX2_90 INVX2_90/A gnd INVX2_90/Y vdd INVX2
XOAI21X1_20 INVX1_20/Y BUFX4_24/Y OAI21X1_20/C gnd OAI21X1_20/Y vdd OAI21X1
XOAI21X1_31 INVX1_31/Y BUFX4_22/Y OAI21X1_31/C gnd OAI21X1_31/Y vdd OAI21X1
XOAI21X1_42 INVX1_42/Y BUFX4_32/Y OAI21X1_42/C gnd OAI21X1_42/Y vdd OAI21X1
XOAI21X1_53 INVX1_53/Y BUFX4_27/Y NAND2X1_53/Y gnd OAI21X1_53/Y vdd OAI21X1
XOAI21X1_75 INVX1_76/Y BUFX4_163/Y NAND2X1_77/Y gnd OAI21X1_75/Y vdd OAI21X1
XOAI21X1_86 INVX1_87/Y BUFX4_161/Y NAND2X1_88/Y gnd OAI21X1_86/Y vdd OAI21X1
XOAI21X1_64 INVX1_64/Y BUFX4_32/Y NAND2X1_64/Y gnd OAI21X1_64/Y vdd OAI21X1
XOAI21X1_97 BUFX4_272/Y BUFX4_195/Y OAI21X1_97/C gnd OAI21X1_98/C vdd OAI21X1
XOAI21X1_201 BUFX4_141/Y INVX1_199/Y AOI22X1_16/Y gnd OAI21X1_201/Y vdd OAI21X1
XOAI21X1_212 BUFX4_145/Y INVX1_210/Y AOI22X1_27/Y gnd OAI21X1_212/Y vdd OAI21X1
XOAI21X1_245 INVX2_8/Y AOI22X1_47/Y OAI21X1_244/Y gnd NAND2X1_142/B vdd OAI21X1
XOAI21X1_256 INVX1_261/A INVX1_260/Y OAI21X1_255/Y gnd NOR2X1_50/A vdd OAI21X1
XOAI21X1_234 AOI21X1_9/Y NOR3X1_50/Y INVX1_243/A gnd NAND2X1_130/B vdd OAI21X1
XOAI21X1_223 BUFX4_141/Y INVX1_221/Y AOI22X1_38/Y gnd OAI21X1_223/Y vdd OAI21X1
XOAI21X1_267 NOR2X1_30/B NOR2X1_30/A NOR2X1_48/Y gnd AOI21X1_29/B vdd OAI21X1
XOAI21X1_278 INVX1_289/Y NOR2X1_62/Y INVX1_292/A gnd INVX1_295/A vdd OAI21X1
XOAI21X1_289 INVX1_313/Y INVX4_4/A NAND2X1_204/Y gnd INVX2_25/A vdd OAI21X1
XAND2X2_12 AND2X2_12/A MUX2X1_13/A gnd AND2X2_12/Y vdd AND2X2
XINVX1_309 OR2X2_53/A gnd INVX1_309/Y vdd INVX1
XAND2X2_34 AND2X2_34/A INVX8_7/A gnd AND2X2_34/Y vdd AND2X2
XAND2X2_45 AND2X2_45/A BUFX4_79/Y gnd AND2X2_45/Y vdd AND2X2
XAND2X2_56 AND2X2_56/A AND2X2_56/B gnd AND2X2_56/Y vdd AND2X2
XAND2X2_23 AND2X2_23/A INVX1_356/Y gnd AND2X2_23/Y vdd AND2X2
XDFFPOSX1_170 BUFX2_13/A CLKBUF1_7/Y XNOR2X1_29/Y gnd vdd DFFPOSX1
XAND2X2_78 AND2X2_78/A AND2X2_78/B gnd AND2X2_78/Y vdd AND2X2
XAND2X2_67 AND2X2_67/A INVX8_3/A gnd AND2X2_67/Y vdd AND2X2
XDFFPOSX1_181 BUFX2_24/A CLKBUF1_35/Y XNOR2X1_42/Y gnd vdd DFFPOSX1
XAND2X2_89 OR2X2_54/A OR2X2_54/B gnd AND2X2_89/Y vdd AND2X2
XDFFPOSX1_192 BUFX2_79/A CLKBUF1_22/Y OR2X2_63/B gnd vdd DFFPOSX1
XNAND2X1_240 NOR2X1_104/Y INVX2_33/Y gnd NOR2X1_143/A vdd NAND2X1
XNAND2X1_262 INVX2_45/A NOR2X1_125/B gnd AND2X2_36/A vdd NAND2X1
XNAND2X1_251 AOI21X1_122/A OAI21X1_588/C gnd OAI22X1_29/A vdd NAND2X1
XNAND2X1_284 INVX8_6/A MUX2X1_30/A gnd OAI22X1_15/B vdd NAND2X1
XNAND2X1_295 INVX8_6/A MUX2X1_17/Y gnd AOI21X1_88/A vdd NAND2X1
XNAND2X1_273 MUX2X1_47/S MUX2X1_21/A gnd NAND2X1_273/Y vdd NAND2X1
XOAI21X1_790 BUFX4_181/Y INVX1_443/Y NAND2X1_613/Y gnd OAI21X1_790/Y vdd OAI21X1
XFILL_6_2 gnd vdd FILL
XFILL_35_0_1 gnd vdd FILL
XCLKBUF1_10 BUFX4_3/Y gnd CLKBUF1_10/Y vdd CLKBUF1
XCLKBUF1_32 BUFX4_6/Y gnd CLKBUF1_32/Y vdd CLKBUF1
XCLKBUF1_21 BUFX4_7/Y gnd CLKBUF1_21/Y vdd CLKBUF1
XCLKBUF1_54 BUFX4_3/Y gnd CLKBUF1_54/Y vdd CLKBUF1
XCLKBUF1_43 BUFX4_4/Y gnd CLKBUF1_43/Y vdd CLKBUF1
XFILL_1_0_1 gnd vdd FILL
XFILL_26_0_1 gnd vdd FILL
XINVX1_106 INVX1_106/A gnd INVX1_106/Y vdd INVX1
XINVX1_139 BUFX2_93/A gnd NOR3X1_2/B vdd INVX1
XINVX1_117 INVX1_117/A gnd INVX1_117/Y vdd INVX1
XINVX1_128 INVX1_128/A gnd INVX1_128/Y vdd INVX1
XFILL_9_1_1 gnd vdd FILL
XFILL_17_0_1 gnd vdd FILL
XINVX1_640 INVX1_640/A gnd INVX1_640/Y vdd INVX1
XINVX1_662 INVX1_662/A gnd INVX1_662/Y vdd INVX1
XINVX1_651 BUFX2_95/A gnd INVX1_651/Y vdd INVX1
XINVX1_673 INVX1_457/A gnd INVX1_673/Y vdd INVX1
XINVX1_684 INVX1_684/A gnd INVX1_684/Y vdd INVX1
XINVX1_695 INVX1_695/A gnd INVX1_695/Y vdd INVX1
XFILL_20_7_0 gnd vdd FILL
XINVX4_14 INVX4_14/A gnd INVX4_14/Y vdd INVX4
XFILL_11_7_0 gnd vdd FILL
XBUFX4_212 INVX8_4/Y gnd MUX2X1_49/S vdd BUFX4
XBUFX4_201 BUFX4_204/A gnd BUFX4_201/Y vdd BUFX4
XBUFX4_245 BUFX4_242/A gnd BUFX4_245/Y vdd BUFX4
XBUFX4_223 INVX8_5/Y gnd BUFX4_223/Y vdd BUFX4
XBUFX4_234 BUFX4_233/A gnd AND2X2_12/A vdd BUFX4
XNOR2X1_316 INVX2_68/Y NOR2X1_316/B gnd NOR2X1_316/Y vdd NOR2X1
XNOR2X1_305 INVX2_45/Y MUX2X1_10/Y gnd NOR2X1_305/Y vdd NOR2X1
XBUFX4_267 BUFX4_264/A gnd BUFX4_267/Y vdd BUFX4
XBUFX4_256 AND2X2_6/Y gnd BUFX4_256/Y vdd BUFX4
XNOR2X1_327 BUFX4_125/Y NOR2X1_327/B gnd NOR2X1_327/Y vdd NOR2X1
XNOR2X1_338 INVX4_9/Y INVX2_66/Y gnd NOR2X1_338/Y vdd NOR2X1
XNOR2X1_349 INVX1_307/A INVX4_3/Y gnd NOR2X1_349/Y vdd NOR2X1
XINVX1_470 INVX1_470/A gnd INVX1_470/Y vdd INVX1
XNAND2X1_806 DFFPOSX1_43/Q INVX2_74/Y gnd OAI21X1_871/C vdd NAND2X1
XINVX1_481 BUFX2_57/A gnd INVX1_481/Y vdd INVX1
XINVX1_492 INVX1_492/A gnd INVX1_492/Y vdd INVX1
XNAND2X1_828 OAI21X1_68/Y BUFX4_62/Y gnd NAND2X1_828/Y vdd NAND2X1
XNAND2X1_817 INVX1_501/A INVX2_76/Y gnd NAND2X1_817/Y vdd NAND2X1
XNAND2X1_839 NAND2X1_837/Y NAND2X1_839/B gnd NAND2X1_39/B vdd NAND2X1
XNAND3X1_12 NAND3X1_12/A BUFX4_111/Y BUFX4_139/Y gnd NAND3X1_13/B vdd NAND3X1
XNAND3X1_23 BUFX4_75/Y NAND3X1_23/B NAND3X1_23/C gnd NAND3X1_23/Y vdd NAND3X1
XNAND3X1_34 NAND3X1_34/A BUFX4_111/Y BUFX4_139/Y gnd NAND3X1_34/Y vdd NAND3X1
XNAND3X1_45 BUFX4_73/Y NAND3X1_45/B NAND3X1_45/C gnd NAND3X1_45/Y vdd NAND3X1
XNAND3X1_56 NAND3X1_56/A AND2X2_2/B BUFX4_136/Y gnd NAND3X1_57/B vdd NAND3X1
XNOR2X1_12 NOR2X1_13/A INVX1_191/Y gnd AND2X2_8/A vdd NOR2X1
XNAND3X1_89 INVX4_10/A NAND3X1_89/B INVX1_328/A gnd INVX2_33/A vdd NAND3X1
XNAND3X1_67 BUFX4_76/Y NAND3X1_67/B NAND3X1_67/C gnd NAND3X1_67/Y vdd NAND3X1
XNAND3X1_78 XNOR2X1_7/B AOI21X1_7/B NAND3X1_78/C gnd NAND3X1_78/Y vdd NAND3X1
XNOR2X1_34 NOR2X1_34/A NOR2X1_34/B gnd NOR2X1_34/Y vdd NOR2X1
XNOR2X1_45 NOR2X1_45/A NOR2X1_45/B gnd NOR2X1_45/Y vdd NOR2X1
XNOR2X1_23 NOR2X1_23/A OR2X2_8/Y gnd AOI21X1_3/B vdd NOR2X1
XNOR2X1_67 NOR2X1_67/A NOR2X1_67/B gnd NOR2X1_67/Y vdd NOR2X1
XNOR2X1_78 NOR2X1_78/A INVX4_3/Y gnd NOR2X1_78/Y vdd NOR2X1
XNOR2X1_56 INVX1_285/Y NOR2X1_56/B gnd INVX1_286/A vdd NOR2X1
XFILL_43_6_0 gnd vdd FILL
XNOR2X1_89 NOR2X1_89/A INVX2_25/A gnd INVX1_433/A vdd NOR2X1
XNOR2X1_124 INVX2_44/Y NOR2X1_249/B gnd NOR2X1_124/Y vdd NOR2X1
XMUX2X1_41 INVX2_53/A MUX2X1_42/A INVX8_8/A gnd MUX2X1_41/Y vdd MUX2X1
XNOR2X1_113 INVX2_39/Y MUX2X1_4/Y gnd OAI22X1_7/C vdd NOR2X1
XMUX2X1_30 MUX2X1_30/A MUX2X1_30/B INVX8_8/A gnd MUX2X1_30/Y vdd MUX2X1
XNOR2X1_102 INVX2_32/Y MUX2X1_44/A gnd NOR2X1_102/Y vdd NOR2X1
XMUX2X1_52 INVX2_60/Y MUX2X1_52/B INVX8_7/A gnd MUX2X1_52/Y vdd MUX2X1
XNOR2X1_146 INVX2_46/Y MUX2X1_16/Y gnd NOR2X1_232/A vdd NOR2X1
XNOR2X1_135 NOR2X1_135/A NOR2X1_135/B gnd INVX1_376/A vdd NOR2X1
XNOR2X1_157 BUFX4_40/Y INVX4_2/Y gnd AOI21X1_53/C vdd NOR2X1
XFILL_30_2 gnd vdd FILL
XFILL_34_6_0 gnd vdd FILL
XNOR2X1_168 INVX2_44/A INVX2_45/A gnd NAND3X1_98/C vdd NOR2X1
XNOR2X1_179 INVX1_347/Y OR2X2_22/A gnd NOR2X1_179/Y vdd NOR2X1
XFILL_23_1 gnd vdd FILL
XOAI21X1_619 NOR2X1_308/B OR2X2_39/A OAI21X1_646/A gnd AND2X2_48/A vdd OAI21X1
XOAI21X1_608 AOI21X1_113/Y NOR2X1_108/B OAI21X1_608/C gnd AOI21X1_146/C vdd OAI21X1
XDFFPOSX1_500 BUFX2_67/A CLKBUF1_47/Y NAND3X1_63/Y gnd vdd DFFPOSX1
XNAND2X1_603 INVX2_28/A OAI21X1_763/Y gnd NAND3X1_174/C vdd NAND2X1
XNAND2X1_625 INVX1_268/A BUFX4_264/Y gnd NAND2X1_625/Y vdd NAND2X1
XNAND2X1_614 INVX2_8/A BUFX4_268/Y gnd NAND2X1_614/Y vdd NAND2X1
XNAND2X1_636 INVX1_296/A BUFX4_267/Y gnd NAND2X1_636/Y vdd NAND2X1
XINVX1_15 gnd gnd INVX1_15/Y vdd INVX1
XNAND2X1_647 INVX8_13/A XNOR2X1_14/Y gnd OAI21X1_822/C vdd NAND2X1
XNAND2X1_669 INVX1_480/Y NOR3X1_65/Y gnd OAI21X1_846/A vdd NAND2X1
XNAND2X1_658 INVX8_13/Y NOR2X1_387/B gnd OAI21X1_833/B vdd NAND2X1
XINVX1_26 gnd gnd INVX1_26/Y vdd INVX1
XINVX1_37 gnd gnd INVX1_37/Y vdd INVX1
XINVX1_48 gnd gnd INVX1_48/Y vdd INVX1
XINVX1_59 gnd gnd INVX1_59/Y vdd INVX1
XFILL_0_6_0 gnd vdd FILL
XFILL_25_6_0 gnd vdd FILL
XAOI21X1_260 AOI21X1_263/A OAI21X1_988/Y OAI22X1_55/Y gnd AOI21X1_260/Y vdd AOI21X1
XAOI21X1_271 AOI21X1_271/A AOI21X1_271/B INVX1_758/Y gnd AOI21X1_271/Y vdd AOI21X1
XFILL_8_7_0 gnd vdd FILL
XFILL_16_6_0 gnd vdd FILL
XNAND3X1_231 BUFX4_221/Y NAND3X1_231/B NAND3X1_231/C gnd NAND2X1_771/B vdd NAND3X1
XNAND3X1_220 INVX1_534/Y BUFX4_206/Y BUFX4_33/Y gnd NAND3X1_221/B vdd NAND3X1
XNAND3X1_253 BUFX4_222/Y NAND3X1_252/Y NAND3X1_253/C gnd NAND2X1_804/B vdd NAND3X1
XNAND3X1_242 INVX1_556/Y BUFX4_208/Y BUFX4_36/Y gnd NAND3X1_242/Y vdd NAND3X1
XNAND3X1_264 INVX1_581/Y BUFX4_102/Y BUFX4_168/Y gnd NAND3X1_264/Y vdd NAND3X1
XNAND3X1_275 BUFX4_119/Y NAND3X1_274/Y NAND3X1_275/C gnd NAND2X1_842/B vdd NAND3X1
XNAND3X1_286 INVX1_603/Y BUFX4_100/Y BUFX4_165/Y gnd NAND3X1_287/B vdd NAND3X1
XNAND3X1_297 BUFX4_122/Y NAND3X1_296/Y NAND2X1_874/Y gnd NAND2X1_875/B vdd NAND3X1
XOAI21X1_405 INVX8_4/A MUX2X1_27/A NAND2X1_389/Y gnd NAND2X1_482/B vdd OAI21X1
XOAI21X1_438 OAI21X1_438/A INVX8_4/A OAI21X1_438/C gnd NOR2X1_271/B vdd OAI21X1
XOAI21X1_416 OAI21X1_416/A INVX8_4/A NAND2X1_401/Y gnd AND2X2_29/A vdd OAI21X1
XOAI21X1_427 AOI21X1_48/Y AOI22X1_79/D AOI21X1_77/B gnd AOI22X1_79/A vdd OAI21X1
XOAI21X1_449 AOI21X1_72/Y NAND2X1_426/Y AOI22X1_80/Y gnd AOI21X1_73/C vdd OAI21X1
XDFFPOSX1_330 INVX1_285/A CLKBUF1_1/Y OAI21X1_898/Y gnd vdd DFFPOSX1
XDFFPOSX1_363 MUX2X1_1/B CLKBUF1_53/Y OAI21X1_20/Y gnd vdd DFFPOSX1
XDFFPOSX1_352 INVX1_681/A CLKBUF1_48/Y OAI21X1_9/Y gnd vdd DFFPOSX1
XDFFPOSX1_374 INVX1_667/A CLKBUF1_48/Y OAI21X1_31/Y gnd vdd DFFPOSX1
XDFFPOSX1_341 XOR2X1_2/A CLKBUF1_59/Y OR2X2_8/A gnd vdd DFFPOSX1
XNAND2X1_411 AOI22X1_81/C AOI22X1_81/D gnd AOI21X1_64/A vdd NAND2X1
XNAND2X1_400 BUFX4_227/Y NAND2X1_400/B gnd NAND2X1_400/Y vdd NAND2X1
XDFFPOSX1_385 INVX2_84/A CLKBUF1_38/Y OAI21X1_42/Y gnd vdd DFFPOSX1
XDFFPOSX1_396 OR2X2_56/B CLKBUF1_62/Y OAI21X1_53/Y gnd vdd DFFPOSX1
XNAND2X1_422 INVX8_3/A OR2X2_41/A gnd OAI21X1_443/C vdd NAND2X1
XNAND2X1_444 NAND2X1_444/A AOI21X1_89/A gnd NAND3X1_114/A vdd NAND2X1
XNAND2X1_433 BUFX4_83/Y AOI22X1_83/A gnd OAI21X1_457/A vdd NAND2X1
XNAND2X1_477 INVX8_3/A NOR2X1_188/B gnd NAND2X1_477/Y vdd NAND2X1
XNAND2X1_488 AOI22X1_96/C AOI22X1_96/D gnd INVX2_59/A vdd NAND2X1
XNAND2X1_455 BUFX4_215/Y NAND2X1_455/B gnd NAND2X1_455/Y vdd NAND2X1
XNAND2X1_466 INVX8_3/A NOR2X1_236/Y gnd OAI21X1_497/C vdd NAND2X1
XNAND2X1_499 INVX2_40/Y MUX2X1_35/B gnd NAND2X1_500/B vdd NAND2X1
XFILL_40_4_0 gnd vdd FILL
XOAI21X1_961 INVX4_14/Y INVX1_722/Y OAI21X1_960/Y gnd OAI21X1_961/Y vdd OAI21X1
XOAI21X1_950 BUFX4_11/Y NOR2X1_470/Y INVX2_88/Y gnd BUFX4_118/A vdd OAI21X1
XOAI21X1_994 OAI21X1_994/A OAI21X1_994/B AOI22X1_140/Y gnd OAI21X1_994/Y vdd OAI21X1
XOAI21X1_972 INVX1_730/Y BUFX4_117/Y OAI21X1_972/C gnd OAI21X1_972/Y vdd OAI21X1
XOAI21X1_983 INVX4_13/Y INVX8_16/Y data_memory_interface_data[25] gnd OAI21X1_984/C
+ vdd OAI21X1
XINVX2_91 data_memory_interface_data[7] gnd INVX2_91/Y vdd INVX2
XINVX2_80 INVX2_80/A gnd INVX2_80/Y vdd INVX2
XOAI21X1_10 INVX1_10/Y BUFX4_23/Y OAI21X1_10/C gnd OAI21X1_10/Y vdd OAI21X1
XOAI21X1_21 INVX1_21/Y BUFX4_18/Y OAI21X1_21/C gnd OAI21X1_21/Y vdd OAI21X1
XOAI21X1_32 INVX1_32/Y BUFX4_20/Y OAI21X1_32/C gnd OAI21X1_32/Y vdd OAI21X1
XOAI21X1_43 INVX1_43/Y BUFX4_30/Y OAI21X1_43/C gnd OAI21X1_43/Y vdd OAI21X1
XFILL_31_4_0 gnd vdd FILL
XOAI21X1_54 INVX1_54/Y BUFX4_30/Y NAND2X1_54/Y gnd OAI21X1_54/Y vdd OAI21X1
XOAI21X1_87 INVX1_88/Y BUFX4_157/Y NAND2X1_89/Y gnd OAI21X1_87/Y vdd OAI21X1
XOAI21X1_65 INVX1_65/Y BUFX4_162/Y NAND2X1_67/Y gnd OAI21X1_65/Y vdd OAI21X1
XOAI21X1_76 INVX1_77/Y BUFX4_159/Y NAND2X1_78/Y gnd OAI21X1_76/Y vdd OAI21X1
XOAI21X1_98 BUFX4_182/Y INVX1_98/Y OAI21X1_98/C gnd INVX1_503/A vdd OAI21X1
XFILL_39_5_0 gnd vdd FILL
XFILL_22_4_0 gnd vdd FILL
XOAI21X1_202 BUFX4_141/Y INVX1_200/Y AOI22X1_17/Y gnd OAI21X1_202/Y vdd OAI21X1
XOAI21X1_213 BUFX4_142/Y INVX1_211/Y AOI22X1_28/Y gnd OAI21X1_213/Y vdd OAI21X1
XOAI21X1_224 OR2X2_4/A INVX1_222/Y AOI22X1_39/Y gnd OAI21X1_224/Y vdd OAI21X1
XOAI21X1_246 NOR2X1_35/B NOR2X1_38/B NAND2X1_142/Y gnd AOI21X1_17/B vdd OAI21X1
XOAI21X1_235 INVX1_243/Y AOI22X1_45/Y OAI21X1_232/Y gnd NAND2X1_131/B vdd OAI21X1
XOAI21X1_268 NOR2X1_50/Y INVX1_269/A AND2X2_15/Y gnd NAND3X1_85/C vdd OAI21X1
XOAI21X1_257 XNOR2X1_9/Y INVX1_233/Y INVX1_262/Y gnd OAI21X1_258/B vdd OAI21X1
XOAI21X1_279 AOI21X1_36/Y INVX1_295/A AND2X2_19/Y gnd NAND3X1_87/C vdd OAI21X1
XAND2X2_13 OR2X2_9/A INVX2_5/Y gnd AND2X2_13/Y vdd AND2X2
XAND2X2_46 AND2X2_46/A INVX2_63/Y gnd AND2X2_46/Y vdd AND2X2
XAND2X2_35 AND2X2_35/A AND2X2_35/B gnd AND2X2_35/Y vdd AND2X2
XAND2X2_24 OR2X2_44/A NOR2X1_6/A gnd AND2X2_24/Y vdd AND2X2
XDFFPOSX1_171 BUFX2_14/A CLKBUF1_26/Y XNOR2X1_30/Y gnd vdd DFFPOSX1
XAND2X2_57 NOR3X1_56/Y AND2X2_57/B gnd NOR3X1_60/B vdd AND2X2
XDFFPOSX1_182 BUFX2_25/A CLKBUF1_6/Y XOR2X1_6/Y gnd vdd DFFPOSX1
XAND2X2_68 NOR3X1_56/Y AND2X2_68/B gnd AND2X2_68/Y vdd AND2X2
XDFFPOSX1_160 BUFX2_3/A CLKBUF1_5/Y XNOR2X1_7/Y gnd vdd DFFPOSX1
XAND2X2_79 AND2X2_79/A AND2X2_79/B gnd AND2X2_79/Y vdd AND2X2
XDFFPOSX1_193 BUFX2_80/A CLKBUF1_8/Y OR2X2_62/B gnd vdd DFFPOSX1
XNAND2X1_230 AOI21X1_37/B INVX1_403/A gnd OR2X2_39/B vdd NAND2X1
XNAND2X1_252 INVX4_4/A MUX2X1_7/A gnd NAND2X1_252/Y vdd NAND2X1
XNAND2X1_241 INVX4_4/A MUX2X1_3/A gnd OAI21X1_307/C vdd NAND2X1
XFILL_5_5_0 gnd vdd FILL
XNAND2X1_263 INVX2_45/Y MUX2X1_10/Y gnd AND2X2_36/B vdd NAND2X1
XNAND2X1_285 BUFX4_77/Y MUX2X1_17/Y gnd AOI21X1_86/A vdd NAND2X1
XNAND2X1_296 INVX8_7/A AND2X2_34/A gnd AOI22X1_88/C vdd NAND2X1
XNAND2X1_274 AOI21X1_63/A NAND2X1_273/Y gnd INVX1_369/A vdd NAND2X1
XFILL_13_4_0 gnd vdd FILL
XOAI21X1_780 AND2X2_56/B MUX2X1_38/Y OAI21X1_780/C gnd OAI21X1_782/B vdd OAI21X1
XOAI21X1_791 BUFX4_177/Y INVX1_444/Y NAND2X1_614/Y gnd OAI21X1_791/Y vdd OAI21X1
XCLKBUF1_33 BUFX4_3/Y gnd CLKBUF1_33/Y vdd CLKBUF1
XCLKBUF1_11 BUFX4_1/Y gnd CLKBUF1_11/Y vdd CLKBUF1
XCLKBUF1_22 BUFX4_2/Y gnd CLKBUF1_22/Y vdd CLKBUF1
XCLKBUF1_44 BUFX4_5/Y gnd CLKBUF1_44/Y vdd CLKBUF1
XCLKBUF1_55 BUFX4_4/Y gnd CLKBUF1_55/Y vdd CLKBUF1
XINVX1_107 INVX1_107/A gnd INVX1_107/Y vdd INVX1
XINVX1_129 INVX1_129/A gnd INVX1_129/Y vdd INVX1
XINVX1_118 INVX1_118/A gnd INVX1_118/Y vdd INVX1
XINVX1_663 NOR2X1_6/B gnd INVX1_663/Y vdd INVX1
XINVX1_652 BUFX2_96/A gnd INVX1_652/Y vdd INVX1
XINVX1_641 BUFX2_87/A gnd INVX1_641/Y vdd INVX1
XINVX1_630 INVX1_557/A gnd INVX1_630/Y vdd INVX1
XINVX1_685 INVX1_685/A gnd INVX1_685/Y vdd INVX1
XINVX1_696 MUX2X1_1/B gnd INVX1_696/Y vdd INVX1
XINVX1_674 INVX1_452/A gnd INVX1_674/Y vdd INVX1
XFILL_36_3_0 gnd vdd FILL
XFILL_20_7_1 gnd vdd FILL
XFILL_2_3_0 gnd vdd FILL
XFILL_27_3_0 gnd vdd FILL
XFILL_11_7_1 gnd vdd FILL
XFILL_10_2_0 gnd vdd FILL
XBUFX4_202 BUFX4_204/A gnd BUFX4_202/Y vdd BUFX4
XBUFX4_213 INVX8_4/Y gnd BUFX4_213/Y vdd BUFX4
XBUFX4_235 BUFX4_233/A gnd BUFX4_235/Y vdd BUFX4
XBUFX4_224 INVX8_5/Y gnd AND2X2_70/B vdd BUFX4
XBUFX4_246 BUFX4_242/A gnd NOR3X1_4/A vdd BUFX4
XNOR2X1_306 INVX2_67/A INVX1_399/A gnd AND2X2_52/A vdd NOR2X1
XFILL_18_3_0 gnd vdd FILL
XBUFX4_268 BUFX4_264/A gnd BUFX4_268/Y vdd BUFX4
XBUFX4_257 AND2X2_6/Y gnd BUFX4_257/Y vdd BUFX4
XNOR2X1_317 INVX2_34/A MUX2X1_1/Y gnd NOR2X1_317/Y vdd NOR2X1
XNOR2X1_339 INVX8_3/A NOR2X1_339/B gnd NOR2X1_339/Y vdd NOR2X1
XNOR2X1_328 OR2X2_33/B NOR2X1_328/B gnd NOR2X1_328/Y vdd NOR2X1
XINVX1_471 INVX1_471/A gnd INVX1_471/Y vdd INVX1
XINVX1_460 INVX1_460/A gnd INVX1_460/Y vdd INVX1
XINVX1_482 BUFX2_58/A gnd INVX1_482/Y vdd INVX1
XINVX1_493 BUFX2_70/A gnd INVX1_493/Y vdd INVX1
XNAND2X1_807 INVX2_1/A INVX1_568/Y gnd NAND2X1_807/Y vdd NAND2X1
XNAND2X1_818 BUFX2_87/A INVX2_78/Y gnd NAND2X1_818/Y vdd NAND2X1
XNAND2X1_829 INVX1_582/Y BUFX4_94/Y gnd NAND3X1_267/C vdd NAND2X1
XNAND3X1_13 BUFX4_72/Y NAND3X1_13/B NAND3X1_13/C gnd NAND3X1_13/Y vdd NAND3X1
XNAND3X1_35 BUFX4_74/Y NAND3X1_34/Y NAND3X1_35/C gnd NAND3X1_35/Y vdd NAND3X1
XNAND3X1_24 NAND3X1_24/A BUFX4_111/Y BUFX4_139/Y gnd NAND3X1_24/Y vdd NAND3X1
XNAND3X1_46 NAND3X1_46/A INVX8_2/A BUFX4_137/Y gnd NAND3X1_47/B vdd NAND3X1
XNAND3X1_57 BUFX4_76/Y NAND3X1_57/B NAND3X1_57/C gnd NAND3X1_57/Y vdd NAND3X1
XNAND3X1_79 INVX1_234/Y NAND3X1_79/B NAND3X1_79/C gnd NAND3X1_79/Y vdd NAND3X1
XNAND3X1_68 NAND3X1_68/A BUFX4_114/Y BUFX4_136/Y gnd NAND3X1_69/B vdd NAND3X1
XNOR2X1_13 NOR2X1_13/A NOR2X1_13/B gnd NOR2X1_13/Y vdd NOR2X1
XNOR2X1_35 NOR2X1_48/A NOR2X1_35/B gnd NOR2X1_35/Y vdd NOR2X1
XNOR2X1_46 NOR2X1_46/A NOR2X1_46/B gnd NOR2X1_46/Y vdd NOR2X1
XNOR2X1_24 INVX1_66/A NOR2X1_1/A gnd NOR2X1_24/Y vdd NOR2X1
XNOR2X1_79 NOR2X1_77/Y NOR2X1_78/Y gnd AND2X2_64/B vdd NOR2X1
XNOR2X1_57 NOR2X1_57/A XOR2X1_7/B gnd NOR2X1_57/Y vdd NOR2X1
XNOR2X1_68 INVX1_230/A NOR2X1_68/B gnd NOR2X1_69/B vdd NOR2X1
XFILL_43_6_1 gnd vdd FILL
XFILL_42_1_0 gnd vdd FILL
XMUX2X1_20 MUX2X1_28/A AND2X2_28/Y MUX2X1_20/S gnd MUX2X1_20/Y vdd MUX2X1
XMUX2X1_42 MUX2X1_42/A MUX2X1_42/B INVX8_8/A gnd MUX2X1_42/Y vdd MUX2X1
XNOR2X1_103 INVX2_36/A INVX2_53/A gnd NOR2X1_103/Y vdd NOR2X1
XMUX2X1_31 MUX2X1_30/B MUX2X1_31/B INVX8_8/A gnd MUX2X1_31/Y vdd MUX2X1
XNOR2X1_114 INVX2_39/A MUX2X1_37/B gnd OAI22X1_7/D vdd NOR2X1
XMUX2X1_53 OR2X2_33/Y MUX2X1_53/B INVX8_7/A gnd MUX2X1_53/Y vdd MUX2X1
XNOR2X1_125 INVX2_45/Y NOR2X1_125/B gnd OAI22X1_24/C vdd NOR2X1
XNOR2X1_147 INVX2_46/A MUX2X1_30/B gnd NOR2X1_147/Y vdd NOR2X1
XNOR2X1_136 AND2X2_93/B INVX2_49/Y gnd INVX1_352/A vdd NOR2X1
XNOR2X1_158 INVX8_8/A INVX2_50/Y gnd NOR2X1_158/Y vdd NOR2X1
XFILL_34_6_1 gnd vdd FILL
XNOR2X1_169 INVX2_34/A INVX2_35/A gnd NAND3X1_99/C vdd NOR2X1
XFILL_23_2 gnd vdd FILL
XFILL_33_1_0 gnd vdd FILL
XOAI21X1_609 NOR2X1_308/B NOR2X1_97/Y INVX1_401/A gnd OAI21X1_609/Y vdd OAI21X1
XFILL_16_1 gnd vdd FILL
XDFFPOSX1_501 BUFX2_68/A CLKBUF1_36/Y NAND3X1_65/Y gnd vdd DFFPOSX1
XNAND2X1_604 AND2X2_56/B MUX2X1_56/Y gnd OAI21X1_780/C vdd NAND2X1
XINVX1_290 AND2X2_17/Y gnd NOR2X1_64/A vdd INVX1
XNAND2X1_626 INVX1_271/A BUFX4_265/Y gnd NAND2X1_626/Y vdd NAND2X1
XNAND2X1_615 INVX1_253/A BUFX4_267/Y gnd NAND2X1_615/Y vdd NAND2X1
XNAND2X1_648 BUFX4_245/Y XNOR2X1_15/Y gnd OAI21X1_825/C vdd NAND2X1
XNAND2X1_659 OR2X2_45/B XNOR2X1_29/Y gnd NAND2X1_659/Y vdd NAND2X1
XNAND2X1_637 NAND2X1_98/A BUFX4_267/Y gnd NAND2X1_637/Y vdd NAND2X1
XINVX1_16 gnd gnd INVX1_16/Y vdd INVX1
XINVX1_27 gnd gnd INVX1_27/Y vdd INVX1
XINVX1_38 gnd gnd INVX1_38/Y vdd INVX1
XINVX1_49 gnd gnd INVX1_49/Y vdd INVX1
XNAND2X1_90 INVX1_276/A BUFX4_161/Y gnd NAND2X1_90/Y vdd NAND2X1
XFILL_0_6_1 gnd vdd FILL
XFILL_25_6_1 gnd vdd FILL
XFILL_24_1_0 gnd vdd FILL
XAOI21X1_261 AOI21X1_263/A AOI21X1_261/B OAI22X1_56/Y gnd OAI21X1_994/A vdd AOI21X1
XAOI21X1_250 NOR2X1_432/Y OAI21X1_931/Y AOI21X1_250/C gnd AOI21X1_250/Y vdd AOI21X1
XFILL_8_7_1 gnd vdd FILL
XFILL_7_2_0 gnd vdd FILL
XFILL_16_6_1 gnd vdd FILL
XFILL_15_1_0 gnd vdd FILL
XNAND3X1_221 BUFX4_218/Y NAND3X1_221/B NAND3X1_221/C gnd NAND2X1_756/B vdd NAND3X1
XNAND3X1_210 INVX1_524/Y BUFX4_209/Y BUFX4_34/Y gnd NAND3X1_210/Y vdd NAND3X1
XNAND3X1_232 INVX1_546/Y BUFX4_210/Y BUFX4_37/Y gnd NAND3X1_232/Y vdd NAND3X1
XNAND3X1_243 BUFX4_221/Y NAND3X1_242/Y NAND3X1_243/C gnd NAND2X1_789/B vdd NAND3X1
XNAND3X1_254 NOR2X1_403/Y NOR2X1_404/Y NAND3X1_254/C gnd NAND3X1_255/B vdd NAND3X1
XNAND3X1_265 BUFX4_120/Y NAND3X1_264/Y NAND3X1_265/C gnd NAND2X1_827/B vdd NAND3X1
XNAND3X1_287 BUFX4_121/Y NAND3X1_287/B NAND3X1_287/C gnd NAND2X1_860/B vdd NAND3X1
XNAND3X1_276 INVX1_593/Y BUFX4_100/Y BUFX4_165/Y gnd NAND3X1_276/Y vdd NAND3X1
XNAND3X1_298 INVX1_615/Y BUFX4_99/Y BUFX4_167/Y gnd NAND3X1_299/B vdd NAND3X1
XOAI21X1_406 INVX8_3/A OAI21X1_398/Y OAI21X1_406/C gnd AOI21X1_59/B vdd OAI21X1
XOAI21X1_417 BUFX4_223/Y OAI21X1_344/Y OAI21X1_417/C gnd OAI21X1_419/B vdd OAI21X1
XOAI21X1_428 AOI21X1_48/Y INVX8_12/Y AOI22X1_79/Y gnd AOI21X1_65/C vdd OAI21X1
XOAI21X1_439 OR2X2_25/A OR2X2_25/B INVX8_5/A gnd OAI21X1_440/C vdd OAI21X1
XDFFPOSX1_331 INVX1_288/A CLKBUF1_1/Y OAI21X1_899/Y gnd vdd DFFPOSX1
XDFFPOSX1_320 INVX1_261/A CLKBUF1_9/Y OAI21X1_888/Y gnd vdd DFFPOSX1
XDFFPOSX1_364 OR2X2_56/A CLKBUF1_58/Y OAI21X1_21/Y gnd vdd DFFPOSX1
XDFFPOSX1_353 MUX2X1_9/B CLKBUF1_48/Y OAI21X1_10/Y gnd vdd DFFPOSX1
XDFFPOSX1_342 INVX2_3/A CLKBUF1_59/Y NOR2X1_23/A gnd vdd DFFPOSX1
XNAND2X1_401 INVX8_4/A NAND2X1_455/B gnd NAND2X1_401/Y vdd NAND2X1
XDFFPOSX1_375 INVX1_664/A CLKBUF1_48/Y OAI21X1_32/Y gnd vdd DFFPOSX1
XDFFPOSX1_386 OR2X2_59/B CLKBUF1_57/Y OAI21X1_43/Y gnd vdd DFFPOSX1
XDFFPOSX1_397 INVX1_457/A CLKBUF1_46/Y OAI21X1_54/Y gnd vdd DFFPOSX1
XNAND2X1_423 NOR2X1_214/A BUFX4_90/Y gnd AOI21X1_71/A vdd NAND2X1
XNAND2X1_434 INVX8_3/A OAI21X1_558/B gnd OAI21X1_461/C vdd NAND2X1
XNAND2X1_445 BUFX4_126/Y NOR2X1_151/B gnd AOI22X1_88/D vdd NAND2X1
XNAND2X1_412 INVX8_5/A MUX2X1_21/A gnd OAI21X1_424/C vdd NAND2X1
XNAND2X1_478 BUFX4_229/Y NAND2X1_496/B gnd OAI21X1_518/C vdd NAND2X1
XNAND2X1_456 BUFX4_78/Y OAI22X1_19/Y gnd NAND3X1_116/B vdd NAND2X1
XNAND2X1_467 BUFX4_82/Y AOI22X1_87/B gnd INVX1_382/A vdd NAND2X1
XNAND2X1_489 INVX8_4/A OAI21X1_485/B gnd NAND2X1_489/Y vdd NAND2X1
XFILL_40_4_1 gnd vdd FILL
XOAI21X1_940 INVX1_681/A INVX1_682/Y AND2X2_87/B gnd NOR3X1_72/C vdd OAI21X1
XOAI21X1_951 AOI21X1_263/A INVX2_87/A BUFX4_118/Y gnd OAI21X1_951/Y vdd OAI21X1
XOAI21X1_962 INVX8_17/Y INVX8_15/Y BUFX2_82/A gnd OAI21X1_963/C vdd OAI21X1
XOAI21X1_973 INVX1_731/Y BUFX4_115/Y OAI21X1_973/C gnd OAI21X1_973/Y vdd OAI21X1
XOAI21X1_984 INVX1_736/Y OAI21X1_992/B OAI21X1_984/C gnd AOI21X1_258/B vdd OAI21X1
XOAI21X1_995 INVX4_13/Y INVX8_16/Y data_memory_interface_data[28] gnd OAI21X1_996/C
+ vdd OAI21X1
XINVX2_70 INVX2_70/A gnd INVX2_70/Y vdd INVX2
XINVX2_81 INVX2_81/A gnd INVX2_81/Y vdd INVX2
XINVX2_92 data_memory_interface_data[8] gnd INVX2_92/Y vdd INVX2
XNAND2X1_990 INVX2_49/A AND2X2_93/B gnd OR2X2_66/A vdd NAND2X1
XOAI21X1_11 INVX1_11/Y BUFX4_22/Y OAI21X1_11/C gnd OAI21X1_11/Y vdd OAI21X1
XOAI21X1_22 INVX1_22/Y BUFX4_18/Y OAI21X1_22/C gnd OAI21X1_22/Y vdd OAI21X1
XOAI21X1_44 INVX1_44/Y BUFX4_26/Y OAI21X1_44/C gnd OAI21X1_44/Y vdd OAI21X1
XFILL_31_4_1 gnd vdd FILL
XOAI21X1_33 INVX1_33/Y BUFX4_28/Y OAI21X1_33/C gnd OAI21X1_33/Y vdd OAI21X1
XOAI21X1_77 INVX1_78/Y BUFX4_162/Y NAND2X1_79/Y gnd OAI21X1_77/Y vdd OAI21X1
XOAI21X1_66 INVX1_67/Y BUFX4_156/Y OAI21X1_66/C gnd OAI21X1_66/Y vdd OAI21X1
XOAI21X1_55 INVX1_55/Y BUFX4_29/Y OAI21X1_55/C gnd OAI21X1_55/Y vdd OAI21X1
XOAI21X1_88 INVX1_89/Y BUFX4_161/Y NAND2X1_90/Y gnd OAI21X1_88/Y vdd OAI21X1
XOAI21X1_99 OR2X2_2/A BUFX4_194/Y OAI21X1_99/C gnd OAI21X1_99/Y vdd OAI21X1
XFILL_39_5_1 gnd vdd FILL
XFILL_38_0_0 gnd vdd FILL
XFILL_22_4_1 gnd vdd FILL
XOAI21X1_203 BUFX4_141/Y INVX1_201/Y AOI22X1_18/Y gnd OAI21X1_203/Y vdd OAI21X1
XOAI21X1_247 NOR2X1_38/A NAND2X1_142/Y AOI21X1_18/Y gnd NOR2X1_36/A vdd OAI21X1
XOAI21X1_236 AOI21X1_11/Y NOR3X1_51/Y INVX1_245/Y gnd AOI21X1_13/B vdd OAI21X1
XOAI21X1_225 NOR2X1_20/B NAND2X1_109/Y NAND2X1_112/Y gnd INVX2_79/A vdd OAI21X1
XOAI21X1_214 BUFX4_142/Y INVX1_212/Y AOI22X1_29/Y gnd OAI21X1_214/Y vdd OAI21X1
XOAI21X1_269 INVX1_276/A INVX1_275/Y INVX1_277/Y gnd NAND3X1_85/A vdd OAI21X1
XOAI21X1_258 NOR3X1_55/Y OAI21X1_258/B NOR2X1_42/Y gnd AOI21X1_26/B vdd OAI21X1
XAND2X2_36 AND2X2_36/A AND2X2_36/B gnd INVX4_8/A vdd AND2X2
XAND2X2_47 AND2X2_47/A INVX2_63/A gnd OR2X2_34/A vdd AND2X2
XAND2X2_14 NOR2X1_43/Y AND2X2_14/B gnd AND2X2_14/Y vdd AND2X2
XAND2X2_25 AND2X2_25/A INVX2_51/Y gnd AND2X2_25/Y vdd AND2X2
XDFFPOSX1_172 BUFX2_15/A CLKBUF1_14/Y XNOR2X1_32/Y gnd vdd DFFPOSX1
XDFFPOSX1_161 BUFX2_4/A CLKBUF1_52/Y XNOR2X1_10/Y gnd vdd DFFPOSX1
XAND2X2_58 AND2X2_58/A INVX2_70/A gnd AND2X2_58/Y vdd AND2X2
XAND2X2_69 AND2X2_69/A AND2X2_69/B gnd AND2X2_69/Y vdd AND2X2
XDFFPOSX1_150 DFFPOSX1_38/D CLKBUF1_12/Y INVX1_296/A gnd vdd DFFPOSX1
XNAND2X1_220 INVX2_32/Y NOR2X1_160/B gnd AND2X2_51/A vdd NAND2X1
XDFFPOSX1_183 BUFX2_26/A CLKBUF1_47/Y XNOR2X1_45/Y gnd vdd DFFPOSX1
XDFFPOSX1_194 BUFX2_81/A CLKBUF1_22/Y OR2X2_61/B gnd vdd DFFPOSX1
XNAND2X1_231 INVX4_4/Y INVX1_325/Y gnd OAI21X1_299/C vdd NAND2X1
XNAND2X1_253 INVX2_42/A MUX2X1_35/A gnd AOI22X1_71/A vdd NAND2X1
XNAND2X1_242 INVX2_38/A MUX2X1_39/A gnd OAI22X1_36/B vdd NAND2X1
XNAND2X1_275 INVX8_3/A MUX2X1_11/Y gnd AOI22X1_81/B vdd NAND2X1
XFILL_5_5_1 gnd vdd FILL
XNAND2X1_264 AOI22X1_71/Y AOI22X1_72/Y gnd NOR2X1_108/A vdd NAND2X1
XNAND2X1_286 AOI21X1_86/A OAI22X1_15/B gnd INVX2_47/A vdd NAND2X1
XNAND2X1_297 INVX2_44/Y NOR2X1_249/B gnd NAND2X1_297/Y vdd NAND2X1
XFILL_4_0_0 gnd vdd FILL
XFILL_29_0_0 gnd vdd FILL
XFILL_13_4_1 gnd vdd FILL
XOAI21X1_770 INVX8_7/A OAI21X1_770/B NOR3X1_56/Y gnd OAI21X1_772/A vdd OAI21X1
XOAI21X1_781 INVX1_432/Y OAI22X1_20/A AOI22X1_109/Y gnd AOI21X1_212/C vdd OAI21X1
XOAI21X1_792 BUFX4_179/Y INVX1_445/Y NAND2X1_615/Y gnd OAI21X1_792/Y vdd OAI21X1
XCLKBUF1_12 BUFX4_6/Y gnd CLKBUF1_12/Y vdd CLKBUF1
XCLKBUF1_23 BUFX4_2/Y gnd CLKBUF1_23/Y vdd CLKBUF1
XCLKBUF1_45 BUFX4_3/Y gnd CLKBUF1_45/Y vdd CLKBUF1
XCLKBUF1_56 BUFX4_5/Y gnd CLKBUF1_56/Y vdd CLKBUF1
XCLKBUF1_34 BUFX4_1/Y gnd CLKBUF1_34/Y vdd CLKBUF1
XINVX1_108 INVX1_108/A gnd INVX1_108/Y vdd INVX1
XINVX1_119 INVX1_119/A gnd INVX1_119/Y vdd INVX1
XINVX1_620 INVX1_547/A gnd INVX1_620/Y vdd INVX1
XINVX1_653 BUFX2_97/A gnd INVX1_653/Y vdd INVX1
XINVX1_642 OAI22X1_6/Y gnd INVX1_642/Y vdd INVX1
XINVX1_631 INVX1_558/A gnd INVX1_631/Y vdd INVX1
XINVX1_686 OR2X2_62/A gnd INVX1_686/Y vdd INVX1
XINVX1_697 INVX1_697/A gnd INVX1_697/Y vdd INVX1
XINVX1_675 MUX2X1_3/B gnd INVX1_675/Y vdd INVX1
XINVX1_664 INVX1_664/A gnd INVX1_664/Y vdd INVX1
XFILL_4_1 gnd vdd FILL
XFILL_36_3_1 gnd vdd FILL
XFILL_2_3_1 gnd vdd FILL
XFILL_27_3_1 gnd vdd FILL
XFILL_10_2_1 gnd vdd FILL
XBUFX4_203 BUFX4_204/A gnd BUFX4_203/Y vdd BUFX4
XBUFX4_214 INVX8_4/Y gnd BUFX4_214/Y vdd BUFX4
XBUFX4_225 INVX8_5/Y gnd BUFX4_225/Y vdd BUFX4
XBUFX4_236 AND2X2_8/Y gnd BUFX4_236/Y vdd BUFX4
XBUFX4_247 BUFX4_242/A gnd INVX8_13/A vdd BUFX4
XNOR2X1_307 BUFX4_275/Y NOR2X1_316/B gnd NOR2X1_307/Y vdd NOR2X1
XFILL_18_3_1 gnd vdd FILL
XBUFX4_258 AND2X2_6/Y gnd BUFX4_258/Y vdd BUFX4
XBUFX4_269 NAND3X1_1/Y gnd BUFX4_269/Y vdd BUFX4
XNOR2X1_318 NOR2X1_318/A NOR2X1_318/B gnd OR2X2_37/B vdd NOR2X1
XNOR2X1_329 BUFX4_56/Y NOR2X1_329/B gnd NOR2X1_329/Y vdd NOR2X1
XINVX1_450 INVX1_450/A gnd INVX1_450/Y vdd INVX1
XINVX1_461 INVX2_81/A gnd INVX1_461/Y vdd INVX1
XINVX1_472 BUFX2_46/A gnd INVX1_472/Y vdd INVX1
XINVX1_483 BUFX2_59/A gnd INVX1_483/Y vdd INVX1
XINVX1_494 BUFX2_69/A gnd NOR3X1_68/A vdd INVX1
XNAND2X1_808 XOR2X1_1/A INVX2_76/Y gnd NAND3X1_256/B vdd NAND2X1
XNAND2X1_819 INVX2_75/A INVX1_568/Y gnd NAND2X1_819/Y vdd NAND2X1
XNAND3X1_14 NAND3X1_14/A BUFX4_111/Y BUFX4_139/Y gnd NAND3X1_15/B vdd NAND3X1
XNAND3X1_36 NAND3X1_36/A BUFX4_111/Y BUFX4_139/Y gnd NAND3X1_36/Y vdd NAND3X1
XNAND3X1_25 BUFX4_74/Y NAND3X1_24/Y NAND3X1_25/C gnd NAND3X1_25/Y vdd NAND3X1
XNAND3X1_47 BUFX4_72/Y NAND3X1_47/B NAND3X1_47/C gnd NAND3X1_47/Y vdd NAND3X1
XNAND3X1_69 BUFX4_73/Y NAND3X1_69/B NAND3X1_69/C gnd NAND3X1_69/Y vdd NAND3X1
XNAND3X1_58 NAND3X1_58/A BUFX4_114/Y BUFX4_136/Y gnd NAND3X1_59/B vdd NAND3X1
XNOR2X1_36 NOR2X1_36/A NOR2X1_35/Y gnd NOR2X1_36/Y vdd NOR2X1
XNOR2X1_25 NOR2X1_6/B OR2X2_1/B gnd NOR2X1_25/Y vdd NOR2X1
XNOR2X1_14 NOR2X1_14/A INVX1_228/A gnd NOR2X1_14/Y vdd NOR2X1
XNOR2X1_47 NOR2X1_47/A NOR2X1_47/B gnd NOR2X1_47/Y vdd NOR2X1
XNOR2X1_69 AOI21X1_5/Y NOR2X1_69/B gnd NOR2X1_69/Y vdd NOR2X1
XNOR2X1_58 INVX1_288/Y NOR2X1_58/B gnd NOR2X1_58/Y vdd NOR2X1
XFILL_42_1_1 gnd vdd FILL
XMUX2X1_10 MUX2X1_10/A INVX1_681/A INVX4_4/A gnd MUX2X1_10/Y vdd MUX2X1
XMUX2X1_21 MUX2X1_21/A MUX2X1_21/B INVX8_8/A gnd MUX2X1_21/Y vdd MUX2X1
XNOR2X1_104 OR2X2_39/B OR2X2_39/A gnd NOR2X1_104/Y vdd NOR2X1
XMUX2X1_43 MUX2X1_42/Y MUX2X1_43/B BUFX4_228/Y gnd MUX2X1_45/B vdd MUX2X1
XNOR2X1_115 INVX2_40/Y MUX2X1_5/Y gnd OAI22X1_8/B vdd NOR2X1
XMUX2X1_54 MUX2X1_54/A MUX2X1_54/B BUFX4_56/Y gnd MUX2X1_54/Y vdd MUX2X1
XMUX2X1_32 MUX2X1_32/A MUX2X1_32/B INVX8_4/A gnd MUX2X1_32/Y vdd MUX2X1
XNOR2X1_126 NOR2X1_126/A OAI22X1_9/Y gnd NOR2X1_126/Y vdd NOR2X1
XNOR2X1_148 BUFX4_77/Y MUX2X1_17/Y gnd NOR2X1_148/Y vdd NOR2X1
XNOR2X1_137 INVX2_20/Y INVX2_21/A gnd NOR2X1_137/Y vdd NOR2X1
XNOR2X1_159 BUFX4_38/Y INVX4_3/Y gnd NOR2X1_159/Y vdd NOR2X1
XFILL_33_1_1 gnd vdd FILL
XFILL_23_3 gnd vdd FILL
XFILL_16_2 gnd vdd FILL
XDFFPOSX1_502 BUFX2_69/A CLKBUF1_6/Y NAND3X1_67/Y gnd vdd DFFPOSX1
XINVX1_280 INVX1_280/A gnd INVX1_280/Y vdd INVX1
XINVX1_291 INVX1_291/A gnd INVX1_291/Y vdd INVX1
XNAND2X1_627 INVX1_273/A BUFX4_264/Y gnd NAND2X1_627/Y vdd NAND2X1
XNAND2X1_605 INVX1_230/A BUFX4_268/Y gnd NAND2X1_605/Y vdd NAND2X1
XNAND2X1_616 INVX2_9/A BUFX4_268/Y gnd NAND2X1_616/Y vdd NAND2X1
XNAND2X1_649 BUFX2_47/A NOR2X1_382/Y gnd XOR2X1_8/A vdd NAND2X1
XNAND2X1_638 NOR2X1_375/A INVX1_436/A gnd NAND2X1_638/Y vdd NAND2X1
XINVX1_17 gnd gnd INVX1_17/Y vdd INVX1
XINVX1_28 gnd gnd INVX1_28/Y vdd INVX1
XINVX1_39 gnd gnd INVX1_39/Y vdd INVX1
XNAND2X1_80 INVX1_258/A BUFX4_163/Y gnd NAND2X1_80/Y vdd NAND2X1
XNAND2X1_91 INVX1_278/A BUFX4_161/Y gnd NAND2X1_91/Y vdd NAND2X1
XFILL_24_1_1 gnd vdd FILL
XAOI21X1_251 AOI21X1_251/A AOI21X1_251/B AOI21X1_251/C gnd AOI21X1_251/Y vdd AOI21X1
XAOI21X1_240 AOI21X1_240/A OAI21X1_909/Y OAI21X1_938/A gnd AOI21X1_240/Y vdd AOI21X1
XAOI21X1_262 AOI21X1_263/A OAI21X1_996/Y OAI22X1_57/Y gnd AOI21X1_262/Y vdd AOI21X1
XFILL_7_2_1 gnd vdd FILL
XFILL_15_1_1 gnd vdd FILL
XNAND3X1_200 INVX1_514/Y BUFX4_208/Y BUFX4_36/Y gnd NAND3X1_201/B vdd NAND3X1
XNAND3X1_211 BUFX4_220/Y NAND3X1_210/Y NAND3X1_211/C gnd NAND2X1_741/B vdd NAND3X1
XNAND3X1_222 INVX1_536/Y BUFX4_208/Y BUFX4_36/Y gnd NAND3X1_223/B vdd NAND3X1
XNAND3X1_255 BUFX4_201/Y NAND3X1_255/B BUFX4_219/Y gnd BUFX4_22/A vdd NAND3X1
XNAND3X1_266 INVX1_583/Y BUFX4_100/Y BUFX4_165/Y gnd NAND3X1_266/Y vdd NAND3X1
XNAND3X1_244 INVX1_558/Y BUFX4_209/Y BUFX4_34/Y gnd NAND3X1_245/B vdd NAND3X1
XNAND3X1_233 BUFX4_222/Y NAND3X1_232/Y NAND3X1_233/C gnd NAND2X1_774/B vdd NAND3X1
XNAND3X1_277 BUFX4_120/Y NAND3X1_276/Y NAND3X1_277/C gnd NAND2X1_845/B vdd NAND3X1
XNAND3X1_288 INVX1_605/Y BUFX4_99/Y BUFX4_167/Y gnd NAND3X1_288/Y vdd NAND3X1
XNAND3X1_299 BUFX4_123/Y NAND3X1_299/B NAND3X1_299/C gnd NAND2X1_878/B vdd NAND3X1
XOAI21X1_418 INVX8_5/A AOI21X1_51/Y OAI21X1_418/C gnd NAND2X1_454/B vdd OAI21X1
XOAI21X1_429 NOR2X1_210/Y AOI22X1_78/Y AOI21X1_65/Y gnd AOI21X1_66/C vdd OAI21X1
XOAI21X1_407 AOI21X1_59/B INVX4_7/Y NAND2X1_394/Y gnd NOR2X1_200/B vdd OAI21X1
XDFFPOSX1_310 INVX1_249/A CLKBUF1_25/Y NOR2X1_415/Y gnd vdd DFFPOSX1
XDFFPOSX1_321 INVX1_264/A CLKBUF1_40/Y OAI21X1_889/Y gnd vdd DFFPOSX1
XDFFPOSX1_365 INVX1_672/A CLKBUF1_58/Y OAI21X1_22/Y gnd vdd DFFPOSX1
XDFFPOSX1_332 NOR2X1_62/A CLKBUF1_1/Y OAI21X1_900/Y gnd vdd DFFPOSX1
XDFFPOSX1_354 OR2X2_59/A CLKBUF1_57/Y OAI21X1_11/Y gnd vdd DFFPOSX1
XDFFPOSX1_343 INVX1_572/A CLKBUF1_40/Y NOR3X1_8/Y gnd vdd DFFPOSX1
XNAND2X1_402 INVX8_5/A INVX1_353/Y gnd NAND2X1_402/Y vdd NAND2X1
XDFFPOSX1_387 OR2X2_58/B CLKBUF1_46/Y OAI21X1_44/Y gnd vdd DFFPOSX1
XDFFPOSX1_376 INVX1_435/A CLKBUF1_29/Y OAI21X1_33/Y gnd vdd DFFPOSX1
XDFFPOSX1_398 INVX1_458/A CLKBUF1_29/Y OAI21X1_55/Y gnd vdd DFFPOSX1
XNAND2X1_424 BUFX4_51/Y MUX2X1_34/B gnd INVX1_374/A vdd NAND2X1
XNAND2X1_413 INVX8_8/A OAI21X1_372/Y gnd OAI21X1_424/B vdd NAND2X1
XNAND2X1_435 INVX2_56/Y NAND2X1_435/B gnd OAI22X1_20/A vdd NAND2X1
XNAND2X1_468 INVX8_4/A OAI21X1_438/A gnd OAI21X1_498/C vdd NAND2X1
XNAND2X1_457 BUFX4_223/Y MUX2X1_30/Y gnd NAND2X1_457/Y vdd NAND2X1
XNAND2X1_446 BUFX4_81/Y AND2X2_55/A gnd NOR2X1_327/B vdd NAND2X1
XNAND2X1_479 BUFX4_214/Y INVX1_395/A gnd NAND2X1_479/Y vdd NAND2X1
XOAI21X1_930 INVX1_689/Y INVX1_443/A OAI21X1_929/Y gnd OAI21X1_930/Y vdd OAI21X1
XOAI21X1_941 NAND3X1_343/Y OAI21X1_941/B INVX1_714/A gnd OAI21X1_941/Y vdd OAI21X1
XOAI21X1_952 INVX1_718/Y OAI21X1_951/Y OAI21X1_952/C gnd OAI21X1_952/Y vdd OAI21X1
XOAI21X1_963 INVX4_14/Y INVX1_723/Y OAI21X1_963/C gnd OAI21X1_963/Y vdd OAI21X1
XOAI21X1_974 INVX1_732/Y BUFX4_116/Y OAI21X1_974/C gnd OAI21X1_974/Y vdd OAI21X1
XOAI21X1_985 INVX1_736/Y OAI21X1_993/B OAI21X1_985/C gnd AOI22X1_138/C vdd OAI21X1
XOAI21X1_996 INVX1_744/Y OAI21X1_992/B OAI21X1_996/C gnd OAI21X1_996/Y vdd OAI21X1
XINVX2_60 INVX2_60/A gnd INVX2_60/Y vdd INVX2
XINVX2_71 INVX2_71/A gnd INVX2_71/Y vdd INVX2
XINVX2_82 INVX2_82/A gnd INVX2_82/Y vdd INVX2
XNAND2X1_991 INVX1_685/A INVX1_707/Y gnd NAND2X1_991/Y vdd NAND2X1
XNAND2X1_980 OR2X2_55/A INVX1_703/Y gnd OAI21X1_920/B vdd NAND2X1
XINVX2_93 INVX2_93/A gnd INVX2_93/Y vdd INVX2
XOAI21X1_23 INVX1_23/Y BUFX4_21/Y OAI21X1_23/C gnd OAI21X1_23/Y vdd OAI21X1
XOAI21X1_12 INVX1_12/Y BUFX4_22/Y OAI21X1_12/C gnd OAI21X1_12/Y vdd OAI21X1
XOAI21X1_45 INVX1_45/Y BUFX4_26/Y OAI21X1_45/C gnd OAI21X1_45/Y vdd OAI21X1
XOAI21X1_34 INVX1_34/Y BUFX4_30/Y OAI21X1_34/C gnd OAI21X1_34/Y vdd OAI21X1
XOAI21X1_78 INVX1_79/Y BUFX4_163/Y NAND2X1_80/Y gnd OAI21X1_78/Y vdd OAI21X1
XOAI21X1_67 INVX1_68/Y BUFX4_160/Y NAND2X1_69/Y gnd OAI21X1_67/Y vdd OAI21X1
XOAI21X1_56 INVX1_56/Y BUFX4_31/Y NAND2X1_56/Y gnd OAI21X1_56/Y vdd OAI21X1
XOAI21X1_89 INVX1_90/Y BUFX4_161/Y NAND2X1_91/Y gnd OAI21X1_89/Y vdd OAI21X1
XFILL_38_0_1 gnd vdd FILL
XOAI21X1_204 OR2X2_4/A INVX1_202/Y AOI22X1_19/Y gnd OAI21X1_204/Y vdd OAI21X1
XOAI21X1_237 AOI21X1_11/Y NOR3X1_51/Y INVX1_245/A gnd OAI21X1_237/Y vdd OAI21X1
XOAI21X1_215 BUFX4_141/Y INVX1_213/Y AOI22X1_30/Y gnd OAI21X1_215/Y vdd OAI21X1
XOAI21X1_226 AOI22X1_41/Y INVX1_225/A NAND3X1_74/Y gnd INVX1_643/A vdd OAI21X1
XOAI21X1_248 NOR2X1_35/Y NOR2X1_36/A NAND3X1_83/C gnd OAI21X1_249/C vdd OAI21X1
XOAI21X1_259 AOI21X1_26/Y OAI21X1_276/B NOR2X1_43/Y gnd OAI21X1_259/Y vdd OAI21X1
XAND2X2_37 MUX2X1_15/Y INVX1_342/A gnd AND2X2_37/Y vdd AND2X2
XAND2X2_15 NOR2X1_49/Y NOR2X1_45/Y gnd AND2X2_15/Y vdd AND2X2
XAND2X2_26 AND2X2_26/A INVX1_356/Y gnd OR2X2_24/B vdd AND2X2
XDFFPOSX1_151 DFFPOSX1_39/D CLKBUF1_51/Y NAND2X1_98/A gnd vdd DFFPOSX1
XAND2X2_48 AND2X2_48/A INVX1_403/A gnd AND2X2_48/Y vdd AND2X2
XDFFPOSX1_162 BUFX2_5/A CLKBUF1_26/Y XNOR2X1_12/Y gnd vdd DFFPOSX1
XDFFPOSX1_173 BUFX2_16/A CLKBUF1_14/Y XNOR2X1_35/Y gnd vdd DFFPOSX1
XAND2X2_59 AND2X2_59/A AND2X2_59/B gnd OR2X2_38/B vdd AND2X2
XDFFPOSX1_140 DFFPOSX1_28/D CLKBUF1_19/Y INVX1_271/A gnd vdd DFFPOSX1
XNAND2X1_210 INVX4_4/A AOI22X1_59/A gnd NAND2X1_210/Y vdd NAND2X1
XDFFPOSX1_184 BUFX2_27/A CLKBUF1_5/Y XNOR2X1_46/Y gnd vdd DFFPOSX1
XDFFPOSX1_195 BUFX2_82/A CLKBUF1_16/Y OR2X2_60/B gnd vdd DFFPOSX1
XNAND2X1_232 INVX4_4/A AOI22X1_53/A gnd OAI21X1_300/C vdd NAND2X1
XNAND2X1_243 INVX2_38/Y MUX2X1_3/Y gnd AOI22X1_70/B vdd NAND2X1
XNAND2X1_221 INVX1_408/A AND2X2_51/A gnd NAND3X1_89/B vdd NAND2X1
XNAND2X1_265 BUFX4_54/Y MUX2X1_11/Y gnd AOI21X1_97/A vdd NAND2X1
XNAND2X1_276 INVX8_4/A MUX2X1_12/Y gnd AOI22X1_81/C vdd NAND2X1
XNAND2X1_254 INVX2_42/Y MUX2X1_7/Y gnd AOI22X1_71/B vdd NAND2X1
XNAND2X1_287 INVX4_4/A INVX1_239/A gnd NAND2X1_287/Y vdd NAND2X1
XNAND2X1_298 INVX2_42/A MUX2X1_7/Y gnd AOI22X1_96/B vdd NAND2X1
XFILL_4_0_1 gnd vdd FILL
XFILL_29_0_1 gnd vdd FILL
XFILL_41_7_0 gnd vdd FILL
XOAI21X1_760 INVX4_7/Y NOR2X1_369/A OAI21X1_760/C gnd NOR3X1_64/B vdd OAI21X1
XOAI21X1_782 OAI22X1_30/C OAI21X1_782/B AOI21X1_212/Y gnd OAI21X1_782/Y vdd OAI21X1
XOAI21X1_771 INVX1_430/Y OAI22X1_20/A AOI22X1_108/Y gnd AOI21X1_209/C vdd OAI21X1
XOAI21X1_793 BUFX4_177/Y INVX1_446/Y NAND2X1_616/Y gnd OAI21X1_793/Y vdd OAI21X1
XFILL_32_7_0 gnd vdd FILL
XCLKBUF1_13 BUFX4_5/Y gnd CLKBUF1_13/Y vdd CLKBUF1
XCLKBUF1_24 BUFX4_1/Y gnd CLKBUF1_24/Y vdd CLKBUF1
XCLKBUF1_35 BUFX4_3/Y gnd CLKBUF1_35/Y vdd CLKBUF1
XCLKBUF1_57 BUFX4_7/Y gnd CLKBUF1_57/Y vdd CLKBUF1
XCLKBUF1_46 BUFX4_7/Y gnd CLKBUF1_46/Y vdd CLKBUF1
XFILL_23_7_0 gnd vdd FILL
XINVX1_109 INVX1_109/A gnd INVX1_109/Y vdd INVX1
XOR2X2_70 OR2X2_70/A OR2X2_70/B gnd OR2X2_70/Y vdd OR2X2
XFILL_14_7_0 gnd vdd FILL
XOAI21X1_590 AOI21X1_114/Y NOR2X1_296/B AOI21X1_129/Y gnd AOI21X1_130/C vdd OAI21X1
XINVX1_610 INVX1_537/A gnd INVX1_610/Y vdd INVX1
XINVX1_654 BUFX2_84/A gnd INVX1_654/Y vdd INVX1
XINVX1_643 INVX1_643/A gnd INVX1_643/Y vdd INVX1
XINVX1_621 INVX1_621/A gnd INVX1_621/Y vdd INVX1
XINVX1_632 INVX1_632/A gnd INVX1_632/Y vdd INVX1
XINVX1_687 OR2X2_63/A gnd OR2X2_65/A vdd INVX1
XINVX1_676 INVX1_451/A gnd INVX1_676/Y vdd INVX1
XINVX1_665 INVX1_467/A gnd INVX1_665/Y vdd INVX1
XINVX1_698 MUX2X1_2/B gnd INVX1_698/Y vdd INVX1
XFILL_4_2 gnd vdd FILL
XFILL_39_1 gnd vdd FILL
XBUFX4_204 BUFX4_204/A gnd BUFX4_204/Y vdd BUFX4
XBUFX4_215 INVX8_4/Y gnd BUFX4_215/Y vdd BUFX4
XBUFX4_226 INVX8_5/Y gnd MUX2X1_40/S vdd BUFX4
XBUFX4_237 AND2X2_8/Y gnd BUFX4_237/Y vdd BUFX4
XBUFX4_248 BUFX4_242/A gnd NOR3X1_9/A vdd BUFX4
XBUFX4_259 AND2X2_6/Y gnd BUFX4_259/Y vdd BUFX4
XNOR2X1_319 INVX2_35/A MUX2X1_2/Y gnd NOR2X1_319/Y vdd NOR2X1
XNOR2X1_308 OR2X2_39/A NOR2X1_308/B gnd NOR2X1_309/A vdd NOR2X1
XINVX1_440 OR2X2_61/B gnd INVX1_440/Y vdd INVX1
XINVX1_451 INVX1_451/A gnd INVX1_451/Y vdd INVX1
XINVX1_462 OR2X2_55/B gnd INVX1_462/Y vdd INVX1
XINVX1_473 OR2X2_46/A gnd INVX1_473/Y vdd INVX1
XINVX1_484 BUFX2_60/A gnd INVX1_484/Y vdd INVX1
XINVX1_495 INVX1_495/A gnd INVX1_495/Y vdd INVX1
XNAND2X1_809 BUFX2_87/A INVX1_569/Y gnd NAND3X1_256/C vdd NAND2X1
XFILL_37_6_0 gnd vdd FILL
XFILL_20_5_0 gnd vdd FILL
XNAND3X1_15 BUFX4_74/Y NAND3X1_15/B NAND3X1_15/C gnd NAND3X1_15/Y vdd NAND3X1
XNAND3X1_26 NAND3X1_26/A BUFX4_110/Y BUFX4_138/Y gnd NAND3X1_27/B vdd NAND3X1
XNAND3X1_37 BUFX4_74/Y NAND3X1_36/Y NAND3X1_37/C gnd NAND3X1_37/Y vdd NAND3X1
XNAND3X1_48 NAND3X1_48/A INVX8_2/A BUFX4_137/Y gnd NAND3X1_49/B vdd NAND3X1
XNAND3X1_59 BUFX4_76/Y NAND3X1_59/B NAND3X1_59/C gnd NAND3X1_59/Y vdd NAND3X1
XFILL_3_6_0 gnd vdd FILL
XNOR2X1_37 INVX2_12/Y NOR2X1_37/B gnd NOR2X1_37/Y vdd NOR2X1
XNOR2X1_26 INVX2_5/Y OR2X2_9/A gnd AOI21X1_6/C vdd NOR2X1
XFILL_28_6_0 gnd vdd FILL
XNOR2X1_15 INVX2_4/A OR2X2_5/B gnd NOR2X1_15/Y vdd NOR2X1
XNOR2X1_48 NOR2X1_48/A NOR2X1_48/B gnd NOR2X1_48/Y vdd NOR2X1
XNOR2X1_59 AND2X2_17/Y NOR2X1_59/B gnd NOR2X1_59/Y vdd NOR2X1
XFILL_11_5_0 gnd vdd FILL
XMUX2X1_11 INVX1_350/A OR2X2_62/A INVX4_4/A gnd MUX2X1_11/Y vdd MUX2X1
XFILL_19_6_0 gnd vdd FILL
XMUX2X1_33 MUX2X1_33/A MUX2X1_33/B INVX8_4/A gnd MUX2X1_33/Y vdd MUX2X1
XMUX2X1_22 MUX2X1_33/B MUX2X1_22/B INVX8_4/A gnd MUX2X1_22/Y vdd MUX2X1
XNOR2X1_105 INVX2_40/Y MUX2X1_35/B gnd OAI22X1_31/A vdd NOR2X1
XMUX2X1_44 MUX2X1_44/A MUX2X1_44/B INVX8_8/A gnd MUX2X1_47/B vdd MUX2X1
XNOR2X1_149 INVX8_6/A MUX2X1_30/A gnd NOR2X1_149/Y vdd NOR2X1
XNOR2X1_116 INVX2_40/A MUX2X1_35/B gnd OAI22X1_8/A vdd NOR2X1
XNOR2X1_127 INVX2_38/A MUX2X1_3/Y gnd OAI22X1_38/B vdd NOR2X1
XMUX2X1_55 MUX2X1_55/A MUX2X1_55/B INVX8_7/A gnd MUX2X1_55/Y vdd MUX2X1
XNOR2X1_138 INVX2_23/Y INVX2_24/A gnd NOR2X1_138/Y vdd NOR2X1
XFILL_16_3 gnd vdd FILL
XDFFPOSX1_503 BUFX2_70/A CLKBUF1_27/Y NAND3X1_69/Y gnd vdd DFFPOSX1
XINVX1_270 INVX1_270/A gnd INVX1_270/Y vdd INVX1
XINVX1_292 INVX1_292/A gnd INVX1_292/Y vdd INVX1
XINVX1_281 INVX1_281/A gnd INVX1_281/Y vdd INVX1
XNAND2X1_606 NOR2X1_375/A INVX1_436/Y gnd NAND2X1_607/A vdd NAND2X1
XNAND2X1_617 INVX2_10/A BUFX4_267/Y gnd NAND2X1_617/Y vdd NAND2X1
XNAND2X1_639 NOR2X1_69/Y NOR3X1_9/A gnd OAI21X1_815/C vdd NAND2X1
XNAND2X1_628 INVX1_274/A BUFX4_264/Y gnd NAND2X1_628/Y vdd NAND2X1
XINVX1_18 gnd gnd INVX1_18/Y vdd INVX1
XINVX1_29 gnd gnd INVX1_29/Y vdd INVX1
XNAND2X1_70 INVX2_7/A BUFX4_157/Y gnd NAND2X1_70/Y vdd NAND2X1
XNAND2X1_92 INVX1_279/A BUFX4_162/Y gnd NAND2X1_92/Y vdd NAND2X1
XNAND2X1_81 INVX2_12/A BUFX4_160/Y gnd NAND2X1_81/Y vdd NAND2X1
XAOI21X1_241 AOI21X1_241/A NOR2X1_448/Y NOR2X1_449/Y gnd INVX1_711/A vdd AOI21X1
XAOI21X1_252 AND2X2_83/A INVX1_711/Y INVX1_712/Y gnd AOI21X1_252/Y vdd AOI21X1
XAOI21X1_230 OAI22X1_6/Y INVX2_79/Y INVX8_14/Y gnd INVX4_11/A vdd AOI21X1
XAOI21X1_263 AOI21X1_263/A AOI21X1_263/B OAI22X1_58/Y gnd AOI21X1_263/Y vdd AOI21X1
XAOI22X1_90 AOI22X1_90/A AOI22X1_90/B AOI22X1_90/C BUFX4_79/Y gnd AOI22X1_90/Y vdd
+ AOI22X1
XFILL_43_4_0 gnd vdd FILL
XNAND3X1_201 BUFX4_221/Y NAND3X1_201/B NAND3X1_201/C gnd NAND2X1_726/B vdd NAND3X1
XNAND3X1_223 BUFX4_221/Y NAND3X1_223/B NAND3X1_223/C gnd NAND2X1_759/B vdd NAND3X1
XNAND3X1_212 INVX1_526/Y BUFX4_210/Y BUFX4_37/Y gnd NAND3X1_212/Y vdd NAND3X1
XNAND3X1_245 BUFX4_220/Y NAND3X1_245/B NAND3X1_245/C gnd NAND2X1_792/B vdd NAND3X1
XNAND3X1_234 INVX1_548/Y BUFX4_207/Y BUFX4_35/Y gnd NAND3X1_235/B vdd NAND3X1
XNAND3X1_256 NAND2X1_807/Y NAND3X1_256/B NAND3X1_256/C gnd NOR2X1_406/A vdd NAND3X1
XNAND3X1_278 INVX1_595/Y BUFX4_100/Y BUFX4_165/Y gnd NAND3X1_278/Y vdd NAND3X1
XNAND3X1_267 BUFX4_121/Y NAND3X1_266/Y NAND3X1_267/C gnd NAND3X1_267/Y vdd NAND3X1
XNAND3X1_289 BUFX4_123/Y NAND3X1_288/Y NAND3X1_289/C gnd NAND2X1_863/B vdd NAND3X1
XFILL_34_4_0 gnd vdd FILL
XOAI21X1_419 INVX8_4/A OAI21X1_419/B NAND2X1_405/Y gnd NOR2X1_205/B vdd OAI21X1
XOAI21X1_408 AOI21X1_53/Y INVX8_5/A OAI21X1_408/C gnd MUX2X1_28/A vdd OAI21X1
XDFFPOSX1_300 NOR2X1_133/A CLKBUF1_47/Y NOR3X1_5/Y gnd vdd DFFPOSX1
XDFFPOSX1_311 INVX2_8/A CLKBUF1_1/Y NOR2X1_416/Y gnd vdd DFFPOSX1
XDFFPOSX1_322 INVX1_268/A CLKBUF1_42/Y OAI21X1_890/Y gnd vdd DFFPOSX1
XDFFPOSX1_344 INVX1_685/A CLKBUF1_48/Y OAI21X1_1/Y gnd vdd DFFPOSX1
XDFFPOSX1_333 INVX1_296/A CLKBUF1_25/Y OAI21X1_901/Y gnd vdd DFFPOSX1
XDFFPOSX1_355 MUX2X1_7/B CLKBUF1_57/Y OAI21X1_12/Y gnd vdd DFFPOSX1
XDFFPOSX1_366 INVX1_700/A CLKBUF1_58/Y OAI21X1_23/Y gnd vdd DFFPOSX1
XDFFPOSX1_388 OR2X2_57/B CLKBUF1_46/Y OAI21X1_45/Y gnd vdd DFFPOSX1
XDFFPOSX1_377 OR2X2_64/B CLKBUF1_37/Y OAI21X1_34/Y gnd vdd DFFPOSX1
XNAND2X1_436 AOI22X1_83/Y AOI21X1_75/Y gnd AOI21X1_80/C vdd NAND2X1
XNAND2X1_425 BUFX4_54/Y MUX2X1_24/B gnd AOI22X1_81/A vdd NAND2X1
XNAND2X1_403 BUFX4_223/Y OAI21X1_343/A gnd OAI21X1_417/C vdd NAND2X1
XNAND2X1_414 BUFX4_82/Y NOR2X1_209/Y gnd INVX1_372/A vdd NAND2X1
XDFFPOSX1_399 INVX1_459/A CLKBUF1_29/Y OAI21X1_56/Y gnd vdd DFFPOSX1
XNAND2X1_458 INVX8_4/A NAND2X1_409/B gnd OAI21X1_485/C vdd NAND2X1
XNAND2X1_469 INVX8_3/A INVX1_384/Y gnd OAI21X1_499/C vdd NAND2X1
XNAND2X1_447 BUFX4_84/Y INVX2_54/A gnd OAI22X1_27/A vdd NAND2X1
XFILL_0_4_0 gnd vdd FILL
XFILL_25_4_0 gnd vdd FILL
XNOR2X1_480 NOR3X1_77/Y NOR3X1_74/Y gnd NOR2X1_480/Y vdd NOR2X1
XOAI21X1_931 AOI21X1_246/Y OR2X2_68/A AOI21X1_247/Y gnd OAI21X1_931/Y vdd OAI21X1
XOAI21X1_920 NOR2X1_451/Y OAI21X1_920/B NAND2X1_979/Y gnd AOI21X1_244/C vdd OAI21X1
XOAI21X1_942 NOR3X1_74/Y NOR3X1_73/Y INVX4_12/Y gnd INVX2_93/A vdd OAI21X1
XOAI21X1_953 INVX1_718/Y INVX4_14/A OAI21X1_953/C gnd OAI21X1_953/Y vdd OAI21X1
XOAI21X1_964 INVX8_17/Y INVX8_15/Y BUFX2_83/A gnd OAI21X1_965/C vdd OAI21X1
XOAI21X1_975 NOR3X1_77/Y NOR3X1_78/Y INVX8_16/A gnd OAI21X1_992/B vdd OAI21X1
XOAI21X1_997 INVX1_744/Y OAI21X1_993/B OAI21X1_997/C gnd AOI22X1_141/C vdd OAI21X1
XOAI21X1_986 OAI21X1_986/A OAI21X1_994/B AOI22X1_138/Y gnd OAI21X1_986/Y vdd OAI21X1
XFILL_8_5_0 gnd vdd FILL
XINVX2_72 INVX2_72/A gnd INVX2_72/Y vdd INVX2
XINVX2_61 INVX2_61/A gnd INVX2_61/Y vdd INVX2
XINVX2_50 INVX2_50/A gnd INVX2_50/Y vdd INVX2
XNAND2X1_992 NOR2X1_461/Y NOR2X1_432/Y gnd NAND2X1_992/Y vdd NAND2X1
XINVX2_83 INVX2_83/A gnd INVX2_83/Y vdd INVX2
XNAND2X1_970 NAND2X1_970/A AOI21X1_245/A gnd NOR2X1_442/A vdd NAND2X1
XNAND2X1_981 AND2X2_81/Y NOR2X1_422/Y gnd NAND2X1_981/Y vdd NAND2X1
XFILL_16_4_0 gnd vdd FILL
XOAI21X1_24 INVX1_24/Y BUFX4_21/Y OAI21X1_24/C gnd OAI21X1_24/Y vdd OAI21X1
XOAI21X1_13 INVX1_13/Y BUFX4_23/Y OAI21X1_13/C gnd OAI21X1_13/Y vdd OAI21X1
XOAI21X1_35 INVX1_35/Y BUFX4_26/Y NAND2X1_35/Y gnd OAI21X1_35/Y vdd OAI21X1
XOAI21X1_68 INVX1_69/Y BUFX4_157/Y NAND2X1_70/Y gnd OAI21X1_68/Y vdd OAI21X1
XOAI21X1_46 INVX1_46/Y BUFX4_32/Y NAND2X1_46/Y gnd OAI21X1_46/Y vdd OAI21X1
XOAI21X1_57 INVX1_57/Y BUFX4_27/Y NAND2X1_57/Y gnd OAI21X1_57/Y vdd OAI21X1
XOAI21X1_79 INVX1_80/Y BUFX4_160/Y NAND2X1_81/Y gnd OAI21X1_79/Y vdd OAI21X1
XOAI21X1_238 AOI21X1_10/Y INVX1_248/Y OAI21X1_237/Y gnd XNOR2X1_15/A vdd OAI21X1
XOAI21X1_227 NAND3X1_76/Y AOI21X1_4/C AOI21X1_8/A gnd BUFX4_148/A vdd OAI21X1
XOAI21X1_216 BUFX4_144/Y INVX1_214/Y AOI22X1_31/Y gnd OAI21X1_216/Y vdd OAI21X1
XOAI21X1_205 BUFX4_144/Y INVX1_203/Y AOI22X1_20/Y gnd OAI21X1_205/Y vdd OAI21X1
XOAI21X1_249 INVX2_11/Y XNOR2X1_28/A OAI21X1_249/C gnd XNOR2X1_30/A vdd OAI21X1
XAND2X2_38 AND2X2_38/A BUFX4_53/Y gnd AND2X2_38/Y vdd AND2X2
XAND2X2_16 AND2X2_16/A AND2X2_16/B gnd AND2X2_16/Y vdd AND2X2
XAND2X2_27 AND2X2_27/A AND2X2_27/B gnd AND2X2_27/Y vdd AND2X2
XDFFPOSX1_130 DFFPOSX1_18/D CLKBUF1_4/Y INVX2_9/A gnd vdd DFFPOSX1
XDFFPOSX1_163 BUFX2_6/A CLKBUF1_35/Y XNOR2X1_13/Y gnd vdd DFFPOSX1
XAND2X2_49 AND2X2_49/A INVX2_65/A gnd NOR3X1_58/B vdd AND2X2
XDFFPOSX1_141 DFFPOSX1_29/D CLKBUF1_40/Y INVX1_273/A gnd vdd DFFPOSX1
XDFFPOSX1_152 INVX2_75/A CLKBUF1_39/Y INVX2_1/A gnd vdd DFFPOSX1
XDFFPOSX1_174 BUFX2_17/A CLKBUF1_41/Y XNOR2X1_36/Y gnd vdd DFFPOSX1
XNAND2X1_211 INVX2_29/Y INVX2_30/Y gnd AOI22X1_69/C vdd NAND2X1
XNAND2X1_200 NOR2X1_80/A INVX2_50/A gnd INVX2_19/A vdd NAND2X1
XDFFPOSX1_185 BUFX2_28/A CLKBUF1_44/Y XOR2X1_7/Y gnd vdd DFFPOSX1
XDFFPOSX1_196 BUFX2_83/A CLKBUF1_16/Y INVX1_442/A gnd vdd DFFPOSX1
XNAND2X1_233 INVX4_4/A AOI22X1_54/A gnd NAND2X1_233/Y vdd NAND2X1
XNAND2X1_244 INVX4_4/A MUX2X1_4/A gnd NAND2X1_244/Y vdd NAND2X1
XNAND2X1_222 INVX4_4/A MUX2X1_1/A gnd NAND2X1_222/Y vdd NAND2X1
XNAND2X1_266 INVX4_4/A INVX1_350/A gnd NAND2X1_266/Y vdd NAND2X1
XNAND2X1_255 INVX4_4/A MUX2X1_8/A gnd NAND2X1_255/Y vdd NAND2X1
XNAND2X1_277 INVX4_4/A INVX1_251/A gnd NAND2X1_277/Y vdd NAND2X1
XNAND2X1_288 INVX8_7/A NOR2X1_151/B gnd OAI21X1_463/A vdd NAND2X1
XNAND2X1_299 INVX2_42/Y MUX2X1_35/A gnd AOI22X1_96/A vdd NAND2X1
XFILL_41_7_1 gnd vdd FILL
XFILL_40_2_0 gnd vdd FILL
XOAI21X1_750 INVX1_305/A OAI21X1_750/B OAI21X1_750/C gnd INVX1_427/A vdd OAI21X1
XOAI21X1_761 OAI21X1_759/Y NOR2X1_368/Y NOR3X1_64/Y gnd OAI21X1_761/Y vdd OAI21X1
XOAI21X1_772 OAI21X1_772/A NOR2X1_373/Y AOI21X1_209/Y gnd AOI21X1_210/C vdd OAI21X1
XOAI21X1_783 OAI21X1_783/A INVX1_434/A INVX2_26/Y gnd NAND3X1_177/C vdd OAI21X1
XOAI21X1_794 BUFX4_178/Y INVX1_447/Y NAND2X1_617/Y gnd OAI21X1_794/Y vdd OAI21X1
XFILL_32_7_1 gnd vdd FILL
XFILL_31_2_0 gnd vdd FILL
XCLKBUF1_14 BUFX4_3/Y gnd CLKBUF1_14/Y vdd CLKBUF1
XCLKBUF1_36 BUFX4_5/Y gnd CLKBUF1_36/Y vdd CLKBUF1
XCLKBUF1_47 BUFX4_5/Y gnd CLKBUF1_47/Y vdd CLKBUF1
XCLKBUF1_25 BUFX4_6/Y gnd CLKBUF1_25/Y vdd CLKBUF1
XCLKBUF1_58 BUFX4_6/Y gnd CLKBUF1_58/Y vdd CLKBUF1
XFILL_39_3_0 gnd vdd FILL
XBUFX4_90 BUFX4_93/A gnd BUFX4_90/Y vdd BUFX4
XFILL_23_7_1 gnd vdd FILL
XFILL_22_2_0 gnd vdd FILL
XOR2X2_60 INVX2_85/A OR2X2_60/B gnd OR2X2_60/Y vdd OR2X2
XFILL_5_3_0 gnd vdd FILL
XFILL_14_7_1 gnd vdd FILL
XFILL_13_2_0 gnd vdd FILL
XOAI21X1_591 INVX1_399/A OAI21X1_694/A AOI21X1_131/Y gnd OAI21X1_591/Y vdd OAI21X1
XOAI21X1_580 OAI22X1_38/A OAI22X1_38/B NOR2X1_293/Y gnd NAND3X1_138/C vdd OAI21X1
XINVX1_611 INVX1_611/A gnd INVX1_611/Y vdd INVX1
XINVX1_600 INVX1_527/A gnd INVX1_600/Y vdd INVX1
XINVX1_644 INVX2_76/A gnd INVX1_644/Y vdd INVX1
XINVX1_622 INVX1_549/A gnd INVX1_622/Y vdd INVX1
XINVX1_633 INVX1_560/A gnd INVX1_633/Y vdd INVX1
XINVX1_688 OR2X2_61/A gnd INVX1_688/Y vdd INVX1
XINVX1_655 BUFX2_85/A gnd INVX1_655/Y vdd INVX1
XINVX1_677 INVX1_450/A gnd INVX1_677/Y vdd INVX1
XINVX1_666 INVX1_666/A gnd INVX1_666/Y vdd INVX1
XINVX1_699 INVX1_699/A gnd INVX1_699/Y vdd INVX1
XFILL_4_3 gnd vdd FILL
XFILL_39_2 gnd vdd FILL
XBUFX4_216 INVX8_4/Y gnd BUFX4_216/Y vdd BUFX4
XBUFX4_227 INVX8_5/Y gnd BUFX4_227/Y vdd BUFX4
XBUFX4_205 BUFX4_204/A gnd BUFX4_205/Y vdd BUFX4
XBUFX4_249 BUFX4_242/A gnd NOR3X1_3/A vdd BUFX4
XBUFX4_238 AND2X2_8/Y gnd BUFX4_238/Y vdd BUFX4
XNOR2X1_309 NOR2X1_309/A NOR2X1_309/B gnd NOR2X1_309/Y vdd NOR2X1
XINVX1_430 NOR2X1_93/B gnd INVX1_430/Y vdd INVX1
XINVX1_441 OR2X2_60/B gnd INVX1_441/Y vdd INVX1
XINVX1_452 INVX1_452/A gnd INVX1_452/Y vdd INVX1
XINVX1_474 BUFX2_49/A gnd INVX1_474/Y vdd INVX1
XINVX1_485 BUFX2_61/A gnd INVX1_485/Y vdd INVX1
XINVX1_463 OR2X2_54/B gnd INVX1_463/Y vdd INVX1
XINVX1_496 INVX2_1/A gnd INVX1_496/Y vdd INVX1
XFILL_37_6_1 gnd vdd FILL
XFILL_36_1_0 gnd vdd FILL
XFILL_20_5_1 gnd vdd FILL
XNAND3X1_38 NAND3X1_38/A INVX8_2/A BUFX4_137/Y gnd NAND3X1_39/B vdd NAND3X1
XNAND3X1_16 NAND3X1_16/A BUFX4_111/Y BUFX4_139/Y gnd NAND3X1_17/B vdd NAND3X1
XNAND3X1_27 BUFX4_75/Y NAND3X1_27/B NAND3X1_27/C gnd NAND3X1_27/Y vdd NAND3X1
XNAND3X1_49 BUFX4_73/Y NAND3X1_49/B NAND3X1_49/C gnd NAND3X1_49/Y vdd NAND3X1
XNOR2X1_27 INVX2_6/Y XNOR2X1_6/A gnd AOI21X1_7/A vdd NOR2X1
XFILL_28_6_1 gnd vdd FILL
XNOR2X1_16 OR2X2_5/B NOR2X1_16/B gnd NOR2X1_16/Y vdd NOR2X1
XNOR2X1_38 NOR2X1_38/A NOR2X1_38/B gnd NOR2X1_38/Y vdd NOR2X1
XFILL_3_6_1 gnd vdd FILL
XFILL_2_1_0 gnd vdd FILL
XNOR2X1_49 XOR2X1_5/B NOR2X1_49/B gnd NOR2X1_49/Y vdd NOR2X1
XFILL_27_1_0 gnd vdd FILL
XFILL_11_5_1 gnd vdd FILL
XFILL_10_0_0 gnd vdd FILL
XFILL_19_6_1 gnd vdd FILL
XMUX2X1_12 INVX1_351/A OR2X2_63/A INVX4_4/A gnd MUX2X1_12/Y vdd MUX2X1
XMUX2X1_34 MUX2X1_34/A MUX2X1_34/B BUFX4_51/Y gnd INVX2_60/A vdd MUX2X1
XMUX2X1_23 MUX2X1_23/A MUX2X1_23/B BUFX4_223/Y gnd INVX1_383/A vdd MUX2X1
XNOR2X1_106 INVX2_40/A MUX2X1_5/Y gnd OAI22X1_31/B vdd NOR2X1
XMUX2X1_45 MUX2X1_45/A MUX2X1_45/B MUX2X1_20/S gnd MUX2X1_45/Y vdd MUX2X1
XFILL_18_1_0 gnd vdd FILL
XNOR2X1_117 INVX2_41/Y MUX2X1_6/Y gnd OAI22X1_8/C vdd NOR2X1
XMUX2X1_56 AND2X2_74/A MUX2X1_56/B BUFX4_55/Y gnd MUX2X1_56/Y vdd MUX2X1
XNOR2X1_128 NOR2X1_1/A OR2X2_16/A gnd NOR2X1_128/Y vdd NOR2X1
XNOR2X1_139 NOR2X1_76/A INVX4_2/Y gnd INVX1_349/A vdd NOR2X1
XINVX1_260 INVX1_260/A gnd INVX1_260/Y vdd INVX1
XINVX1_271 INVX1_271/A gnd OR2X2_12/B vdd INVX1
XINVX1_293 INVX1_293/A gnd INVX1_293/Y vdd INVX1
XINVX1_282 INVX1_282/A gnd INVX1_282/Y vdd INVX1
XNAND2X1_607 NAND2X1_607/A INVX1_437/Y gnd BUFX4_178/A vdd NAND2X1
XNAND2X1_618 INVX2_11/A BUFX4_267/Y gnd NAND2X1_618/Y vdd NAND2X1
XNAND2X1_629 INVX1_276/A BUFX4_264/Y gnd NAND2X1_629/Y vdd NAND2X1
XINVX1_19 gnd gnd INVX1_19/Y vdd INVX1
XNAND2X1_60 BUFX4_28/Y NAND2X1_60/B gnd OAI21X1_60/C vdd NAND2X1
XNAND2X1_71 INVX1_234/A BUFX4_160/Y gnd NAND2X1_71/Y vdd NAND2X1
XNAND2X1_82 INVX2_13/A BUFX4_159/Y gnd OAI21X1_80/C vdd NAND2X1
XNAND2X1_93 INVX1_283/A BUFX4_160/Y gnd OAI21X1_91/C vdd NAND2X1
XAOI21X1_220 BUFX2_65/A NOR3X1_66/Y BUFX2_66/A gnd AOI21X1_220/Y vdd AOI21X1
XAOI21X1_242 NAND2X1_939/Y NOR2X1_450/Y INVX1_699/A gnd INVX1_712/A vdd AOI21X1
XAOI21X1_231 OAI22X1_6/Y NOR2X1_412/Y NOR2X1_411/Y gnd AOI21X1_231/Y vdd AOI21X1
XAOI21X1_264 AOI21X1_263/A AOI21X1_264/B OAI22X1_59/Y gnd AOI21X1_264/Y vdd AOI21X1
XAOI21X1_253 NOR2X1_442/Y OAI21X1_935/Y INVX1_705/A gnd OAI21X1_936/C vdd AOI21X1
XAOI22X1_80 AOI22X1_80/A BUFX4_153/Y NOR2X1_194/Y AOI22X1_80/D gnd AOI22X1_80/Y vdd
+ AOI22X1
XAOI22X1_91 INVX4_5/Y AOI22X1_91/B AOI22X1_91/C BUFX4_79/Y gnd AOI22X1_91/Y vdd AOI22X1
XFILL_43_4_1 gnd vdd FILL
XNAND3X1_202 INVX1_516/Y BUFX4_209/Y BUFX4_34/Y gnd NAND3X1_203/B vdd NAND3X1
XNAND3X1_213 BUFX4_222/Y NAND3X1_212/Y NAND2X1_743/Y gnd NAND2X1_744/B vdd NAND3X1
XNAND3X1_235 BUFX4_219/Y NAND3X1_235/B NAND3X1_235/C gnd NAND2X1_777/B vdd NAND3X1
XNAND3X1_224 INVX1_538/Y BUFX4_207/Y BUFX4_35/Y gnd NAND3X1_224/Y vdd NAND3X1
XNAND3X1_257 NAND3X1_257/A NAND3X1_257/B AOI21X1_226/Y gnd NOR2X1_406/B vdd NAND3X1
XNAND3X1_246 INVX1_560/Y BUFX4_210/Y BUFX4_37/Y gnd NAND3X1_246/Y vdd NAND3X1
XNAND3X1_279 BUFX4_121/Y NAND3X1_278/Y NAND3X1_279/C gnd NAND2X1_848/B vdd NAND3X1
XNAND3X1_268 INVX1_585/Y BUFX4_100/Y BUFX4_165/Y gnd NAND3X1_269/B vdd NAND3X1
XFILL_34_4_1 gnd vdd FILL
XOAI21X1_409 NOR2X1_158/Y NOR2X1_159/Y INVX8_5/A gnd OAI21X1_410/C vdd OAI21X1
XDFFPOSX1_301 OR2X2_22/B CLKBUF1_58/Y NOR3X1_6/Y gnd vdd DFFPOSX1
XDFFPOSX1_312 INVX1_253/A CLKBUF1_25/Y NOR2X1_417/Y gnd vdd DFFPOSX1
XDFFPOSX1_334 NAND2X1_98/A CLKBUF1_12/Y INVX8_14/A gnd vdd DFFPOSX1
XDFFPOSX1_345 OR2X2_64/A CLKBUF1_48/Y OAI21X1_2/Y gnd vdd DFFPOSX1
XDFFPOSX1_356 OR2X2_57/A CLKBUF1_48/Y OAI21X1_13/Y gnd vdd DFFPOSX1
XDFFPOSX1_323 INVX1_271/A CLKBUF1_1/Y OAI21X1_891/Y gnd vdd DFFPOSX1
XDFFPOSX1_367 INVX2_82/A CLKBUF1_4/Y OAI21X1_24/Y gnd vdd DFFPOSX1
XDFFPOSX1_378 OR2X2_63/B CLKBUF1_46/Y OAI21X1_35/Y gnd vdd DFFPOSX1
XDFFPOSX1_389 INVX1_449/A CLKBUF1_8/Y OAI21X1_46/Y gnd vdd DFFPOSX1
XNAND2X1_426 AOI22X1_81/B AOI22X1_81/A gnd NAND2X1_426/Y vdd NAND2X1
XNAND2X1_415 INVX8_5/A INVX1_366/A gnd NAND2X1_415/Y vdd NAND2X1
XNAND2X1_404 INVX8_5/A OR2X2_19/A gnd OAI21X1_418/C vdd NAND2X1
XNAND2X1_437 INVX8_5/A MUX2X1_25/B gnd OAI21X1_470/C vdd NAND2X1
XNAND2X1_448 INVX2_46/Y MUX2X1_30/B gnd AOI22X1_89/D vdd NAND2X1
XNAND2X1_459 BUFX4_57/Y AOI22X1_98/A gnd NOR2X1_229/B vdd NAND2X1
XFILL_0_4_1 gnd vdd FILL
XFILL_25_4_1 gnd vdd FILL
XNOR2X1_470 AND2X2_99/B INVX8_15/Y gnd NOR2X1_470/Y vdd NOR2X1
XNOR2X1_481 NOR3X1_73/Y NOR3X1_74/Y gnd NOR2X1_481/Y vdd NOR2X1
XOAI21X1_943 AOI21X1_259/B INVX4_12/Y NAND3X1_352/Y gnd NOR2X1_475/A vdd OAI21X1
XOAI21X1_932 OAI21X1_932/A INVX1_691/A AOI21X1_249/Y gnd AOI21X1_250/C vdd OAI21X1
XOAI21X1_910 NOR2X1_431/Y AND2X2_87/A AND2X2_87/B gnd OAI21X1_910/Y vdd OAI21X1
XOAI21X1_921 INVX1_668/A INVX2_80/Y NOR2X1_453/Y gnd AND2X2_92/A vdd OAI21X1
XOAI21X1_954 INVX8_17/Y INVX8_15/Y BUFX2_78/A gnd OAI21X1_955/C vdd OAI21X1
XOAI21X1_965 INVX4_14/Y INVX1_724/Y OAI21X1_965/C gnd OAI21X1_965/Y vdd OAI21X1
XOAI21X1_976 INVX4_13/Y INVX8_16/Y data_memory_interface_data[24] gnd OAI21X1_977/C
+ vdd OAI21X1
XOAI21X1_998 AOI21X1_262/Y OAI21X1_994/B OAI21X1_998/C gnd OAI21X1_998/Y vdd OAI21X1
XOAI21X1_987 INVX4_13/Y INVX8_16/Y data_memory_interface_data[26] gnd OAI21X1_987/Y
+ vdd OAI21X1
XFILL_8_5_1 gnd vdd FILL
XFILL_7_0_0 gnd vdd FILL
XINVX2_40 INVX2_40/A gnd INVX2_40/Y vdd INVX2
XINVX2_62 OR2X2_40/A gnd INVX2_62/Y vdd INVX2
XINVX2_51 INVX2_51/A gnd INVX2_51/Y vdd INVX2
XINVX2_73 INVX2_73/A gnd INVX2_73/Y vdd INVX2
XNAND2X1_960 OR2X2_62/B INVX1_686/Y gnd AOI21X1_234/A vdd NAND2X1
XNAND2X1_971 AND2X2_81/A AND2X2_81/B gnd NOR2X1_442/B vdd NAND2X1
XNAND2X1_982 INVX1_668/A INVX2_80/Y gnd AND2X2_92/B vdd NAND2X1
XINVX2_84 INVX2_84/A gnd INVX2_84/Y vdd INVX2
XNAND2X1_993 NAND2X1_993/A OAI21X1_938/Y gnd NAND2X1_993/Y vdd NAND2X1
XFILL_16_4_1 gnd vdd FILL
XOAI21X1_25 INVX1_25/Y BUFX4_21/Y OAI21X1_25/C gnd OAI21X1_25/Y vdd OAI21X1
XOAI21X1_14 INVX1_14/Y BUFX4_23/Y OAI21X1_14/C gnd OAI21X1_14/Y vdd OAI21X1
XOAI21X1_69 INVX1_70/Y BUFX4_160/Y NAND2X1_71/Y gnd OAI21X1_69/Y vdd OAI21X1
XOAI21X1_47 INVX1_47/Y BUFX4_29/Y OAI21X1_47/C gnd OAI21X1_47/Y vdd OAI21X1
XOAI21X1_58 INVX1_58/Y BUFX4_26/Y NAND2X1_58/Y gnd OAI21X1_58/Y vdd OAI21X1
XOAI21X1_36 INVX1_36/Y BUFX4_27/Y NAND2X1_36/Y gnd OAI21X1_36/Y vdd OAI21X1
XOAI21X1_228 AOI21X1_6/Y XNOR2X1_8/Y INVX1_233/Y gnd XNOR2X1_10/A vdd OAI21X1
XOAI21X1_217 BUFX4_144/Y INVX1_215/Y AOI22X1_32/Y gnd OAI21X1_217/Y vdd OAI21X1
XOAI21X1_206 BUFX4_145/Y INVX1_204/Y AOI22X1_21/Y gnd OAI21X1_206/Y vdd OAI21X1
XOAI21X1_239 AOI21X1_12/Y NOR3X1_52/Y INVX1_249/A gnd OAI21X1_239/Y vdd OAI21X1
XAND2X2_28 MUX2X1_19/A AND2X2_70/B gnd AND2X2_28/Y vdd AND2X2
XAND2X2_17 INVX1_289/Y AND2X2_17/B gnd AND2X2_17/Y vdd AND2X2
XDFFPOSX1_120 DFFPOSX1_8/D CLKBUF1_32/Y INVX1_230/A gnd vdd DFFPOSX1
XDFFPOSX1_153 INVX1_501/A CLKBUF1_43/Y XOR2X1_1/A gnd vdd DFFPOSX1
XDFFPOSX1_164 BUFX2_7/A CLKBUF1_35/Y XNOR2X1_14/Y gnd vdd DFFPOSX1
XAND2X2_39 AND2X2_38/Y BUFX4_84/Y gnd AND2X2_39/Y vdd AND2X2
XDFFPOSX1_142 DFFPOSX1_30/D CLKBUF1_32/Y INVX1_274/A gnd vdd DFFPOSX1
XDFFPOSX1_131 DFFPOSX1_19/D CLKBUF1_32/Y INVX2_10/A gnd vdd DFFPOSX1
XDFFPOSX1_175 BUFX2_18/A CLKBUF1_54/Y XOR2X1_3/Y gnd vdd DFFPOSX1
XDFFPOSX1_186 BUFX2_29/A CLKBUF1_5/Y NOR2X1_60/Y gnd vdd DFFPOSX1
XNAND2X1_201 NOR2X1_82/Y INVX1_305/Y gnd OR2X2_15/B vdd NAND2X1
XDFFPOSX1_197 OAI21X1_966/C CLKBUF1_38/Y INVX1_443/A gnd vdd DFFPOSX1
XNAND2X1_223 INVX4_4/A MUX2X1_2/A gnd NAND2X1_223/Y vdd NAND2X1
XNAND2X1_234 AND2X2_59/B AND2X2_59/A gnd AOI21X1_38/B vdd NAND2X1
XNAND2X1_212 INVX2_29/A INVX2_30/A gnd INVX1_412/A vdd NAND2X1
XNAND2X1_267 INVX8_3/A MUX2X1_24/B gnd AOI22X1_73/A vdd NAND2X1
XNAND2X1_256 INVX2_43/A NOR2X1_123/B gnd OAI22X1_25/C vdd NAND2X1
XNAND2X1_278 INVX1_342/A MUX2X1_31/B gnd AOI22X1_74/A vdd NAND2X1
XNAND2X1_245 INVX2_39/A MUX2X1_37/B gnd AOI22X1_70/C vdd NAND2X1
XNAND2X1_289 BUFX4_126/Y AND2X2_34/A gnd AOI22X1_82/A vdd NAND2X1
XFILL_40_2_1 gnd vdd FILL
XOAI21X1_740 OAI22X1_30/C MUX2X1_51/Y NOR2X1_352/Y gnd AOI21X1_198/C vdd OAI21X1
XOAI21X1_751 OAI21X1_698/B OR2X2_15/B INVX1_427/Y gnd NOR2X1_362/B vdd OAI21X1
XOAI21X1_762 INVX1_428/Y NOR2X1_138/Y INVX2_22/A gnd INVX1_429/A vdd OAI21X1
XOAI21X1_784 BUFX4_177/Y INVX1_435/Y NAND2X1_605/Y gnd OAI21X1_784/Y vdd OAI21X1
XOAI21X1_773 NOR2X1_366/B INVX1_311/A OAI21X1_773/C gnd OR2X2_43/A vdd OAI21X1
XOAI21X1_795 BUFX4_179/Y INVX1_448/Y NAND2X1_618/Y gnd OAI21X1_795/Y vdd OAI21X1
XNAND2X1_790 OAI21X1_92/Y BUFX4_131/Y gnd NAND2X1_790/Y vdd NAND2X1
XFILL_31_2_1 gnd vdd FILL
XCLKBUF1_15 BUFX4_7/Y gnd CLKBUF1_15/Y vdd CLKBUF1
XCLKBUF1_26 BUFX4_3/Y gnd CLKBUF1_26/Y vdd CLKBUF1
XCLKBUF1_48 BUFX4_7/Y gnd CLKBUF1_48/Y vdd CLKBUF1
XCLKBUF1_37 BUFX4_7/Y gnd CLKBUF1_37/Y vdd CLKBUF1
XCLKBUF1_59 BUFX4_1/Y gnd CLKBUF1_59/Y vdd CLKBUF1
XFILL_39_3_1 gnd vdd FILL
XBUFX4_80 INVX8_6/Y gnd BUFX4_80/Y vdd BUFX4
XBUFX4_91 BUFX4_93/A gnd BUFX4_91/Y vdd BUFX4
XFILL_22_2_1 gnd vdd FILL
XOR2X2_50 OR2X2_50/A OR2X2_50/B gnd OR2X2_50/Y vdd OR2X2
XOR2X2_61 OR2X2_61/A OR2X2_61/B gnd OR2X2_61/Y vdd OR2X2
XXNOR2X1_1 XOR2X1_2/A BUFX2_90/A gnd AND2X2_3/A vdd XNOR2X1
XFILL_5_3_1 gnd vdd FILL
XFILL_13_2_1 gnd vdd FILL
XINVX1_1 gnd gnd INVX1_1/Y vdd INVX1
XOAI21X1_570 BUFX4_52/Y NOR2X1_222/B OAI21X1_570/C gnd NOR2X1_368/B vdd OAI21X1
XOAI21X1_592 OAI22X1_9/Y OAI21X1_529/C AOI21X1_132/Y gnd AOI21X1_134/B vdd OAI21X1
XOAI21X1_581 AND2X2_46/Y NOR2X1_293/A INVX2_64/Y gnd NAND3X1_138/B vdd OAI21X1
XINVX1_601 INVX1_601/A gnd INVX1_601/Y vdd INVX1
XINVX1_634 INVX1_561/A gnd INVX1_634/Y vdd INVX1
XINVX1_645 OR2X2_52/B gnd INVX1_645/Y vdd INVX1
XINVX1_623 INVX1_623/A gnd INVX1_623/Y vdd INVX1
XINVX1_612 INVX1_539/A gnd INVX1_612/Y vdd INVX1
XINVX1_678 MUX2X1_4/B gnd INVX1_678/Y vdd INVX1
XINVX1_656 BUFX2_86/A gnd INVX1_656/Y vdd INVX1
XINVX1_667 INVX1_667/A gnd INVX1_667/Y vdd INVX1
XINVX1_689 INVX1_689/A gnd INVX1_689/Y vdd INVX1
XFILL_39_3 gnd vdd FILL
XBUFX4_228 INVX8_5/Y gnd BUFX4_228/Y vdd BUFX4
XBUFX4_217 INVX8_4/Y gnd BUFX4_217/Y vdd BUFX4
XBUFX4_206 BUFX4_210/A gnd BUFX4_206/Y vdd BUFX4
XBUFX4_239 AND2X2_8/Y gnd AOI22X1_9/B vdd BUFX4
XAND2X2_1 AND2X2_1/A AND2X2_1/B gnd AND2X2_1/Y vdd AND2X2
XINVX1_420 MUX2X1_48/Y gnd INVX1_420/Y vdd INVX1
XINVX1_431 NOR2X1_93/A gnd INVX1_431/Y vdd INVX1
XINVX1_442 INVX1_442/A gnd INVX1_442/Y vdd INVX1
XINVX1_453 INVX2_83/A gnd INVX1_453/Y vdd INVX1
XINVX1_475 BUFX2_50/A gnd INVX1_475/Y vdd INVX1
XINVX1_486 NOR3X1_66/B gnd INVX1_486/Y vdd INVX1
XINVX1_464 OR2X2_53/B gnd INVX1_464/Y vdd INVX1
XINVX1_497 XOR2X1_1/A gnd INVX1_497/Y vdd INVX1
XFILL_2_1 gnd vdd FILL
XFILL_44_1 gnd vdd FILL
XFILL_36_1_1 gnd vdd FILL
XNAND3X1_39 BUFX4_72/Y NAND3X1_39/B NAND3X1_39/C gnd NAND3X1_39/Y vdd NAND3X1
XNAND3X1_17 BUFX4_74/Y NAND3X1_17/B NAND3X1_17/C gnd NAND3X1_17/Y vdd NAND3X1
XNAND3X1_28 NAND3X1_28/A BUFX4_110/Y BUFX4_138/Y gnd NAND3X1_29/B vdd NAND3X1
XNOR2X1_28 INVX2_7/Y XNOR2X1_9/A gnd NOR2X1_28/Y vdd NOR2X1
XNOR2X1_17 OR2X2_6/B OR2X2_6/A gnd NOR2X1_17/Y vdd NOR2X1
XNOR2X1_39 NOR2X1_39/A NOR2X1_39/B gnd NOR2X1_39/Y vdd NOR2X1
XFILL_2_1_1 gnd vdd FILL
XFILL_27_1_1 gnd vdd FILL
XFILL_10_0_1 gnd vdd FILL
XMUX2X1_24 MUX2X1_21/B MUX2X1_24/B INVX8_8/A gnd MUX2X1_25/B vdd MUX2X1
XMUX2X1_35 MUX2X1_35/A MUX2X1_35/B INVX8_8/A gnd INVX1_396/A vdd MUX2X1
XFILL_18_1_1 gnd vdd FILL
XMUX2X1_13 MUX2X1_13/A INVX1_685/A INVX4_4/A gnd MUX2X1_13/Y vdd MUX2X1
XNOR2X1_118 INVX2_41/A MUX2X1_37/A gnd OAI22X1_8/D vdd NOR2X1
XNOR2X1_107 OAI22X1_31/B OAI22X1_31/A gnd OR2X2_32/B vdd NOR2X1
XMUX2X1_46 INVX2_30/A MUX2X1_46/B INVX8_8/A gnd MUX2X1_47/A vdd MUX2X1
XNOR2X1_129 NOR2X1_6/A NOR2X1_131/A gnd NOR2X1_129/Y vdd NOR2X1
XINVX1_261 INVX1_261/A gnd INVX1_261/Y vdd INVX1
XINVX1_250 INVX1_689/A gnd INVX1_250/Y vdd INVX1
XINVX1_272 INVX1_272/A gnd INVX1_272/Y vdd INVX1
XINVX1_294 INVX1_294/A gnd INVX1_294/Y vdd INVX1
XINVX1_283 INVX1_283/A gnd INVX1_283/Y vdd INVX1
XNAND2X1_608 INVX2_5/A BUFX4_268/Y gnd OAI21X1_785/C vdd NAND2X1
XNAND2X1_619 INVX1_258/A BUFX4_268/Y gnd NAND2X1_619/Y vdd NAND2X1
XNAND2X1_50 BUFX4_28/Y NAND2X1_50/B gnd OAI21X1_50/C vdd NAND2X1
XNAND2X1_61 BUFX4_32/Y NAND2X1_61/B gnd OAI21X1_61/C vdd NAND2X1
XNAND2X1_83 INVX2_14/A BUFX4_157/Y gnd NAND2X1_83/Y vdd NAND2X1
XNAND2X1_94 INVX1_285/A BUFX4_159/Y gnd NAND2X1_94/Y vdd NAND2X1
XNAND2X1_72 INVX1_243/A BUFX4_158/Y gnd OAI21X1_70/C vdd NAND2X1
XAOI21X1_210 INVX2_65/A AOI21X1_210/B AOI21X1_210/C gnd AOI21X1_210/Y vdd AOI21X1
XAOI21X1_221 INVX1_490/A NOR3X1_67/Y BUFX2_69/A gnd OAI21X1_866/B vdd AOI21X1
XAOI21X1_243 AND2X2_83/Y NAND2X1_977/Y OAI21X1_918/Y gnd AOI21X1_243/Y vdd AOI21X1
XAOI21X1_232 INVX1_669/Y INVX1_460/A NOR2X1_423/Y gnd NAND3X1_331/B vdd AOI21X1
XAOI21X1_254 NOR2X1_424/Y OAI21X1_934/Y AOI21X1_254/C gnd OAI21X1_937/C vdd AOI21X1
XAOI21X1_265 OAI22X1_58/C AOI21X1_265/B NOR2X1_482/Y gnd AOI21X1_265/Y vdd AOI21X1
XAOI22X1_81 AOI22X1_81/A AOI22X1_81/B AOI22X1_81/C AOI22X1_81/D gnd AOI21X1_74/A vdd
+ AOI22X1
XAOI22X1_92 INVX8_11/Y AOI22X1_92/B AOI22X1_92/C AOI22X1_92/D gnd AOI22X1_92/Y vdd
+ AOI22X1
XAOI22X1_70 OAI22X1_36/B AOI22X1_70/B AOI22X1_70/C AOI22X1_70/D gnd AOI22X1_70/Y vdd
+ AOI22X1
XNAND3X1_214 INVX1_528/Y BUFX4_209/Y BUFX4_34/Y gnd NAND3X1_214/Y vdd NAND3X1
XNAND3X1_203 BUFX4_220/Y NAND3X1_203/B NAND3X1_203/C gnd NAND2X1_729/B vdd NAND3X1
XNAND3X1_236 INVX1_550/Y BUFX4_207/Y BUFX4_35/Y gnd NAND3X1_236/Y vdd NAND3X1
XNAND3X1_225 BUFX4_219/Y NAND3X1_224/Y NAND3X1_225/C gnd NAND2X1_762/B vdd NAND3X1
XNAND3X1_247 BUFX4_222/Y NAND3X1_246/Y NAND3X1_247/C gnd NAND2X1_795/B vdd NAND3X1
XNAND3X1_269 BUFX4_120/Y NAND3X1_269/B NAND3X1_269/C gnd NAND2X1_833/B vdd NAND3X1
XNAND3X1_258 BUFX4_99/Y NOR2X1_407/Y AOI21X1_227/Y gnd BUFX4_98/A vdd NAND3X1
XDFFPOSX1_302 INVX2_48/A CLKBUF1_17/Y NOR3X1_7/Y gnd vdd DFFPOSX1
XDFFPOSX1_313 INVX2_9/A CLKBUF1_25/Y NOR2X1_418/Y gnd vdd DFFPOSX1
XDFFPOSX1_346 OR2X2_63/A CLKBUF1_4/Y OAI21X1_3/Y gnd vdd DFFPOSX1
XDFFPOSX1_324 INVX1_273/A CLKBUF1_56/Y OAI21X1_892/Y gnd vdd DFFPOSX1
XDFFPOSX1_335 NAND2X1_927/B CLKBUF1_13/Y INVX1_643/A gnd vdd DFFPOSX1
XDFFPOSX1_368 INVX1_669/A CLKBUF1_4/Y OAI21X1_25/Y gnd vdd DFFPOSX1
XDFFPOSX1_357 MUX2X1_6/B CLKBUF1_48/Y OAI21X1_14/Y gnd vdd DFFPOSX1
XDFFPOSX1_379 OR2X2_62/B CLKBUF1_62/Y OAI21X1_36/Y gnd vdd DFFPOSX1
XNAND2X1_427 BUFX4_215/Y NAND2X1_427/B gnd NAND2X1_427/Y vdd NAND2X1
XNAND2X1_405 INVX8_4/A NAND2X1_454/B gnd NAND2X1_405/Y vdd NAND2X1
XNAND2X1_416 BUFX4_227/Y NAND2X1_416/B gnd NAND2X1_416/Y vdd NAND2X1
XNAND2X1_438 BUFX4_216/Y NAND2X1_438/B gnd NAND2X1_438/Y vdd NAND2X1
XNAND2X1_449 AOI22X1_89/C AOI22X1_89/D gnd INVX2_57/A vdd NAND2X1
XNOR2X1_460 INVX2_51/A OR2X2_66/A gnd NOR2X1_460/Y vdd NOR2X1
XNOR2X1_471 NOR3X1_78/C NOR2X1_471/B gnd NOR2X1_471/Y vdd NOR2X1
XNOR2X1_482 INVX2_91/Y OAI22X1_58/C gnd NOR2X1_482/Y vdd NOR2X1
XOAI21X1_900 INVX8_14/Y AOI21X1_231/Y AOI22X1_124/Y gnd OAI21X1_900/Y vdd OAI21X1
XOAI21X1_933 INVX1_696/Y INVX2_86/A AND2X2_91/A gnd AOI21X1_251/C vdd OAI21X1
XOAI21X1_922 NOR2X1_422/B AND2X2_81/A NAND2X1_970/A gnd INVX1_705/A vdd OAI21X1
XOAI21X1_911 MUX2X1_7/B INVX1_692/Y NOR2X1_439/Y gnd AND2X2_88/A vdd OAI21X1
XOAI21X1_944 AOI21X1_259/A INVX4_12/Y NAND3X1_354/Y gnd NOR2X1_475/B vdd OAI21X1
XOAI21X1_955 INVX4_14/Y INVX1_719/Y OAI21X1_955/C gnd OAI21X1_955/Y vdd OAI21X1
XOAI21X1_966 INVX8_17/Y INVX8_15/Y OAI21X1_966/C gnd OAI21X1_967/C vdd OAI21X1
XOAI21X1_999 INVX4_13/Y INVX8_16/Y data_memory_interface_data[29] gnd OAI21X1_999/Y
+ vdd OAI21X1
XOAI21X1_977 INVX1_734/Y OAI21X1_992/B OAI21X1_977/C gnd AOI21X1_257/B vdd OAI21X1
XOAI21X1_988 INVX1_738/Y OAI21X1_992/B OAI21X1_987/Y gnd OAI21X1_988/Y vdd OAI21X1
XINVX2_30 INVX2_30/A gnd INVX2_30/Y vdd INVX2
XINVX2_52 INVX2_52/A gnd INVX2_52/Y vdd INVX2
XFILL_7_0_1 gnd vdd FILL
XINVX2_63 INVX2_63/A gnd INVX2_63/Y vdd INVX2
XINVX2_41 INVX2_41/A gnd INVX2_41/Y vdd INVX2
XINVX2_85 INVX2_85/A gnd INVX2_85/Y vdd INVX2
XNAND2X1_961 AND2X2_95/A AND2X2_95/B gnd NAND2X1_961/Y vdd NAND2X1
XNAND2X1_983 AND2X2_93/B NOR2X1_455/Y gnd NAND2X1_983/Y vdd NAND2X1
XNAND2X1_972 MUX2X1_1/B INVX2_86/A gnd AOI22X1_134/A vdd NAND2X1
XNAND2X1_950 MUX2X1_7/B OR2X2_58/B gnd AOI22X1_130/B vdd NAND2X1
XINVX2_74 INVX2_74/A gnd INVX2_74/Y vdd INVX2
XNAND2X1_994 NAND3X1_1/B AND2X2_100/A gnd NOR3X1_80/A vdd NAND2X1
XOAI21X1_15 INVX1_15/Y BUFX4_19/Y OAI21X1_15/C gnd OAI21X1_15/Y vdd OAI21X1
XOAI21X1_26 INVX1_26/Y BUFX4_17/Y OAI21X1_26/C gnd OAI21X1_26/Y vdd OAI21X1
XOAI21X1_59 INVX1_59/Y BUFX4_26/Y OAI21X1_59/C gnd OAI21X1_59/Y vdd OAI21X1
XOAI21X1_37 INVX1_37/Y BUFX4_28/Y OAI21X1_37/C gnd OAI21X1_37/Y vdd OAI21X1
XOAI21X1_48 INVX1_48/Y BUFX4_25/Y NAND2X1_48/Y gnd OAI21X1_48/Y vdd OAI21X1
XFILL_35_7_0 gnd vdd FILL
XOAI21X1_229 AND2X2_11/Y AND2X2_12/Y INVX1_230/A gnd OAI21X1_230/B vdd OAI21X1
XOAI21X1_218 BUFX4_144/Y INVX1_216/Y AOI22X1_33/Y gnd OAI21X1_218/Y vdd OAI21X1
XOAI21X1_207 BUFX4_145/Y INVX1_205/Y AOI22X1_22/Y gnd OAI21X1_207/Y vdd OAI21X1
XAND2X2_18 AND2X2_14/Y AND2X2_15/Y gnd AND2X2_18/Y vdd AND2X2
XAND2X2_29 AND2X2_29/A BUFX4_85/Y gnd AND2X2_29/Y vdd AND2X2
XDFFPOSX1_121 DFFPOSX1_9/D CLKBUF1_30/Y INVX2_5/A gnd vdd DFFPOSX1
XDFFPOSX1_110 NAND3X1_1/B CLKBUF1_3/Y AND2X2_1/B gnd vdd DFFPOSX1
XDFFPOSX1_132 DFFPOSX1_20/D CLKBUF1_12/Y INVX2_11/A gnd vdd DFFPOSX1
XDFFPOSX1_143 DFFPOSX1_31/D CLKBUF1_49/Y INVX1_276/A gnd vdd DFFPOSX1
XDFFPOSX1_154 OR2X2_50/A CLKBUF1_9/Y INVX2_2/A gnd vdd DFFPOSX1
XDFFPOSX1_165 BUFX2_8/A CLKBUF1_26/Y XNOR2X1_15/Y gnd vdd DFFPOSX1
XDFFPOSX1_176 BUFX2_19/A CLKBUF1_35/Y XNOR2X1_39/Y gnd vdd DFFPOSX1
XDFFPOSX1_187 BUFX2_30/A CLKBUF1_5/Y XNOR2X1_47/Y gnd vdd DFFPOSX1
XNAND2X1_202 INVX4_4/A AOI22X1_65/A gnd NAND2X1_202/Y vdd NAND2X1
XDFFPOSX1_198 INVX1_726/A CLKBUF1_16/Y INVX1_444/A gnd vdd DFFPOSX1
XNAND2X1_224 INVX2_34/A NOR2X1_94/B gnd OAI22X1_39/B vdd NAND2X1
XNAND2X1_235 INVX2_31/Y MUX2X1_44/B gnd INVX1_411/A vdd NAND2X1
XNAND2X1_213 INVX4_4/A AOI22X1_58/A gnd OAI21X1_294/C vdd NAND2X1
XNAND2X1_268 BUFX4_213/Y MUX2X1_12/Y gnd AOI22X1_73/C vdd NAND2X1
XNAND2X1_257 INVX2_43/Y MUX2X1_8/Y gnd AOI22X1_71/D vdd NAND2X1
XNAND2X1_246 INVX2_39/Y MUX2X1_4/Y gnd AOI22X1_70/D vdd NAND2X1
XNAND2X1_279 INVX1_342/Y MUX2X1_15/Y gnd AOI21X1_98/A vdd NAND2X1
XFILL_26_7_0 gnd vdd FILL
XFILL_1_7_0 gnd vdd FILL
XNOR2X1_290 OAI22X1_34/Y NOR2X1_290/B gnd NOR2X1_290/Y vdd NOR2X1
XOAI21X1_730 NOR2X1_314/B BUFX4_56/Y BUFX4_129/Y gnd OAI21X1_730/Y vdd OAI21X1
XOAI21X1_741 NOR2X1_355/B NOR2X1_354/Y INVX1_422/Y gnd OAI21X1_741/Y vdd OAI21X1
XOAI21X1_785 BUFX4_177/Y INVX1_438/Y OAI21X1_785/C gnd OAI21X1_785/Y vdd OAI21X1
XOAI21X1_774 NOR2X1_370/B NOR2X1_93/B INVX2_26/A gnd NAND3X1_175/C vdd OAI21X1
XOAI21X1_752 INVX2_22/A NOR2X1_366/B NOR2X1_363/Y gnd NAND3X1_169/B vdd OAI21X1
XOAI21X1_763 NOR2X1_357/B INVX1_429/A OAI21X1_763/C gnd OAI21X1_763/Y vdd OAI21X1
XOAI21X1_796 BUFX4_177/Y INVX1_449/Y NAND2X1_619/Y gnd OAI21X1_796/Y vdd OAI21X1
XNAND2X1_780 NAND2X1_780/A NAND2X1_780/B gnd NAND2X1_24/B vdd NAND2X1
XNAND2X1_791 INVX1_557/Y BUFX4_205/Y gnd NAND3X1_245/C vdd NAND2X1
XFILL_17_7_0 gnd vdd FILL
XCLKBUF1_27 BUFX4_5/Y gnd CLKBUF1_27/Y vdd CLKBUF1
XCLKBUF1_16 BUFX4_2/Y gnd CLKBUF1_16/Y vdd CLKBUF1
XCLKBUF1_38 BUFX4_2/Y gnd CLKBUF1_38/Y vdd CLKBUF1
XCLKBUF1_49 BUFX4_1/Y gnd CLKBUF1_49/Y vdd CLKBUF1
XBUFX4_70 BUFX4_69/A gnd BUFX4_70/Y vdd BUFX4
XBUFX4_92 BUFX4_93/A gnd BUFX4_92/Y vdd BUFX4
XBUFX4_81 INVX8_9/Y gnd BUFX4_81/Y vdd BUFX4
XOR2X2_40 OR2X2_40/A OR2X2_40/B gnd OR2X2_40/Y vdd OR2X2
XOR2X2_51 OR2X2_49/A BUFX2_91/A gnd OR2X2_51/Y vdd OR2X2
XOR2X2_62 OR2X2_62/A OR2X2_62/B gnd OR2X2_62/Y vdd OR2X2
XXNOR2X1_2 XOR2X1_1/A INVX2_76/A gnd XNOR2X1_2/Y vdd XNOR2X1
XFILL_41_5_0 gnd vdd FILL
XINVX1_2 gnd gnd INVX1_2/Y vdd INVX1
XOAI21X1_582 INVX2_64/Y NOR2X1_294/Y AOI21X1_125/Y gnd OAI21X1_582/Y vdd OAI21X1
XOAI21X1_560 OAI22X1_8/A INVX8_12/Y AOI22X1_97/Y gnd OAI21X1_560/Y vdd OAI21X1
XOAI21X1_593 OAI22X1_7/Y OAI21X1_593/B OAI21X1_593/C gnd OAI21X1_593/Y vdd OAI21X1
XOAI21X1_571 NOR2X1_281/B NOR2X1_281/A OAI21X1_593/B gnd AND2X2_46/A vdd OAI21X1
XINVX1_602 INVX1_529/A gnd INVX1_602/Y vdd INVX1
XINVX1_624 INVX1_551/A gnd INVX1_624/Y vdd INVX1
XINVX1_613 INVX1_613/A gnd INVX1_613/Y vdd INVX1
XINVX1_635 INVX1_635/A gnd INVX1_635/Y vdd INVX1
XINVX1_679 MUX2X1_6/B gnd INVX1_679/Y vdd INVX1
XINVX1_668 INVX1_668/A gnd INVX1_668/Y vdd INVX1
XINVX1_646 BUFX2_90/A gnd INVX1_646/Y vdd INVX1
XINVX1_657 INVX1_495/A gnd INVX1_657/Y vdd INVX1
XFILL_39_4 gnd vdd FILL
XFILL_32_5_0 gnd vdd FILL
XFILL_23_5_0 gnd vdd FILL
XFILL_6_6_0 gnd vdd FILL
XBUFX4_207 BUFX4_210/A gnd BUFX4_207/Y vdd BUFX4
XBUFX4_218 BUFX4_222/A gnd BUFX4_218/Y vdd BUFX4
XBUFX4_229 INVX8_5/Y gnd BUFX4_229/Y vdd BUFX4
XFILL_14_5_0 gnd vdd FILL
XOAI21X1_390 INVX8_4/A OAI21X1_390/B NAND2X1_374/Y gnd INVX1_365/A vdd OAI21X1
XINVX1_410 INVX1_410/A gnd INVX1_410/Y vdd INVX1
XAND2X2_2 AND2X2_2/A AND2X2_2/B gnd BUFX4_46/A vdd AND2X2
XINVX1_421 INVX1_421/A gnd INVX1_421/Y vdd INVX1
XINVX1_432 INVX1_432/A gnd INVX1_432/Y vdd INVX1
XINVX1_443 INVX1_443/A gnd INVX1_443/Y vdd INVX1
XINVX1_476 INVX1_476/A gnd INVX1_476/Y vdd INVX1
XINVX1_487 INVX1_487/A gnd NOR3X1_67/B vdd INVX1
XINVX1_454 INVX1_454/A gnd INVX1_454/Y vdd INVX1
XINVX1_465 INVX2_80/A gnd INVX1_465/Y vdd INVX1
XINVX1_498 XOR2X1_2/A gnd INVX1_498/Y vdd INVX1
XFILL_2_2 gnd vdd FILL
XFILL_37_1 gnd vdd FILL
XNAND3X1_18 NAND3X1_18/A BUFX4_110/Y BUFX4_138/Y gnd NAND3X1_18/Y vdd NAND3X1
XNAND3X1_29 BUFX4_75/Y NAND3X1_29/B NAND3X1_29/C gnd NAND3X1_29/Y vdd NAND3X1
XNOR2X1_18 NOR2X1_18/A OR2X2_5/B gnd NOR2X1_18/Y vdd NOR2X1
XNOR2X1_29 NOR2X1_29/A NOR2X1_29/B gnd NOR2X1_29/Y vdd NOR2X1
XMUX2X1_25 MUX2X1_25/A MUX2X1_25/B INVX8_5/A gnd AND2X2_32/A vdd MUX2X1
XMUX2X1_36 MUX2X1_36/A MUX2X1_36/B BUFX4_229/Y gnd MUX2X1_36/Y vdd MUX2X1
XMUX2X1_14 MUX2X1_14/A OR2X2_64/A INVX4_4/A gnd MUX2X1_14/Y vdd MUX2X1
XNOR2X1_119 OAI22X1_7/Y OAI22X1_8/Y gnd NAND3X1_93/C vdd NOR2X1
XNOR2X1_108 NOR2X1_108/A NOR2X1_108/B gnd NOR2X1_108/Y vdd NOR2X1
XMUX2X1_47 MUX2X1_47/A MUX2X1_47/B MUX2X1_47/S gnd MUX2X1_47/Y vdd MUX2X1
XINVX1_240 INVX1_240/A gnd INVX1_240/Y vdd INVX1
XINVX1_251 INVX1_251/A gnd INVX1_251/Y vdd INVX1
XINVX1_262 NOR2X1_28/Y gnd INVX1_262/Y vdd INVX1
XINVX1_273 INVX1_273/A gnd OR2X2_13/B vdd INVX1
XINVX1_295 INVX1_295/A gnd INVX1_295/Y vdd INVX1
XINVX1_284 NOR2X1_55/Y gnd INVX1_284/Y vdd INVX1
XNAND2X1_609 INVX2_7/A BUFX4_264/Y gnd NAND2X1_609/Y vdd NAND2X1
XNAND2X1_51 BUFX4_31/Y NAND2X1_51/B gnd NAND2X1_51/Y vdd NAND2X1
XNAND2X1_40 BUFX4_27/Y NAND2X1_40/B gnd NAND2X1_40/Y vdd NAND2X1
XNAND2X1_73 INVX1_245/A BUFX4_159/Y gnd NAND2X1_73/Y vdd NAND2X1
XNAND2X1_84 INVX1_261/A BUFX4_161/Y gnd NAND2X1_84/Y vdd NAND2X1
XNAND2X1_62 BUFX4_25/Y NAND2X1_62/B gnd OAI21X1_62/C vdd NAND2X1
XNAND2X1_95 INVX1_288/A BUFX4_156/Y gnd NAND2X1_95/Y vdd NAND2X1
XFILL_37_4_0 gnd vdd FILL
XAOI21X1_200 INVX1_423/A AOI21X1_200/B INVX1_424/A gnd NOR2X1_357/B vdd AOI21X1
XFILL_20_3_0 gnd vdd FILL
XAOI21X1_211 NOR2X1_367/Y INVX2_71/Y INVX1_428/Y gnd OAI21X1_773/C vdd AOI21X1
XAOI21X1_233 INVX1_681/Y INVX1_444/A NOR2X1_431/Y gnd NAND3X1_334/B vdd AOI21X1
XAOI21X1_222 INVX2_74/A INVX1_498/Y INVX1_499/Y gnd AOI21X1_222/Y vdd AOI21X1
XAOI21X1_255 INVX2_49/A INVX1_713/Y INVX1_714/Y gnd AOI21X1_255/Y vdd AOI21X1
XAOI21X1_244 AOI22X1_127/Y OAI21X1_919/Y AOI21X1_244/C gnd NOR2X1_452/B vdd AOI21X1
XAOI21X1_266 OAI22X1_58/C AOI21X1_266/B NOR2X1_482/Y gnd BUFX4_65/A vdd AOI21X1
XAOI22X1_60 AOI22X1_60/A AND2X2_12/A BUFX4_146/Y INVX2_82/A gnd INVX1_275/A vdd AOI22X1
XAOI22X1_71 AOI22X1_71/A AOI22X1_71/B OAI22X1_25/C AOI22X1_71/D gnd AOI22X1_71/Y vdd
+ AOI22X1
XAOI22X1_82 AOI22X1_82/A BUFX4_189/Y OR2X2_24/Y INVX1_378/Y gnd AOI22X1_82/Y vdd AOI22X1
XAOI22X1_93 AND2X2_26/A INVX2_56/Y AND2X2_42/A AOI22X1_94/D gnd AOI22X1_93/Y vdd AOI22X1
XFILL_3_4_0 gnd vdd FILL
XFILL_28_4_0 gnd vdd FILL
XNAND3X1_204 INVX1_518/Y BUFX4_209/Y BUFX4_34/Y gnd NAND3X1_204/Y vdd NAND3X1
XNAND3X1_237 BUFX4_219/Y NAND3X1_236/Y NAND3X1_237/C gnd NAND2X1_780/B vdd NAND3X1
XNAND3X1_215 BUFX4_220/Y NAND3X1_214/Y NAND3X1_215/C gnd NAND2X1_747/B vdd NAND3X1
XNAND3X1_226 INVX1_540/Y BUFX4_208/Y BUFX4_36/Y gnd NAND3X1_227/B vdd NAND3X1
XNAND3X1_248 INVX1_562/Y BUFX4_210/Y BUFX4_37/Y gnd NAND3X1_248/Y vdd NAND3X1
XFILL_11_3_0 gnd vdd FILL
XNAND3X1_259 NAND2X1_817/Y NAND2X1_818/Y NAND2X1_819/Y gnd NOR2X1_408/A vdd NAND3X1
XFILL_19_4_0 gnd vdd FILL
XDFFPOSX1_303 INVX1_230/A CLKBUF1_56/Y OAI22X1_49/Y gnd vdd DFFPOSX1
XDFFPOSX1_347 OR2X2_62/A CLKBUF1_58/Y OAI21X1_4/Y gnd vdd DFFPOSX1
XDFFPOSX1_336 NAND2X1_927/A CLKBUF1_13/Y INVX2_79/A gnd vdd DFFPOSX1
XDFFPOSX1_325 INVX1_274/A CLKBUF1_1/Y OAI21X1_893/Y gnd vdd DFFPOSX1
XDFFPOSX1_314 INVX2_10/A CLKBUF1_49/Y NAND3X1_327/Y gnd vdd DFFPOSX1
XDFFPOSX1_358 MUX2X1_4/B CLKBUF1_53/Y OAI21X1_15/Y gnd vdd DFFPOSX1
XDFFPOSX1_369 INVX1_306/A CLKBUF1_53/Y OAI21X1_26/Y gnd vdd DFFPOSX1
XNAND2X1_417 BUFX4_215/Y MUX2X1_33/A gnd NAND2X1_417/Y vdd NAND2X1
XNAND2X1_406 BUFX4_78/Y NAND2X1_406/B gnd NAND3X1_110/A vdd NAND2X1
XNAND2X1_428 BUFX4_81/Y OAI21X1_558/B gnd OAI22X1_14/C vdd NAND2X1
XNAND2X1_439 MUX2X1_49/S INVX1_364/Y gnd OAI21X1_472/C vdd NAND2X1
XNOR2X1_450 INVX1_458/A INVX1_700/Y gnd NOR2X1_450/Y vdd NOR2X1
XNOR2X1_461 OR2X2_68/A OR2X2_68/B gnd NOR2X1_461/Y vdd NOR2X1
XNOR2X1_483 INVX8_15/A INVX8_17/Y gnd AND2X2_101/B vdd NOR2X1
XNOR2X1_472 INVX2_87/A INVX4_12/Y gnd INVX8_16/A vdd NOR2X1
XOAI21X1_934 AOI21X1_251/Y NAND2X1_989/Y AOI21X1_252/Y gnd OAI21X1_934/Y vdd OAI21X1
XOAI21X1_912 NOR2X1_429/Y AND2X2_86/A OAI21X1_912/C gnd INVX1_695/A vdd OAI21X1
XOAI21X1_901 INVX8_14/Y AOI21X1_231/Y AOI22X1_125/Y gnd OAI21X1_901/Y vdd OAI21X1
XOAI21X1_923 AND2X2_92/Y NAND2X1_981/Y INVX1_705/Y gnd NOR2X1_454/A vdd OAI21X1
XOAI21X1_945 INVX4_13/Y INVX8_16/Y NOR2X1_475/Y gnd BUFX2_35/A vdd OAI21X1
XOAI21X1_956 INVX8_17/Y INVX8_15/Y BUFX2_79/A gnd OAI21X1_956/Y vdd OAI21X1
XOAI21X1_967 INVX4_14/Y INVX1_725/Y OAI21X1_967/C gnd OAI21X1_967/Y vdd OAI21X1
XOAI21X1_978 INVX8_17/Y INVX8_15/Y NOR3X1_73/B gnd OAI21X1_994/B vdd OAI21X1
XOAI21X1_989 INVX1_738/Y OAI21X1_993/B OAI21X1_989/C gnd OAI21X1_989/Y vdd OAI21X1
XINVX2_20 INVX2_20/A gnd INVX2_20/Y vdd INVX2
XINVX2_42 INVX2_42/A gnd INVX2_42/Y vdd INVX2
XINVX2_53 INVX2_53/A gnd INVX2_53/Y vdd INVX2
XINVX2_31 INVX2_31/A gnd INVX2_31/Y vdd INVX2
XNAND2X1_940 INVX1_672/A INVX1_457/A gnd NAND2X1_940/Y vdd NAND2X1
XINVX2_75 INVX2_75/A gnd INVX2_75/Y vdd INVX2
XINVX2_64 INVX2_64/A gnd INVX2_64/Y vdd INVX2
XNAND2X1_962 OR2X2_60/B INVX2_85/Y gnd NAND2X1_962/Y vdd NAND2X1
XNAND2X1_973 INVX1_696/Y INVX2_86/Y gnd AOI22X1_134/B vdd NAND2X1
XINVX2_86 INVX2_86/A gnd INVX2_86/Y vdd INVX2
XNAND2X1_951 OR2X2_59/A OR2X2_59/B gnd NAND2X1_951/Y vdd NAND2X1
XNAND2X1_984 NAND2X1_962/Y NOR2X1_435/Y gnd NAND2X1_984/Y vdd NAND2X1
XNAND2X1_995 INVX2_89/Y NOR2X1_471/Y gnd NAND3X1_349/A vdd NAND2X1
XFILL_43_2_0 gnd vdd FILL
XOAI21X1_16 INVX1_16/Y BUFX4_23/Y OAI21X1_16/C gnd OAI21X1_16/Y vdd OAI21X1
XOAI21X1_27 INVX1_27/Y BUFX4_19/Y OAI21X1_27/C gnd OAI21X1_27/Y vdd OAI21X1
XOAI21X1_38 INVX1_38/Y BUFX4_29/Y OAI21X1_38/C gnd OAI21X1_38/Y vdd OAI21X1
XOAI21X1_49 INVX1_49/Y BUFX4_29/Y OAI21X1_49/C gnd OAI21X1_49/Y vdd OAI21X1
XFILL_35_7_1 gnd vdd FILL
XFILL_34_2_0 gnd vdd FILL
XOAI21X1_208 BUFX4_141/Y INVX1_206/Y AOI22X1_23/Y gnd OAI21X1_208/Y vdd OAI21X1
XOAI21X1_219 BUFX4_142/Y INVX1_217/Y AOI22X1_34/Y gnd OAI21X1_219/Y vdd OAI21X1
XAND2X2_19 INVX1_297/Y AND2X2_19/B gnd AND2X2_19/Y vdd AND2X2
XDFFPOSX1_100 INVX1_213/A CLKBUF1_50/Y OAI21X1_141/C gnd vdd DFFPOSX1
XDFFPOSX1_111 INVX1_715/A CLKBUF1_61/Y AND2X2_1/A gnd vdd DFFPOSX1
XDFFPOSX1_133 DFFPOSX1_21/D CLKBUF1_2/Y INVX1_258/A gnd vdd DFFPOSX1
XDFFPOSX1_144 DFFPOSX1_32/D CLKBUF1_32/Y INVX1_278/A gnd vdd DFFPOSX1
XDFFPOSX1_122 DFFPOSX1_10/D CLKBUF1_49/Y INVX2_6/A gnd vdd DFFPOSX1
XDFFPOSX1_155 INVX1_502/A CLKBUF1_9/Y XOR2X1_2/A gnd vdd DFFPOSX1
XDFFPOSX1_177 BUFX2_20/A CLKBUF1_54/Y XOR2X1_4/Y gnd vdd DFFPOSX1
XDFFPOSX1_166 BUFX2_9/A CLKBUF1_33/Y XNOR2X1_18/Y gnd vdd DFFPOSX1
XDFFPOSX1_188 BUFX2_31/A CLKBUF1_6/Y NOR2X1_67/Y gnd vdd DFFPOSX1
XNAND2X1_225 INVX2_34/Y MUX2X1_1/Y gnd AOI21X1_153/A vdd NAND2X1
XNAND2X1_214 INVX2_31/Y INVX1_321/Y gnd INVX1_410/A vdd NAND2X1
XNAND2X1_203 INVX4_4/A AOI22X1_66/A gnd NAND2X1_203/Y vdd NAND2X1
XDFFPOSX1_199 INVX1_727/A CLKBUF1_16/Y INVX2_84/A gnd vdd DFFPOSX1
XNAND2X1_269 INVX4_4/A INVX1_351/A gnd OAI21X1_316/C vdd NAND2X1
XNAND2X1_258 INVX4_4/A MUX2X1_9/A gnd NAND2X1_258/Y vdd NAND2X1
XNAND2X1_247 INVX4_4/A MUX2X1_5/A gnd OAI21X1_309/C vdd NAND2X1
XNAND2X1_236 INVX2_37/A MUX2X1_42/A gnd INVX2_68/A vdd NAND2X1
XFILL_0_2_0 gnd vdd FILL
XFILL_1_7_1 gnd vdd FILL
XFILL_25_2_0 gnd vdd FILL
XFILL_26_7_1 gnd vdd FILL
XNOR2X1_291 INVX2_38/Y MUX2X1_39/A gnd OAI22X1_38/A vdd NOR2X1
XNOR2X1_280 BUFX4_53/Y OR2X2_30/B gnd INVX4_9/A vdd NOR2X1
XOAI21X1_731 NOR2X1_265/Y BUFX4_129/Y INVX2_65/A gnd NOR2X1_348/B vdd OAI21X1
XOAI21X1_720 INVX1_307/A INVX4_3/A INVX8_12/A gnd NAND3X1_162/B vdd OAI21X1
XOAI21X1_742 OAI21X1_722/C NOR2X1_356/B AOI21X1_199/Y gnd INVX1_424/A vdd OAI21X1
XOAI21X1_753 NOR2X1_357/B INVX2_22/Y NOR2X1_365/Y gnd OAI21X1_753/Y vdd OAI21X1
XOAI21X1_775 AND2X2_70/A AND2X2_70/B INVX1_381/Y gnd OAI21X1_775/Y vdd OAI21X1
XOAI21X1_764 INVX2_28/A OAI21X1_763/Y NOR2X1_370/Y gnd NAND3X1_173/A vdd OAI21X1
XOAI21X1_786 BUFX4_180/Y INVX1_439/Y NAND2X1_609/Y gnd OAI21X1_786/Y vdd OAI21X1
XOAI21X1_797 BUFX4_179/Y INVX1_450/Y NAND2X1_620/Y gnd OAI21X1_797/Y vdd OAI21X1
XFILL_8_3_0 gnd vdd FILL
XNAND2X1_770 INVX1_543/Y BUFX4_203/Y gnd NAND3X1_231/C vdd NAND2X1
XNAND2X1_781 OAI21X1_89/Y BUFX4_134/Y gnd NAND2X1_783/A vdd NAND2X1
XNAND2X1_792 NAND2X1_790/Y NAND2X1_792/B gnd NAND2X1_28/B vdd NAND2X1
XFILL_16_2_0 gnd vdd FILL
XFILL_17_7_1 gnd vdd FILL
XCLKBUF1_17 BUFX4_6/Y gnd CLKBUF1_17/Y vdd CLKBUF1
XCLKBUF1_28 BUFX4_2/Y gnd CLKBUF1_28/Y vdd CLKBUF1
XCLKBUF1_39 BUFX4_1/Y gnd CLKBUF1_39/Y vdd CLKBUF1
XBUFX4_60 BUFX4_62/A gnd BUFX4_60/Y vdd BUFX4
XBUFX4_71 BUFX4_69/A gnd BUFX4_71/Y vdd BUFX4
XBUFX4_82 INVX8_9/Y gnd BUFX4_82/Y vdd BUFX4
XBUFX4_93 BUFX4_93/A gnd BUFX4_93/Y vdd BUFX4
XOR2X2_30 OR2X2_30/A OR2X2_30/B gnd OR2X2_30/Y vdd OR2X2
XOR2X2_41 OR2X2_41/A INVX8_3/A gnd OR2X2_41/Y vdd OR2X2
XOR2X2_52 OR2X2_50/A OR2X2_52/B gnd OR2X2_52/Y vdd OR2X2
XOR2X2_63 OR2X2_63/A OR2X2_63/B gnd OR2X2_63/Y vdd OR2X2
XOR2X2_1 OR2X2_1/A OR2X2_1/B gnd OR2X2_1/Y vdd OR2X2
XXNOR2X1_3 XOR2X1_1/A INVX2_73/A gnd AND2X2_4/A vdd XNOR2X1
XFILL_41_5_1 gnd vdd FILL
XFILL_40_0_0 gnd vdd FILL
XINVX1_3 gnd gnd INVX1_3/Y vdd INVX1
XOAI21X1_550 OAI22X1_37/A AOI22X1_96/D AOI22X1_96/A gnd AOI21X1_113/C vdd OAI21X1
XOAI21X1_572 INVX2_63/Y AND2X2_46/A NOR2X1_286/Y gnd OAI21X1_572/Y vdd OAI21X1
XOAI21X1_561 INVX2_40/A MUX2X1_5/Y NOR2X1_281/B gnd OAI21X1_561/Y vdd OAI21X1
XOAI21X1_583 BUFX4_43/Y MUX2X1_4/Y OAI21X1_583/C gnd OAI21X1_612/A vdd OAI21X1
XINVX1_614 INVX1_614/A gnd INVX1_614/Y vdd INVX1
XOAI21X1_594 OAI21X1_551/A NAND3X1_93/Y OAI21X1_594/C gnd AOI21X1_180/B vdd OAI21X1
XINVX1_636 INVX1_636/A gnd INVX1_636/Y vdd INVX1
XINVX1_603 INVX1_603/A gnd INVX1_603/Y vdd INVX1
XINVX1_625 INVX1_625/A gnd INVX1_625/Y vdd INVX1
XINVX1_669 INVX1_669/A gnd INVX1_669/Y vdd INVX1
XINVX1_647 BUFX2_91/A gnd INVX1_647/Y vdd INVX1
XINVX1_658 INVX2_73/A gnd INVX1_658/Y vdd INVX1
XFILL_32_5_1 gnd vdd FILL
XFILL_31_0_0 gnd vdd FILL
XFILL_39_1_0 gnd vdd FILL
XFILL_22_0_0 gnd vdd FILL
XFILL_23_5_1 gnd vdd FILL
XFILL_6_6_1 gnd vdd FILL
XFILL_5_1_0 gnd vdd FILL
XBUFX4_219 BUFX4_222/A gnd BUFX4_219/Y vdd BUFX4
XBUFX4_208 BUFX4_210/A gnd BUFX4_208/Y vdd BUFX4
XFILL_13_0_0 gnd vdd FILL
XFILL_14_5_1 gnd vdd FILL
XOAI21X1_391 BUFX4_52/Y NOR2X1_251/B NAND2X1_375/Y gnd OAI21X1_391/Y vdd OAI21X1
XINVX1_400 INVX1_400/A gnd INVX1_400/Y vdd INVX1
XINVX1_411 INVX1_411/A gnd INVX1_411/Y vdd INVX1
XOAI21X1_380 INVX1_361/Y AND2X2_70/B NAND2X1_366/Y gnd OAI21X1_380/Y vdd OAI21X1
XAND2X2_3 AND2X2_3/A AND2X2_3/B gnd AND2X2_3/Y vdd AND2X2
XINVX1_422 INVX1_422/A gnd INVX1_422/Y vdd INVX1
XINVX1_433 INVX1_433/A gnd INVX1_433/Y vdd INVX1
XINVX1_444 INVX1_444/A gnd INVX1_444/Y vdd INVX1
XINVX1_477 BUFX2_52/A gnd INVX1_477/Y vdd INVX1
XINVX1_455 INVX2_86/A gnd INVX1_455/Y vdd INVX1
XINVX1_466 INVX1_666/A gnd INVX1_466/Y vdd INVX1
XINVX1_488 BUFX2_67/A gnd INVX1_488/Y vdd INVX1
XINVX1_499 INVX1_572/A gnd INVX1_499/Y vdd INVX1
XFILL_2_3 gnd vdd FILL
XFILL_37_2 gnd vdd FILL
XNAND3X1_19 BUFX4_72/Y NAND3X1_18/Y NAND3X1_19/C gnd NAND3X1_19/Y vdd NAND3X1
XNOR2X1_19 INVX2_4/A INVX1_228/Y gnd INVX1_229/A vdd NOR2X1
XMUX2X1_15 INVX1_251/A INVX1_689/A INVX4_4/A gnd MUX2X1_15/Y vdd MUX2X1
XMUX2X1_26 MUX2X1_26/A MUX2X1_26/B INVX8_4/A gnd MUX2X1_26/Y vdd MUX2X1
XNOR2X1_109 INVX8_8/A MUX2X1_13/Y gnd INVX2_52/A vdd NOR2X1
XMUX2X1_37 MUX2X1_37/A MUX2X1_37/B INVX8_8/A gnd MUX2X1_37/Y vdd MUX2X1
XMUX2X1_48 INVX2_50/A INVX4_3/A INVX8_8/A gnd MUX2X1_48/Y vdd MUX2X1
XINVX1_252 INVX1_252/A gnd INVX1_252/Y vdd INVX1
XINVX1_241 INVX2_85/A gnd AOI21X1_9/C vdd INVX1
XINVX1_230 INVX1_230/A gnd INVX1_230/Y vdd INVX1
XINVX1_263 INVX1_263/A gnd INVX1_263/Y vdd INVX1
XINVX1_274 INVX1_274/A gnd OR2X2_14/B vdd INVX1
XINVX1_285 INVX1_285/A gnd INVX1_285/Y vdd INVX1
XINVX1_296 INVX1_296/A gnd INVX1_296/Y vdd INVX1
XNAND2X1_30 BUFX4_20/Y NAND2X1_30/B gnd OAI21X1_30/C vdd NAND2X1
XNAND2X1_41 BUFX4_31/Y NAND2X1_41/B gnd NAND2X1_41/Y vdd NAND2X1
XNAND2X1_52 BUFX4_31/Y NAND2X1_52/B gnd OAI21X1_52/C vdd NAND2X1
XNAND2X1_74 INVX1_249/A BUFX4_157/Y gnd NAND2X1_74/Y vdd NAND2X1
XNAND2X1_63 BUFX4_30/Y NAND2X1_63/B gnd OAI21X1_63/C vdd NAND2X1
XNAND2X1_85 INVX1_264/A BUFX4_158/Y gnd NAND2X1_85/Y vdd NAND2X1
XFILL_37_4_1 gnd vdd FILL
XNAND2X1_96 NOR2X1_62/A BUFX4_156/Y gnd OAI21X1_94/C vdd NAND2X1
XAOI21X1_223 INVX2_75/Y INVX1_495/A OAI22X1_45/Y gnd AOI21X1_223/Y vdd AOI21X1
XAOI21X1_212 AOI21X1_89/A INVX1_397/Y AOI21X1_212/C gnd AOI21X1_212/Y vdd AOI21X1
XAOI21X1_201 INVX2_65/A MUX2X1_53/Y AOI21X1_201/C gnd AOI21X1_201/Y vdd AOI21X1
XAOI21X1_234 AOI21X1_234/A NOR2X1_434/Y INVX1_708/A gnd AOI21X1_234/Y vdd AOI21X1
XFILL_20_3_1 gnd vdd FILL
XAOI21X1_245 AOI21X1_245/A OAI21X1_925/Y NAND2X1_983/Y gnd OAI21X1_941/B vdd AOI21X1
XAOI21X1_267 INVX2_92/Y INVX2_93/Y AOI21X1_267/C gnd NOR2X1_485/B vdd AOI21X1
XAOI21X1_256 NOR3X1_79/A NOR3X1_80/A NOR3X1_80/C gnd INVX4_13/A vdd AOI21X1
XAOI22X1_50 MUX2X1_5/A BUFX4_235/Y BUFX4_151/Y OR2X2_57/A gnd XNOR2X1_28/A vdd AOI22X1
XAOI22X1_83 AOI22X1_83/A AOI22X1_87/A AOI22X1_83/C AOI21X1_79/Y gnd AOI22X1_83/Y vdd
+ AOI22X1
XAOI22X1_72 AOI22X1_72/A AOI22X1_72/B AND2X2_36/A AND2X2_36/B gnd AOI22X1_72/Y vdd
+ AOI22X1
XAOI22X1_61 AOI22X1_61/A BUFX4_233/Y BUFX4_148/Y INVX1_669/A gnd NOR2X1_52/B vdd AOI22X1
XAOI22X1_94 INVX1_377/A INVX2_56/Y AOI21X1_49/B AOI22X1_94/D gnd AOI22X1_94/Y vdd
+ AOI22X1
XFILL_28_4_1 gnd vdd FILL
XFILL_3_4_1 gnd vdd FILL
XNAND3X1_205 BUFX4_218/Y NAND3X1_204/Y NAND3X1_205/C gnd NAND2X1_732/B vdd NAND3X1
XNAND3X1_238 INVX1_552/Y BUFX4_207/Y BUFX4_35/Y gnd NAND3X1_238/Y vdd NAND3X1
XNAND3X1_216 INVX1_530/Y BUFX4_206/Y BUFX4_33/Y gnd NAND3X1_217/B vdd NAND3X1
XNAND3X1_227 BUFX4_221/Y NAND3X1_227/B NAND3X1_227/C gnd NAND2X1_765/B vdd NAND3X1
XNAND3X1_249 BUFX4_222/Y NAND3X1_248/Y NAND3X1_249/C gnd NAND2X1_798/B vdd NAND3X1
XFILL_11_3_1 gnd vdd FILL
XOAI22X1_1 OAI22X1_1/A OAI22X1_1/B OAI22X1_1/C OAI22X1_1/D gnd OAI22X1_1/Y vdd OAI22X1
XFILL_19_4_1 gnd vdd FILL
XDFFPOSX1_304 INVX2_5/A CLKBUF1_40/Y OAI21X1_877/Y gnd vdd DFFPOSX1
XDFFPOSX1_315 INVX2_11/A CLKBUF1_56/Y OAI21X1_883/Y gnd vdd DFFPOSX1
XDFFPOSX1_337 NOR2X1_419/A CLKBUF1_56/Y OAI22X1_6/Y gnd vdd DFFPOSX1
XDFFPOSX1_326 INVX1_276/A CLKBUF1_49/Y OAI21X1_894/Y gnd vdd DFFPOSX1
XDFFPOSX1_348 OR2X2_61/A CLKBUF1_58/Y OAI21X1_5/Y gnd vdd DFFPOSX1
XDFFPOSX1_359 MUX2X1_3/B CLKBUF1_53/Y OAI21X1_16/Y gnd vdd DFFPOSX1
XNAND2X1_407 NAND2X1_407/A NOR2X1_208/Y gnd NAND3X1_110/B vdd NAND2X1
XNAND2X1_418 INVX8_5/A OAI21X1_379/Y gnd OAI21X1_436/C vdd NAND2X1
XNAND2X1_429 INVX8_4/A OAI21X1_353/B gnd OAI21X1_451/C vdd NAND2X1
XNOR2X1_440 OR2X2_57/B INVX1_694/Y gnd NOR2X1_440/Y vdd NOR2X1
XNOR2X1_451 OR2X2_54/A INVX1_702/Y gnd NOR2X1_451/Y vdd NOR2X1
XNOR2X1_462 NOR2X1_462/A NOR2X1_462/B gnd NOR2X1_462/Y vdd NOR2X1
XNOR2X1_473 AND2X2_99/B INVX2_88/A gnd INVX8_17/A vdd NOR2X1
XNOR2X1_484 INVX1_753/Y AND2X2_101/B gnd BUFX4_69/A vdd NOR2X1
XOAI21X1_902 NAND3X1_328/Y OAI21X1_902/B INVX1_662/Y gnd BUFX4_242/A vdd OAI21X1
XOAI21X1_913 OAI21X1_913/A INVX1_710/A INVX1_695/Y gnd OAI21X1_913/Y vdd OAI21X1
XOAI21X1_924 AOI21X1_243/Y NOR2X1_462/A NOR2X1_454/Y gnd OAI21X1_925/B vdd OAI21X1
XOAI21X1_935 INVX1_668/Y INVX2_80/A AND2X2_92/A gnd OAI21X1_935/Y vdd OAI21X1
XOAI21X1_957 INVX4_14/Y INVX1_720/Y OAI21X1_956/Y gnd OAI21X1_957/Y vdd OAI21X1
XOAI21X1_946 NOR3X1_77/Y NOR3X1_78/Y NOR2X1_476/Y gnd INVX1_759/A vdd OAI21X1
XOAI21X1_968 INVX1_726/Y BUFX4_118/Y OAI21X1_968/C gnd OAI21X1_968/Y vdd OAI21X1
XOAI21X1_979 NOR3X1_79/A NAND3X1_356/Y AOI21X1_259/A gnd OAI21X1_979/Y vdd OAI21X1
XINVX2_10 INVX2_10/A gnd INVX2_10/Y vdd INVX2
XINVX2_21 INVX2_21/A gnd INVX2_21/Y vdd INVX2
XINVX2_43 INVX2_43/A gnd INVX2_43/Y vdd INVX2
XINVX2_54 INVX2_54/A gnd INVX2_54/Y vdd INVX2
XINVX2_32 INVX2_32/A gnd INVX2_32/Y vdd INVX2
XNAND2X1_930 INVX1_666/A INVX1_667/Y gnd AND2X2_81/B vdd NAND2X1
XINVX2_65 INVX2_65/A gnd INVX2_65/Y vdd INVX2
XNAND2X1_941 INVX1_672/Y INVX1_673/Y gnd NAND2X1_941/Y vdd NAND2X1
XNAND2X1_963 AOI22X1_130/Y OAI21X1_910/Y gnd NAND2X1_963/Y vdd NAND2X1
XNAND2X1_952 INVX1_681/A INVX1_682/Y gnd AND2X2_87/A vdd NAND2X1
XINVX2_87 INVX2_87/A gnd INVX2_87/Y vdd INVX2
XINVX2_76 INVX2_76/A gnd INVX2_76/Y vdd INVX2
XNAND2X1_974 MUX2X1_2/B INVX1_454/A gnd NAND2X1_974/Y vdd NAND2X1
XNAND2X1_985 AND2X2_88/B AND2X2_88/A gnd AOI21X1_248/C vdd NAND2X1
XNAND2X1_996 AND2X2_99/B INVX8_15/Y gnd NOR3X1_73/B vdd NAND2X1
XFILL_43_2_1 gnd vdd FILL
XOAI21X1_17 INVX1_17/Y BUFX4_24/Y OAI21X1_17/C gnd OAI21X1_17/Y vdd OAI21X1
XOAI21X1_28 INVX1_28/Y BUFX4_22/Y OAI21X1_28/C gnd OAI21X1_28/Y vdd OAI21X1
XOAI21X1_39 INVX1_39/Y BUFX4_32/Y OAI21X1_39/C gnd OAI21X1_39/Y vdd OAI21X1
XFILL_34_2_1 gnd vdd FILL
XFILL_12_1 gnd vdd FILL
XOAI21X1_209 BUFX4_142/Y INVX1_207/Y AOI22X1_24/Y gnd OAI21X1_209/Y vdd OAI21X1
XDFFPOSX1_101 INVX1_214/A CLKBUF1_23/Y OAI21X1_143/C gnd vdd DFFPOSX1
XDFFPOSX1_112 OR2X2_69/A CLKBUF1_60/Y INVX1_66/A gnd vdd DFFPOSX1
XDFFPOSX1_145 DFFPOSX1_33/D CLKBUF1_32/Y INVX1_279/A gnd vdd DFFPOSX1
XDFFPOSX1_134 DFFPOSX1_22/D CLKBUF1_49/Y INVX2_12/A gnd vdd DFFPOSX1
XDFFPOSX1_123 DFFPOSX1_11/D CLKBUF1_24/Y INVX2_7/A gnd vdd DFFPOSX1
XDFFPOSX1_167 BUFX2_10/A CLKBUF1_14/Y XNOR2X1_19/Y gnd vdd DFFPOSX1
XDFFPOSX1_178 BUFX2_21/A CLKBUF1_35/Y XNOR2X1_40/Y gnd vdd DFFPOSX1
XDFFPOSX1_189 BUFX2_32/A CLKBUF1_6/Y NAND2X1_192/Y gnd vdd DFFPOSX1
XDFFPOSX1_156 OR2X2_49/A CLKBUF1_39/Y INVX2_3/A gnd vdd DFFPOSX1
XNAND2X1_226 AOI21X1_153/A OAI22X1_39/B gnd AOI21X1_37/B vdd NAND2X1
XNAND2X1_215 INVX2_31/A MUX2X1_44/B gnd INVX2_69/A vdd NAND2X1
XNAND2X1_204 INVX4_4/A AOI22X1_68/A gnd NAND2X1_204/Y vdd NAND2X1
XNAND2X1_248 INVX4_4/A MUX2X1_6/A gnd OAI21X1_310/C vdd NAND2X1
XNAND2X1_237 INVX2_37/Y NOR2X1_96/B gnd NAND2X1_237/Y vdd NAND2X1
XNAND2X1_259 INVX2_44/A NOR2X1_249/B gnd AOI22X1_72/A vdd NAND2X1
XFILL_25_2_1 gnd vdd FILL
XNOR2X1_270 INVX8_3/A NOR2X1_270/B gnd NOR2X1_270/Y vdd NOR2X1
XFILL_0_2_1 gnd vdd FILL
XNOR2X1_281 NOR2X1_281/A NOR2X1_281/B gnd NOR2X1_281/Y vdd NOR2X1
XNOR2X1_292 INVX2_39/A MUX2X1_4/Y gnd NOR2X1_293/A vdd NOR2X1
XOAI21X1_732 OAI21X1_732/A AND2X2_64/B OAI21X1_750/B gnd OAI21X1_732/Y vdd OAI21X1
XOAI21X1_721 AND2X2_64/Y OAI21X1_721/B AOI21X1_190/Y gnd INVX1_91/A vdd OAI21X1
XOAI21X1_710 AND2X2_64/A AND2X2_64/B INVX8_11/Y gnd OAI21X1_721/B vdd OAI21X1
XOAI21X1_776 OAI21X1_775/Y AND2X2_73/Y MUX2X1_49/S gnd OAI21X1_776/Y vdd OAI21X1
XOAI21X1_765 INVX2_24/Y BUFX4_40/Y NAND2X1_335/Y gnd NOR2X1_372/B vdd OAI21X1
XOAI21X1_743 OAI21X1_743/A INVX1_423/Y INVX1_424/Y gnd OAI21X1_744/B vdd OAI21X1
XOAI21X1_754 NOR2X1_357/Y NOR2X1_85/B INVX2_71/A gnd NAND3X1_170/C vdd OAI21X1
XOAI21X1_787 BUFX4_181/Y INVX1_440/Y NAND2X1_610/Y gnd OAI21X1_787/Y vdd OAI21X1
XOAI21X1_798 BUFX4_178/Y INVX1_451/Y NAND2X1_621/Y gnd OAI21X1_798/Y vdd OAI21X1
XFILL_8_3_1 gnd vdd FILL
XNAND2X1_760 OAI21X1_82/Y BUFX4_134/Y gnd NAND2X1_762/A vdd NAND2X1
XNAND2X1_771 NAND2X1_769/Y NAND2X1_771/B gnd NAND2X1_21/B vdd NAND2X1
XNAND2X1_782 INVX1_551/Y BUFX4_203/Y gnd NAND3X1_239/C vdd NAND2X1
XNAND2X1_793 OAI21X1_93/Y BUFX4_131/Y gnd NAND2X1_795/A vdd NAND2X1
XFILL_16_2_1 gnd vdd FILL
XCLKBUF1_18 BUFX4_6/Y gnd CLKBUF1_18/Y vdd CLKBUF1
XCLKBUF1_29 BUFX4_2/Y gnd CLKBUF1_29/Y vdd CLKBUF1
XBUFX4_50 BUFX4_46/A gnd NOR3X1_4/C vdd BUFX4
XBUFX4_61 BUFX4_62/A gnd BUFX4_61/Y vdd BUFX4
XBUFX4_72 INVX8_1/Y gnd BUFX4_72/Y vdd BUFX4
XBUFX4_83 INVX8_9/Y gnd BUFX4_83/Y vdd BUFX4
XBUFX4_94 BUFX4_98/A gnd BUFX4_94/Y vdd BUFX4
XOR2X2_20 OR2X2_20/A OR2X2_20/B gnd OR2X2_20/Y vdd OR2X2
XOR2X2_42 OR2X2_42/A OR2X2_42/B gnd OR2X2_42/Y vdd OR2X2
XOR2X2_31 OR2X2_31/A OR2X2_31/B gnd OR2X2_31/Y vdd OR2X2
XOR2X2_64 OR2X2_64/A OR2X2_64/B gnd OR2X2_64/Y vdd OR2X2
XOR2X2_53 OR2X2_53/A OR2X2_53/B gnd OR2X2_53/Y vdd OR2X2
XOR2X2_2 OR2X2_2/A OR2X2_2/B gnd OR2X2_2/Y vdd OR2X2
XXNOR2X1_4 XOR2X1_2/A INVX2_74/A gnd NAND3X1_3/C vdd XNOR2X1
XFILL_40_0_1 gnd vdd FILL
XINVX1_4 gnd gnd INVX1_4/Y vdd INVX1
XOAI21X1_540 INVX1_392/Y OAI22X1_9/C INVX1_393/A gnd NAND3X1_130/C vdd OAI21X1
XOAI21X1_551 OAI21X1_551/A NOR2X1_108/A AOI21X1_113/Y gnd OR2X2_32/A vdd OAI21X1
XOAI21X1_573 INVX2_61/Y NOR2X1_304/A OAI21X1_602/B gnd AND2X2_47/A vdd OAI21X1
XOAI21X1_562 NAND2X1_500/B NOR2X1_281/A BUFX4_92/Y gnd NOR2X1_282/A vdd OAI21X1
XOAI21X1_584 INVX8_5/A OAI21X1_612/A NAND2X1_526/Y gnd NAND2X1_547/B vdd OAI21X1
XOAI21X1_595 INVX1_399/A AOI21X1_180/B OAI21X1_595/C gnd OAI21X1_595/Y vdd OAI21X1
XINVX1_626 INVX1_553/A gnd INVX1_626/Y vdd INVX1
XINVX1_604 INVX1_604/A gnd INVX1_604/Y vdd INVX1
XINVX1_615 INVX1_542/A gnd INVX1_615/Y vdd INVX1
XINVX1_648 BUFX2_92/A gnd INVX1_648/Y vdd INVX1
XINVX1_637 INVX1_637/A gnd INVX1_637/Y vdd INVX1
XINVX1_659 OR2X2_50/B gnd INVX1_659/Y vdd INVX1
XNAND2X1_590 MUX2X1_49/S NAND2X1_590/B gnd OAI21X1_738/C vdd NAND2X1
XFILL_31_0_1 gnd vdd FILL
XFILL_39_1_1 gnd vdd FILL
XFILL_22_0_1 gnd vdd FILL
XBUFX4_209 BUFX4_210/A gnd BUFX4_209/Y vdd BUFX4
XFILL_5_1_1 gnd vdd FILL
XFILL_13_0_1 gnd vdd FILL
XOAI21X1_392 INVX8_8/A MUX2X1_14/Y OAI21X1_392/C gnd OAI21X1_394/B vdd OAI21X1
XINVX1_401 INVX1_401/A gnd INVX1_401/Y vdd INVX1
XOAI21X1_370 AOI21X1_54/Y INVX1_357/Y OAI21X1_370/C gnd AOI21X1_57/B vdd OAI21X1
XOAI21X1_381 INVX2_25/Y INVX8_8/A INVX8_5/A gnd OAI21X1_381/Y vdd OAI21X1
XAND2X2_4 AND2X2_4/A AND2X2_4/B gnd AND2X2_4/Y vdd AND2X2
XINVX1_412 INVX1_412/A gnd INVX1_412/Y vdd INVX1
XINVX1_423 INVX1_423/A gnd INVX1_423/Y vdd INVX1
XINVX1_434 INVX1_434/A gnd INVX1_434/Y vdd INVX1
XINVX1_478 BUFX2_55/A gnd INVX1_478/Y vdd INVX1
XINVX1_456 OR2X2_56/B gnd INVX1_456/Y vdd INVX1
XINVX1_467 INVX1_467/A gnd INVX1_467/Y vdd INVX1
XINVX1_445 INVX2_84/A gnd INVX1_445/Y vdd INVX1
XINVX1_489 BUFX2_68/A gnd INVX1_489/Y vdd INVX1
XFILL_2_4 gnd vdd FILL
XFILL_37_3 gnd vdd FILL
XMUX2X1_27 MUX2X1_27/A MUX2X1_27/B INVX8_4/A gnd MUX2X1_27/Y vdd MUX2X1
XMUX2X1_16 INVX1_247/A INVX1_690/A INVX4_4/A gnd MUX2X1_16/Y vdd MUX2X1
XMUX2X1_38 MUX2X1_38/A MUX2X1_38/B BUFX4_51/Y gnd MUX2X1_38/Y vdd MUX2X1
XMUX2X1_49 MUX2X1_49/A MUX2X1_49/B MUX2X1_49/S gnd MUX2X1_49/Y vdd MUX2X1
XINVX1_253 INVX1_253/A gnd INVX1_253/Y vdd INVX1
XINVX1_242 INVX1_242/A gnd NOR3X1_50/A vdd INVX1
XINVX1_231 NOR2X1_6/B gnd INVX1_231/Y vdd INVX1
XINVX1_220 INVX1_220/A gnd INVX1_220/Y vdd INVX1
XINVX1_275 INVX1_275/A gnd INVX1_275/Y vdd INVX1
XINVX1_264 INVX1_264/A gnd OR2X2_10/B vdd INVX1
XINVX1_286 INVX1_286/A gnd INVX1_286/Y vdd INVX1
XINVX1_297 INVX1_297/A gnd INVX1_297/Y vdd INVX1
XNAND2X1_20 BUFX4_24/Y NAND2X1_20/B gnd OAI21X1_20/C vdd NAND2X1
XNAND2X1_31 BUFX4_20/Y NAND2X1_31/B gnd OAI21X1_31/C vdd NAND2X1
XNAND2X1_42 BUFX4_32/Y NAND2X1_42/B gnd OAI21X1_42/C vdd NAND2X1
XNAND2X1_75 INVX2_8/A BUFX4_162/Y gnd NAND2X1_75/Y vdd NAND2X1
XNAND2X1_86 INVX1_268/A BUFX4_158/Y gnd NAND2X1_86/Y vdd NAND2X1
XNAND2X1_64 BUFX4_32/Y NAND2X1_64/B gnd NAND2X1_64/Y vdd NAND2X1
XNAND2X1_53 BUFX4_27/Y NAND2X1_53/B gnd NAND2X1_53/Y vdd NAND2X1
XNAND2X1_97 INVX1_296/A BUFX4_163/Y gnd NAND2X1_97/Y vdd NAND2X1
XAOI21X1_213 INVX2_65/A OAI21X1_779/Y OAI21X1_782/Y gnd AOI21X1_213/Y vdd AOI21X1
XAOI21X1_202 OAI21X1_334/C NOR2X1_354/Y INVX1_349/A gnd OAI21X1_750/C vdd AOI21X1
XAOI21X1_224 INVX2_74/A INVX1_502/Y INVX1_504/Y gnd AOI21X1_224/Y vdd AOI21X1
XAOI21X1_257 AOI21X1_263/A AOI21X1_257/B OAI22X1_53/Y gnd OAI21X1_982/A vdd AOI21X1
XAOI21X1_246 OAI21X1_907/C AOI21X1_246/B OAI21X1_927/Y gnd AOI21X1_246/Y vdd AOI21X1
XAOI21X1_235 AOI21X1_234/Y OAI21X1_907/Y OR2X2_68/A gnd AOI21X1_235/Y vdd AOI21X1
XAOI21X1_268 OAI21X1_992/B NOR2X1_475/Y BUFX2_37/A gnd AOI21X1_271/A vdd AOI21X1
XAOI22X1_40 INVX1_224/Y AND2X2_8/B INVX1_223/Y NOR2X1_13/Y gnd AOI22X1_40/Y vdd AOI22X1
XAOI22X1_51 MUX2X1_4/A BUFX4_235/Y BUFX4_151/Y MUX2X1_4/B gnd NOR2X1_37/B vdd AOI22X1
XAOI22X1_73 AOI22X1_73/A AOI21X1_97/A AOI22X1_73/C AOI22X1_73/D gnd AOI21X1_77/A vdd
+ AOI22X1
XAOI22X1_84 OR2X2_28/Y AOI21X1_84/Y AOI22X1_84/C BUFX4_77/Y gnd AOI22X1_84/Y vdd AOI22X1
XAOI22X1_62 AOI22X1_62/A BUFX4_233/Y BUFX4_148/Y INVX1_306/A gnd NOR2X1_53/B vdd AOI22X1
XAOI22X1_95 AND2X2_43/Y AOI22X1_95/B AOI22X1_95/C BUFX4_78/Y gnd AOI22X1_95/Y vdd
+ AOI22X1
XNAND3X1_217 BUFX4_218/Y NAND3X1_217/B NAND3X1_217/C gnd NAND2X1_750/B vdd NAND3X1
XNAND3X1_206 INVX1_520/Y BUFX4_206/Y BUFX4_33/Y gnd NAND3X1_207/B vdd NAND3X1
XNAND3X1_239 BUFX4_219/Y NAND3X1_238/Y NAND3X1_239/C gnd NAND2X1_783/B vdd NAND3X1
XNAND3X1_228 INVX1_542/Y BUFX4_208/Y BUFX4_36/Y gnd NAND3X1_228/Y vdd NAND3X1
XOAI22X1_2 INVX2_2/Y OR2X2_52/B INVX2_3/A AOI22X1_3/D gnd NOR3X1_16/A vdd OAI22X1
XFILL_30_6_0 gnd vdd FILL
XDFFPOSX1_316 INVX1_258/A CLKBUF1_12/Y OAI21X1_884/Y gnd vdd DFFPOSX1
XDFFPOSX1_327 INVX1_278/A CLKBUF1_1/Y OAI21X1_895/Y gnd vdd DFFPOSX1
XDFFPOSX1_305 INVX2_6/A CLKBUF1_49/Y OAI21X1_878/Y gnd vdd DFFPOSX1
XDFFPOSX1_338 INVX2_1/A CLKBUF1_9/Y NOR2X1_22/B gnd vdd DFFPOSX1
XDFFPOSX1_349 INVX2_85/A CLKBUF1_58/Y OAI21X1_6/Y gnd vdd DFFPOSX1
XNAND2X1_408 INVX8_5/A INVX2_52/A gnd NAND2X1_408/Y vdd NAND2X1
XNAND2X1_419 INVX8_4/A MUX2X1_32/B gnd OAI21X1_438/C vdd NAND2X1
XFILL_38_7_0 gnd vdd FILL
XNOR2X1_430 NOR2X1_428/Y NOR2X1_429/Y gnd NOR2X1_430/Y vdd NOR2X1
XNOR2X1_441 INVX1_449/A INVX1_679/Y gnd NOR2X1_441/Y vdd NOR2X1
XNOR2X1_452 NOR2X1_424/B NOR2X1_452/B gnd NOR2X1_454/B vdd NOR2X1
XNOR2X1_463 MUX2X1_7/B OR2X2_58/B gnd NOR2X1_463/Y vdd NOR2X1
XNOR2X1_485 OAI22X1_60/Y NOR2X1_485/B gnd NOR2X1_485/Y vdd NOR2X1
XNOR2X1_474 INVX8_17/Y NOR2X1_474/B gnd NOR2X1_474/Y vdd NOR2X1
XOAI21X1_903 INVX2_82/Y INVX1_459/A NAND3X1_337/A gnd NOR2X1_425/A vdd OAI21X1
XFILL_21_6_0 gnd vdd FILL
XOAI21X1_925 AOI21X1_240/Y OAI21X1_925/B NOR2X1_422/Y gnd OAI21X1_925/Y vdd OAI21X1
XOAI21X1_914 INVX1_669/A INVX1_670/Y AND2X2_82/A gnd NOR3X1_71/A vdd OAI21X1
XOAI21X1_936 NOR2X1_424/B NOR2X1_452/B OAI21X1_936/C gnd AOI21X1_254/C vdd OAI21X1
XOAI21X1_958 INVX8_17/Y INVX8_15/Y BUFX2_80/A gnd OAI21X1_959/C vdd OAI21X1
XOAI21X1_947 NOR3X1_77/Y NOR3X1_78/Y NOR2X1_477/Y gnd OAI22X1_58/B vdd OAI21X1
XOAI21X1_969 INVX1_727/Y BUFX4_116/Y OAI21X1_969/C gnd OAI21X1_969/Y vdd OAI21X1
XINVX2_11 INVX2_11/A gnd INVX2_11/Y vdd INVX2
XINVX2_33 INVX2_33/A gnd INVX2_33/Y vdd INVX2
XINVX2_44 INVX2_44/A gnd INVX2_44/Y vdd INVX2
XINVX2_22 INVX2_22/A gnd INVX2_22/Y vdd INVX2
XNAND2X1_931 OR2X2_53/A OR2X2_53/B gnd AOI22X1_126/A vdd NAND2X1
XNAND2X1_920 NOR2X1_22/B INVX1_643/Y gnd OAI22X1_49/B vdd NAND2X1
XINVX2_66 INVX2_66/A gnd INVX2_66/Y vdd INVX2
XINVX2_55 INVX2_55/A gnd INVX2_55/Y vdd INVX2
XNAND2X1_942 OR2X2_56/A OR2X2_56/B gnd AOI22X1_128/A vdd NAND2X1
XNAND2X1_964 MUX2X1_7/B INVX1_692/Y gnd AND2X2_88/B vdd NAND2X1
XNAND2X1_953 MUX2X1_9/B INVX2_84/Y gnd AND2X2_87/B vdd NAND2X1
XINVX2_77 BUFX2_90/A gnd INVX2_77/Y vdd INVX2
XINVX2_88 INVX2_88/A gnd INVX2_88/Y vdd INVX2
XNAND2X1_975 AOI21X1_251/B AOI21X1_251/A gnd NAND2X1_975/Y vdd NAND2X1
XNAND2X1_986 INVX1_451/A INVX1_675/Y gnd NAND2X1_987/B vdd NAND2X1
XNAND2X1_997 NAND3X1_1/B NOR2X1_3/A gnd NOR3X1_75/C vdd NAND2X1
XFILL_4_7_0 gnd vdd FILL
XFILL_29_7_0 gnd vdd FILL
XOAI21X1_18 INVX1_18/Y BUFX4_18/Y OAI21X1_18/C gnd OAI21X1_18/Y vdd OAI21X1
XOAI21X1_29 INVX1_29/Y BUFX4_22/Y OAI21X1_29/C gnd OAI21X1_29/Y vdd OAI21X1
XFILL_12_6_0 gnd vdd FILL
XFILL_12_2 gnd vdd FILL
XDFFPOSX1_102 INVX1_215/A CLKBUF1_63/Y OAI21X1_145/C gnd vdd DFFPOSX1
XDFFPOSX1_135 DFFPOSX1_23/D CLKBUF1_18/Y INVX2_13/A gnd vdd DFFPOSX1
XDFFPOSX1_146 DFFPOSX1_34/D CLKBUF1_24/Y INVX1_283/A gnd vdd DFFPOSX1
XDFFPOSX1_124 DFFPOSX1_12/D CLKBUF1_42/Y INVX1_234/A gnd vdd DFFPOSX1
XDFFPOSX1_113 OR2X2_69/B CLKBUF1_62/Y NOR2X1_1/A gnd vdd DFFPOSX1
XDFFPOSX1_168 BUFX2_11/A CLKBUF1_26/Y XNOR2X1_22/Y gnd vdd DFFPOSX1
XDFFPOSX1_179 BUFX2_22/A CLKBUF1_35/Y XNOR2X1_41/Y gnd vdd DFFPOSX1
XDFFPOSX1_157 INVX1_504/A CLKBUF1_43/Y INVX1_572/A gnd vdd DFFPOSX1
XNAND2X1_216 INVX2_69/A INVX1_410/A gnd INVX4_10/A vdd NAND2X1
XNAND2X1_205 INVX4_4/A AOI22X1_67/A gnd NAND2X1_205/Y vdd NAND2X1
XNAND2X1_227 INVX2_35/A MUX2X1_42/B gnd INVX1_402/A vdd NAND2X1
XNAND2X1_238 INVX2_68/A NAND2X1_237/Y gnd INVX2_67/A vdd NAND2X1
XNAND2X1_249 INVX2_41/A MUX2X1_37/A gnd OAI21X1_588/C vdd NAND2X1
XNOR2X1_260 BUFX4_58/Y AND2X2_44/A gnd NOR2X1_260/Y vdd NOR2X1
XNOR2X1_271 BUFX4_52/Y NOR2X1_271/B gnd NOR2X1_271/Y vdd NOR2X1
XNOR2X1_293 NOR2X1_293/A AND2X2_46/Y gnd NOR2X1_293/Y vdd NOR2X1
XNOR2X1_282 NOR2X1_282/A NOR2X1_281/Y gnd NOR2X1_282/Y vdd NOR2X1
XOAI21X1_711 INVX1_328/Y INVX1_413/Y AND2X2_62/B gnd AOI21X1_186/C vdd OAI21X1
XOAI21X1_700 OAI21X1_700/A BUFX4_225/Y OAI21X1_700/C gnd NAND2X1_595/B vdd OAI21X1
XOAI21X1_733 INVX2_18/Y OAI21X1_732/Y NOR2X1_350/Y gnd NAND3X1_165/B vdd OAI21X1
XOAI21X1_722 OAI21X1_743/A NOR2X1_356/A OAI21X1_722/C gnd OAI21X1_722/Y vdd OAI21X1
XOAI21X1_766 OAI21X1_745/Y AND2X2_70/B MUX2X1_20/S gnd OAI22X1_44/B vdd OAI21X1
XOAI21X1_755 INVX2_20/A INVX2_21/Y INVX2_71/A gnd OAI21X1_755/Y vdd OAI21X1
XOAI21X1_744 INVX2_22/A OAI21X1_744/B NOR2X1_358/Y gnd NAND3X1_169/A vdd OAI21X1
XOAI21X1_777 MUX2X1_49/S NAND2X1_590/B OAI21X1_776/Y gnd AND2X2_74/A vdd OAI21X1
XOAI21X1_788 BUFX4_180/Y INVX1_441/Y NAND2X1_611/Y gnd OAI21X1_788/Y vdd OAI21X1
XOAI21X1_799 BUFX4_181/Y INVX1_452/Y NAND2X1_622/Y gnd OAI21X1_799/Y vdd OAI21X1
XNAND2X1_772 OAI21X1_86/Y BUFX4_134/Y gnd NAND2X1_774/A vdd NAND2X1
XNAND2X1_750 NAND2X1_750/A NAND2X1_750/B gnd NAND2X1_14/B vdd NAND2X1
XNAND2X1_761 INVX1_537/Y BUFX4_201/Y gnd NAND3X1_225/C vdd NAND2X1
XNAND2X1_783 NAND2X1_783/A NAND2X1_783/B gnd NAND2X1_25/B vdd NAND2X1
XNAND2X1_794 INVX1_559/Y BUFX4_204/Y gnd NAND3X1_247/C vdd NAND2X1
XCLKBUF1_19 BUFX4_4/Y gnd CLKBUF1_19/Y vdd CLKBUF1
XBUFX4_51 INVX8_3/Y gnd BUFX4_51/Y vdd BUFX4
XBUFX4_40 INVX8_8/Y gnd BUFX4_40/Y vdd BUFX4
XBUFX4_62 BUFX4_62/A gnd BUFX4_62/Y vdd BUFX4
XBUFX4_84 INVX8_9/Y gnd BUFX4_84/Y vdd BUFX4
XBUFX4_73 INVX8_1/Y gnd BUFX4_73/Y vdd BUFX4
XBUFX4_95 BUFX4_98/A gnd BUFX4_95/Y vdd BUFX4
XFILL_35_5_0 gnd vdd FILL
XOR2X2_32 OR2X2_32/A OR2X2_32/B gnd OR2X2_32/Y vdd OR2X2
XOR2X2_21 OR2X2_21/A OR2X2_21/B gnd OR2X2_21/Y vdd OR2X2
XOR2X2_10 OR2X2_10/A OR2X2_10/B gnd OR2X2_10/Y vdd OR2X2
XOR2X2_65 OR2X2_65/A OR2X2_63/B gnd OR2X2_65/Y vdd OR2X2
XOR2X2_43 OR2X2_43/A INVX2_28/Y gnd OR2X2_43/Y vdd OR2X2
XOR2X2_54 OR2X2_54/A OR2X2_54/B gnd OR2X2_54/Y vdd OR2X2
XOR2X2_3 OR2X2_3/A OR2X2_3/B gnd OR2X2_3/Y vdd OR2X2
XXNOR2X1_5 XNOR2X1_5/A AOI21X1_5/Y gnd XNOR2X1_5/Y vdd XNOR2X1
XFILL_26_5_0 gnd vdd FILL
XFILL_1_5_0 gnd vdd FILL
XINVX8_10 INVX8_10/A gnd BUFX4_93/A vdd INVX8
XINVX1_5 gnd gnd INVX1_5/Y vdd INVX1
XOAI21X1_530 AND2X2_41/A INVX2_59/Y BUFX4_92/Y gnd NOR2X1_255/A vdd OAI21X1
XOAI21X1_541 INVX1_393/A NOR2X1_269/Y OAI21X1_541/C gnd OAI21X1_541/Y vdd OAI21X1
XOAI21X1_574 AND2X2_47/A INVX2_63/A INVX8_11/Y gnd OR2X2_34/B vdd OAI21X1
XOAI21X1_552 OAI22X1_8/B OAI22X1_8/A OR2X2_32/A gnd NOR2X1_281/B vdd OAI21X1
XOAI21X1_563 OAI22X1_29/A OAI21X1_561/Y NOR2X1_282/Y gnd OAI21X1_563/Y vdd OAI21X1
XINVX1_616 INVX1_543/A gnd INVX1_616/Y vdd INVX1
XOAI21X1_596 INVX1_398/Y BUFX4_217/Y OAI21X1_596/C gnd INVX2_66/A vdd OAI21X1
XOAI21X1_585 BUFX4_214/Y NAND2X1_497/B NAND2X1_527/Y gnd MUX2X1_38/A vdd OAI21X1
XINVX1_627 INVX1_554/A gnd INVX1_627/Y vdd INVX1
XINVX1_605 INVX1_532/A gnd INVX1_605/Y vdd INVX1
XINVX1_638 INVX1_565/A gnd INVX1_638/Y vdd INVX1
XINVX1_649 BUFX2_93/A gnd INVX1_649/Y vdd INVX1
.ends

