module AXI4_read 
(
    input axi_clk,
    input resetn   //axi is reset low

);
    
endmodule