module Control_Unit 
(
      input [6 : 0] opcode,
      input [2 : 0] funct3,
      input [6 : 0] funct7


      // Outputs :)))
);
      
endmodule