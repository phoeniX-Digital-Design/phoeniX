magic
tech scmos
timestamp 1693479267
<< metal1 >>
rect 496 4403 498 4407
rect 502 4403 505 4407
rect 509 4403 512 4407
rect 1520 4403 1522 4407
rect 1526 4403 1529 4407
rect 1533 4403 1536 4407
rect 2544 4403 2546 4407
rect 2550 4403 2553 4407
rect 2557 4403 2560 4407
rect 3568 4403 3570 4407
rect 3574 4403 3577 4407
rect 3581 4403 3584 4407
rect 4045 4378 4046 4382
rect 3018 4368 3033 4371
rect 3597 4368 3598 4372
rect 4202 4368 4203 4372
rect 42 4357 44 4361
rect 778 4358 782 4362
rect 2530 4358 2537 4361
rect 2894 4358 2905 4361
rect 3306 4358 3313 4361
rect 3622 4361 3625 4368
rect 54 4348 70 4351
rect 646 4348 665 4351
rect 794 4348 801 4351
rect 846 4348 854 4351
rect 918 4348 926 4351
rect 1478 4351 1482 4353
rect 1478 4348 1489 4351
rect 1558 4348 1577 4351
rect 1622 4348 1638 4351
rect 1718 4348 1726 4351
rect 1734 4348 1742 4351
rect 1790 4348 1809 4351
rect 2942 4348 2961 4351
rect 3166 4348 3174 4351
rect 3274 4348 3281 4351
rect 3582 4351 3585 4361
rect 3614 4358 3625 4361
rect 3718 4358 3737 4361
rect 3946 4358 3950 4362
rect 3978 4358 3982 4362
rect 3550 4348 3585 4351
rect 3738 4348 3745 4351
rect 3798 4348 3806 4351
rect 4030 4351 4033 4361
rect 4014 4348 4033 4351
rect 4218 4348 4225 4351
rect 4282 4348 4289 4351
rect 14 4338 22 4341
rect 126 4338 153 4341
rect 466 4338 490 4341
rect 686 4338 694 4341
rect 486 4336 490 4338
rect 70 4328 78 4331
rect 886 4331 890 4336
rect 874 4328 890 4331
rect 902 4331 906 4333
rect 1134 4332 1137 4342
rect 1190 4338 1202 4341
rect 1678 4338 1697 4341
rect 2222 4338 2233 4341
rect 2358 4338 2369 4341
rect 2390 4338 2401 4341
rect 2438 4338 2446 4341
rect 2470 4338 2481 4341
rect 2502 4338 2513 4341
rect 2550 4338 2577 4341
rect 2622 4338 2633 4341
rect 2650 4338 2657 4341
rect 2918 4338 2929 4341
rect 3606 4338 3617 4341
rect 3854 4338 3865 4341
rect 3898 4338 3905 4341
rect 4302 4341 4305 4348
rect 4302 4338 4313 4341
rect 4502 4338 4518 4341
rect 1678 4336 1682 4338
rect 1270 4332 1274 4336
rect 902 4328 913 4331
rect 1822 4331 1826 4333
rect 1814 4328 1826 4331
rect 2214 4328 2217 4338
rect 2374 4328 2385 4331
rect 2486 4328 2497 4331
rect 2582 4328 2593 4331
rect 2638 4328 2649 4331
rect 2878 4331 2882 4333
rect 2926 4332 2929 4338
rect 2878 4328 2886 4331
rect 2994 4328 3001 4331
rect 4098 4328 4105 4331
rect 378 4318 380 4322
rect 444 4318 446 4322
rect 626 4318 627 4322
rect 994 4318 1009 4321
rect 2186 4318 2187 4322
rect 2349 4318 2350 4322
rect 2410 4318 2411 4322
rect 2461 4318 2462 4322
rect 2522 4318 2523 4322
rect 2541 4318 2542 4322
rect 2613 4318 2614 4322
rect 2909 4318 2910 4322
rect 4069 4318 4070 4322
rect 1000 4303 1002 4307
rect 1006 4303 1009 4307
rect 1013 4303 1016 4307
rect 2024 4303 2026 4307
rect 2030 4303 2033 4307
rect 2037 4303 2040 4307
rect 3048 4303 3050 4307
rect 3054 4303 3057 4307
rect 3061 4303 3064 4307
rect 4080 4303 4082 4307
rect 4086 4303 4089 4307
rect 4093 4303 4096 4307
rect 332 4288 334 4292
rect 2246 4288 2254 4291
rect 3245 4288 3246 4292
rect 3517 4288 3518 4292
rect 70 4278 78 4281
rect 466 4278 482 4281
rect 1046 4278 1054 4282
rect 1182 4278 1193 4281
rect 478 4277 482 4278
rect 1046 4272 1049 4278
rect 1478 4272 1481 4281
rect 2418 4278 2425 4281
rect 3332 4278 3334 4282
rect 3390 4278 3401 4281
rect 3558 4278 3585 4281
rect 14 4268 22 4271
rect 582 4268 609 4271
rect 58 4258 70 4261
rect 294 4258 302 4261
rect 866 4258 873 4261
rect 902 4258 910 4261
rect 990 4258 1025 4261
rect 1030 4258 1038 4261
rect 1086 4261 1089 4271
rect 1374 4268 1386 4271
rect 1486 4268 1494 4271
rect 1670 4271 1674 4274
rect 1670 4268 1689 4271
rect 2042 4268 2057 4271
rect 2860 4268 2862 4272
rect 3598 4268 3625 4271
rect 3674 4268 3689 4271
rect 3822 4268 3841 4271
rect 4158 4268 4166 4271
rect 1086 4258 1102 4261
rect 1122 4258 1137 4261
rect 1958 4258 1977 4261
rect 2030 4258 2065 4261
rect 2542 4258 2558 4261
rect 3022 4258 3033 4261
rect 3062 4258 3089 4261
rect 3110 4258 3121 4261
rect 3770 4258 3777 4261
rect 3902 4261 3905 4268
rect 3894 4258 3905 4261
rect 3922 4258 3929 4261
rect 3934 4258 3953 4261
rect 3966 4258 3974 4261
rect 4030 4258 4038 4261
rect 4070 4258 4086 4261
rect 4174 4261 4177 4271
rect 4230 4268 4249 4271
rect 4414 4268 4433 4271
rect 4522 4268 4529 4271
rect 4166 4258 4177 4261
rect 4190 4258 4198 4261
rect 4222 4258 4230 4261
rect 4286 4258 4294 4261
rect 4382 4258 4390 4261
rect 4434 4258 4441 4261
rect 4510 4258 4529 4261
rect 1066 4248 1073 4251
rect 2014 4248 2022 4251
rect 2222 4248 2230 4251
rect 2238 4248 2249 4251
rect 2334 4248 2342 4251
rect 2438 4251 2441 4258
rect 2398 4248 2409 4251
rect 2430 4248 2441 4251
rect 2462 4248 2473 4251
rect 2510 4248 2521 4251
rect 2622 4248 2630 4251
rect 2734 4248 2745 4251
rect 2898 4248 2905 4251
rect 3270 4248 3281 4251
rect 3354 4248 3358 4252
rect 3750 4248 3769 4251
rect 3950 4248 3953 4258
rect 4526 4248 4529 4258
rect 251 4238 254 4242
rect 818 4238 833 4241
rect 2454 4241 2457 4248
rect 2446 4238 2457 4241
rect 2626 4238 2649 4241
rect 2746 4238 2761 4241
rect 2794 4238 2825 4241
rect 454 4228 470 4231
rect 1826 4218 1827 4222
rect 496 4203 498 4207
rect 502 4203 505 4207
rect 509 4203 512 4207
rect 1520 4203 1522 4207
rect 1526 4203 1529 4207
rect 1533 4203 1536 4207
rect 2544 4203 2546 4207
rect 2550 4203 2553 4207
rect 2557 4203 2560 4207
rect 3568 4203 3570 4207
rect 3574 4203 3577 4207
rect 3581 4203 3584 4207
rect 941 4188 942 4192
rect 1794 4188 1795 4192
rect 1826 4188 1827 4192
rect 2022 4188 2030 4191
rect 3373 4188 3374 4192
rect 3469 4188 3470 4192
rect 3898 4188 3899 4192
rect 878 4172 881 4181
rect 2198 4168 2209 4171
rect 2978 4168 2985 4171
rect 3002 4168 3005 4172
rect 3314 4168 3345 4171
rect 113 4158 118 4162
rect 246 4158 254 4161
rect 558 4161 561 4168
rect 2206 4162 2209 4168
rect 494 4158 521 4161
rect 550 4158 561 4161
rect 578 4158 585 4161
rect 590 4158 598 4161
rect 622 4158 633 4161
rect 654 4158 665 4161
rect 266 4148 273 4151
rect 758 4148 777 4151
rect 846 4148 857 4151
rect 886 4151 890 4154
rect 1750 4152 1753 4161
rect 1990 4158 2001 4161
rect 2070 4158 2081 4161
rect 2150 4158 2161 4161
rect 2342 4158 2353 4161
rect 2942 4161 2945 4168
rect 2942 4158 2953 4161
rect 3146 4157 3148 4161
rect 3322 4158 3329 4161
rect 3758 4158 3766 4161
rect 3954 4158 3958 4162
rect 886 4148 905 4151
rect 910 4148 926 4151
rect 998 4148 1006 4151
rect 1054 4148 1073 4151
rect 1094 4148 1105 4151
rect 854 4142 857 4148
rect 14 4138 22 4141
rect 258 4138 265 4141
rect 458 4138 465 4141
rect 538 4138 545 4141
rect 750 4138 761 4141
rect 778 4138 785 4141
rect 910 4138 913 4148
rect 1270 4148 1278 4151
rect 1310 4148 1318 4151
rect 1462 4148 1481 4151
rect 1510 4148 1545 4151
rect 1766 4148 1774 4151
rect 1778 4148 1793 4151
rect 2226 4148 2233 4151
rect 950 4138 985 4141
rect 1274 4138 1289 4141
rect 1710 4138 1713 4148
rect 2878 4148 2889 4151
rect 2918 4148 2937 4151
rect 3118 4148 3126 4151
rect 3198 4148 3209 4151
rect 3214 4148 3225 4151
rect 3422 4148 3446 4151
rect 3470 4148 3486 4151
rect 3506 4148 3513 4151
rect 3586 4148 3617 4151
rect 3682 4148 3737 4151
rect 3790 4148 3814 4151
rect 3926 4148 3945 4151
rect 4030 4148 4038 4151
rect 4142 4148 4150 4151
rect 4166 4148 4174 4151
rect 4206 4151 4209 4161
rect 4250 4158 4254 4162
rect 4282 4158 4286 4162
rect 4190 4148 4209 4151
rect 4286 4148 4294 4151
rect 4338 4148 4345 4151
rect 4370 4148 4377 4151
rect 4382 4148 4401 4151
rect 4466 4148 4473 4151
rect 4522 4148 4529 4151
rect 2878 4142 2881 4148
rect 2974 4146 2978 4148
rect 3222 4142 3225 4148
rect 1774 4138 1782 4141
rect 1874 4138 1881 4141
rect 2294 4138 2305 4141
rect 2374 4138 2385 4141
rect 2402 4138 2409 4141
rect 2542 4138 2569 4141
rect 2630 4138 2641 4141
rect 3070 4138 3078 4141
rect 3082 4138 3094 4141
rect 3174 4138 3201 4141
rect 3302 4138 3310 4141
rect 3382 4138 3390 4141
rect 3578 4138 3625 4141
rect 3686 4138 3726 4141
rect 3878 4138 3889 4141
rect 3942 4138 3945 4148
rect 3998 4138 4006 4141
rect 4318 4138 4337 4141
rect 4422 4138 4438 4141
rect 4454 4141 4457 4148
rect 4454 4138 4465 4141
rect 70 4128 78 4131
rect 446 4131 450 4133
rect 446 4128 457 4131
rect 542 4128 545 4138
rect 998 4128 1025 4131
rect 1558 4131 1562 4133
rect 1550 4128 1562 4131
rect 2894 4131 2897 4138
rect 2894 4128 2905 4131
rect 3090 4128 3097 4131
rect 3174 4128 3177 4138
rect 3582 4128 3590 4131
rect 3682 4128 3689 4131
rect 4462 4128 4465 4138
rect 525 4118 526 4122
rect 618 4118 619 4122
rect 669 4118 670 4122
rect 821 4118 822 4122
rect 1949 4118 1950 4122
rect 2054 4118 2062 4121
rect 2180 4118 2182 4122
rect 2452 4118 2454 4122
rect 2502 4118 2510 4121
rect 3841 4118 3846 4122
rect 1000 4103 1002 4107
rect 1006 4103 1009 4107
rect 1013 4103 1016 4107
rect 2024 4103 2026 4107
rect 2030 4103 2033 4107
rect 2037 4103 2040 4107
rect 3048 4103 3050 4107
rect 3054 4103 3057 4107
rect 3061 4103 3064 4107
rect 4080 4103 4082 4107
rect 4086 4103 4089 4107
rect 4093 4103 4096 4107
rect 3309 4088 3310 4092
rect 3397 4088 3398 4092
rect 3562 4088 3577 4091
rect 876 4078 889 4081
rect 1010 4078 1022 4081
rect 1062 4078 1073 4081
rect 2158 4078 2169 4081
rect 3054 4078 3070 4081
rect 3236 4078 3238 4082
rect 4058 4078 4065 4081
rect 886 4072 889 4078
rect 178 4068 185 4071
rect 234 4068 241 4071
rect 274 4068 281 4071
rect 294 4068 302 4071
rect 318 4068 337 4071
rect 942 4068 958 4071
rect 990 4068 1001 4071
rect 1446 4068 1462 4071
rect 1498 4068 1505 4071
rect 1858 4068 1865 4071
rect 2326 4071 2330 4072
rect 2334 4071 2337 4078
rect 1890 4068 1897 4071
rect 2142 4068 2153 4071
rect 2230 4068 2241 4071
rect 2326 4068 2337 4071
rect 2438 4071 2442 4072
rect 2446 4071 2449 4078
rect 2438 4068 2449 4071
rect 2596 4068 2598 4072
rect 2658 4068 2665 4071
rect 3166 4068 3174 4071
rect 3270 4068 3289 4071
rect 3518 4068 3545 4071
rect 3630 4068 3641 4071
rect 3994 4068 4001 4071
rect 4022 4068 4041 4071
rect 4046 4068 4054 4071
rect 4090 4068 4113 4071
rect 4362 4068 4369 4071
rect 262 4058 270 4061
rect 302 4058 310 4061
rect 990 4062 993 4068
rect 662 4058 682 4061
rect 766 4058 782 4061
rect 790 4058 806 4061
rect 838 4058 858 4061
rect 1062 4061 1065 4068
rect 1054 4058 1065 4061
rect 1426 4058 1433 4061
rect 1466 4058 1473 4061
rect 1526 4058 1542 4061
rect 1782 4058 1801 4061
rect 1814 4058 1833 4061
rect 2774 4061 2777 4068
rect 2766 4058 2777 4061
rect 3202 4058 3209 4061
rect 3294 4058 3302 4061
rect 3542 4058 3558 4061
rect 3678 4058 3697 4061
rect 3790 4058 3806 4061
rect 3822 4058 3830 4061
rect 3970 4058 3977 4061
rect 3986 4058 4009 4061
rect 4086 4058 4094 4061
rect 4246 4058 4262 4061
rect 4330 4058 4337 4061
rect 4382 4058 4390 4061
rect 4406 4058 4422 4061
rect 678 4056 682 4058
rect 854 4056 858 4058
rect 478 4048 486 4051
rect 778 4048 785 4051
rect 802 4048 809 4051
rect 929 4048 934 4052
rect 1814 4048 1817 4058
rect 2910 4056 2914 4058
rect 1974 4048 1985 4051
rect 2022 4048 2049 4051
rect 2338 4048 2345 4051
rect 2390 4048 2401 4051
rect 2454 4048 2465 4051
rect 2566 4048 2577 4051
rect 3678 4048 3681 4058
rect 3926 4056 3930 4058
rect 4274 4048 4278 4052
rect 378 4038 385 4041
rect 428 4038 430 4042
rect 610 4038 617 4041
rect 682 4038 697 4041
rect 814 4038 830 4041
rect 858 4038 873 4041
rect 1171 4038 1174 4042
rect 2134 4038 2142 4041
rect 2222 4038 2230 4041
rect 2738 4038 2745 4041
rect 2886 4038 2910 4041
rect 2962 4038 2965 4042
rect 3045 4038 3046 4042
rect 3098 4038 3101 4042
rect 3198 4041 3201 4048
rect 3190 4038 3201 4041
rect 3302 4041 3306 4044
rect 3390 4041 3394 4044
rect 3294 4038 3306 4041
rect 3382 4038 3394 4041
rect 4469 4038 4470 4042
rect 213 4018 214 4022
rect 3621 4018 3622 4022
rect 3853 4018 3854 4022
rect 4338 4018 4339 4022
rect 496 4003 498 4007
rect 502 4003 505 4007
rect 509 4003 512 4007
rect 1520 4003 1522 4007
rect 1526 4003 1529 4007
rect 1533 4003 1536 4007
rect 2544 4003 2546 4007
rect 2550 4003 2553 4007
rect 2557 4003 2560 4007
rect 3568 4003 3570 4007
rect 3574 4003 3577 4007
rect 3581 4003 3584 4007
rect 570 3988 572 3992
rect 990 3988 1006 3991
rect 1781 3988 1782 3992
rect 1813 3988 1814 3992
rect 3034 3988 3049 3991
rect 1234 3968 1237 3972
rect 2346 3968 2353 3971
rect 2822 3968 2830 3971
rect 4546 3968 4547 3972
rect 750 3958 769 3961
rect 774 3958 785 3961
rect 878 3958 889 3961
rect 1410 3958 1417 3961
rect 1518 3958 1526 3961
rect 2854 3958 2862 3961
rect 3366 3958 3377 3961
rect 3542 3958 3550 3961
rect 3586 3958 3593 3961
rect 4078 3958 4086 3961
rect 4338 3958 4345 3961
rect 198 3948 222 3951
rect 390 3948 401 3951
rect 718 3948 729 3951
rect 814 3951 817 3958
rect 806 3948 817 3951
rect 1574 3948 1582 3951
rect 2094 3951 2097 3958
rect 3374 3952 3378 3954
rect 2086 3948 2097 3951
rect 2510 3948 2518 3951
rect 2562 3948 2569 3951
rect 14 3938 41 3941
rect 94 3938 121 3941
rect 238 3938 249 3941
rect 294 3938 302 3941
rect 350 3938 369 3941
rect 422 3938 441 3941
rect 502 3938 537 3941
rect 1854 3938 1862 3941
rect 1894 3941 1897 3948
rect 3098 3948 3105 3951
rect 3246 3948 3262 3951
rect 3382 3948 3385 3958
rect 3534 3948 3542 3951
rect 3558 3948 3590 3951
rect 3638 3948 3657 3951
rect 3834 3948 3849 3951
rect 4070 3948 4102 3951
rect 4282 3948 4289 3951
rect 4490 3948 4497 3951
rect 4558 3951 4561 3961
rect 4582 3961 4585 3968
rect 4582 3958 4593 3961
rect 4558 3948 4577 3951
rect 3654 3942 3657 3948
rect 1894 3938 1905 3941
rect 1942 3938 1953 3941
rect 2062 3938 2070 3941
rect 2102 3938 2113 3941
rect 2162 3938 2169 3941
rect 2262 3938 2273 3941
rect 2294 3938 2305 3941
rect 2534 3938 2550 3941
rect 2646 3938 2657 3941
rect 2758 3938 2769 3941
rect 2810 3938 2817 3941
rect 2870 3938 2881 3941
rect 3306 3938 3318 3941
rect 3894 3938 3902 3941
rect 3942 3938 3950 3941
rect 4046 3938 4057 3941
rect 4118 3938 4126 3941
rect 4230 3938 4238 3941
rect 4270 3938 4294 3941
rect 4390 3938 4409 3941
rect 74 3928 89 3931
rect 106 3928 113 3931
rect 790 3928 798 3931
rect 2078 3928 2081 3938
rect 2278 3928 2289 3931
rect 2662 3928 2665 3938
rect 2774 3928 2777 3938
rect 2830 3928 2833 3938
rect 3702 3928 3713 3931
rect 137 3918 142 3922
rect 850 3918 851 3922
rect 874 3918 875 3922
rect 1933 3918 1934 3922
rect 1974 3918 1982 3921
rect 2253 3918 2254 3922
rect 2637 3918 2638 3922
rect 2677 3918 2678 3922
rect 2716 3918 2718 3922
rect 4189 3918 4190 3922
rect 4269 3918 4270 3922
rect 4298 3918 4299 3922
rect 1000 3903 1002 3907
rect 1006 3903 1009 3907
rect 1013 3903 1016 3907
rect 2024 3903 2026 3907
rect 2030 3903 2033 3907
rect 2037 3903 2040 3907
rect 3048 3903 3050 3907
rect 3054 3903 3057 3907
rect 3061 3903 3064 3907
rect 4080 3903 4082 3907
rect 4086 3903 4089 3907
rect 4093 3903 4096 3907
rect 234 3888 236 3892
rect 434 3888 436 3892
rect 612 3888 614 3892
rect 726 3878 737 3881
rect 806 3878 817 3881
rect 982 3876 986 3878
rect 1718 3872 1721 3881
rect 2498 3878 2505 3881
rect 2958 3878 2969 3881
rect 3150 3878 3161 3881
rect 3330 3878 3346 3881
rect 262 3868 270 3871
rect 702 3868 710 3871
rect 750 3868 769 3871
rect 830 3868 849 3871
rect 938 3868 945 3871
rect 1194 3868 1201 3871
rect 1274 3868 1289 3871
rect 1302 3868 1326 3871
rect 1382 3868 1393 3871
rect 1762 3868 1769 3871
rect 1918 3868 1926 3871
rect 2012 3868 2022 3871
rect 2172 3868 2174 3872
rect 2442 3868 2449 3871
rect 2460 3868 2462 3872
rect 2742 3871 2746 3872
rect 2750 3871 2753 3878
rect 3342 3874 3346 3878
rect 3358 3878 3369 3881
rect 3678 3878 3689 3881
rect 3694 3878 3702 3881
rect 3950 3878 3961 3881
rect 3358 3877 3362 3878
rect 3678 3872 3681 3878
rect 2742 3868 2753 3871
rect 2942 3868 2953 3871
rect 3262 3868 3274 3871
rect 3374 3868 3385 3871
rect 3402 3868 3417 3871
rect 300 3858 302 3862
rect 406 3861 410 3864
rect 406 3858 436 3861
rect 1382 3862 1385 3868
rect 886 3858 897 3861
rect 1094 3858 1102 3861
rect 1246 3858 1265 3861
rect 1466 3858 1473 3861
rect 1654 3858 1662 3861
rect 1750 3858 1774 3861
rect 665 3848 670 3852
rect 1982 3848 1993 3851
rect 1790 3838 1801 3841
rect 2054 3841 2057 3861
rect 2258 3848 2265 3851
rect 2398 3848 2409 3851
rect 2478 3848 2489 3851
rect 2506 3848 2513 3851
rect 2054 3838 2073 3841
rect 2266 3838 2281 3841
rect 2554 3838 2585 3841
rect 2670 3841 2673 3861
rect 2894 3861 2897 3868
rect 2942 3862 2945 3868
rect 3718 3868 3729 3871
rect 2894 3858 2905 3861
rect 3718 3862 3721 3868
rect 4162 3868 4185 3871
rect 4338 3868 4345 3871
rect 4422 3868 4430 3871
rect 4482 3868 4502 3871
rect 4518 3868 4534 3871
rect 4538 3868 4545 3871
rect 3706 3858 3713 3861
rect 3850 3858 3857 3861
rect 3886 3858 3894 3861
rect 3926 3858 3934 3861
rect 3998 3858 4017 3861
rect 4082 3858 4113 3861
rect 4118 3858 4137 3861
rect 4262 3858 4270 3861
rect 4326 3858 4334 3861
rect 4338 3858 4353 3861
rect 4530 3858 4537 3861
rect 4566 3858 4590 3861
rect 2710 3848 2721 3851
rect 2754 3848 2761 3851
rect 2990 3848 3001 3851
rect 4014 3848 4017 3858
rect 4066 3848 4073 3851
rect 2670 3838 2689 3841
rect 2694 3838 2702 3841
rect 3074 3838 3097 3841
rect 496 3803 498 3807
rect 502 3803 505 3807
rect 509 3803 512 3807
rect 1520 3803 1522 3807
rect 1526 3803 1529 3807
rect 1533 3803 1536 3807
rect 2544 3803 2546 3807
rect 2550 3803 2553 3807
rect 2557 3803 2560 3807
rect 3568 3803 3570 3807
rect 3574 3803 3577 3807
rect 3581 3803 3584 3807
rect 1882 3788 1883 3792
rect 1962 3788 1963 3792
rect 2266 3768 2273 3771
rect 2958 3768 2966 3771
rect 3414 3768 3426 3771
rect 3414 3762 3417 3768
rect 3422 3766 3426 3768
rect 3718 3766 3722 3768
rect 42 3757 44 3761
rect 649 3758 654 3762
rect 1682 3758 1689 3761
rect 54 3748 94 3751
rect 118 3748 126 3751
rect 130 3748 142 3751
rect 958 3748 966 3751
rect 1230 3751 1234 3753
rect 1222 3748 1234 3751
rect 1342 3748 1369 3751
rect 1462 3748 1478 3751
rect 1670 3748 1678 3751
rect 1830 3751 1833 3761
rect 1830 3748 1849 3751
rect 1894 3751 1897 3761
rect 2610 3758 2617 3761
rect 2718 3758 2729 3761
rect 2782 3758 2793 3761
rect 2838 3758 2849 3761
rect 3126 3752 3129 3761
rect 3146 3758 3153 3761
rect 3158 3758 3177 3761
rect 3266 3758 3270 3762
rect 3398 3752 3401 3761
rect 1894 3748 1913 3751
rect 1942 3748 1961 3751
rect 2006 3748 2014 3751
rect 2082 3748 2089 3751
rect 2422 3748 2433 3751
rect 2458 3748 2465 3751
rect 2546 3748 2561 3751
rect 2422 3742 2425 3748
rect 3450 3748 3457 3751
rect 3702 3751 3706 3752
rect 3718 3751 3721 3761
rect 3546 3748 3553 3751
rect 3702 3748 3721 3751
rect 3726 3748 3734 3751
rect 4046 3748 4054 3751
rect 4338 3748 4345 3751
rect 4542 3748 4566 3751
rect 14 3738 22 3741
rect 742 3738 758 3741
rect 778 3738 785 3741
rect 870 3732 873 3742
rect 1350 3738 1358 3741
rect 1378 3738 1385 3741
rect 1926 3738 1934 3741
rect 2202 3738 2209 3741
rect 2246 3738 2262 3741
rect 2582 3738 2593 3741
rect 2630 3738 2641 3741
rect 2662 3738 2673 3741
rect 3054 3738 3081 3741
rect 3142 3738 3150 3741
rect 3198 3738 3209 3741
rect 3238 3738 3246 3741
rect 3278 3738 3289 3741
rect 3470 3738 3481 3741
rect 3774 3738 3809 3741
rect 4042 3738 4065 3741
rect 4210 3738 4217 3741
rect 4242 3738 4249 3741
rect 4390 3738 4398 3741
rect 4490 3738 4497 3741
rect 4554 3738 4561 3741
rect 70 3728 86 3731
rect 1486 3728 1494 3731
rect 1710 3731 1714 3733
rect 1702 3728 1714 3731
rect 2566 3728 2577 3731
rect 2646 3728 2657 3731
rect 2886 3728 2889 3738
rect 2942 3728 2945 3738
rect 3806 3732 3809 3738
rect 708 3718 710 3722
rect 2501 3718 2502 3722
rect 2621 3718 2622 3722
rect 2682 3718 2683 3722
rect 2901 3718 2902 3722
rect 3429 3718 3430 3722
rect 3582 3718 3590 3721
rect 3957 3718 3958 3722
rect 3997 3718 3998 3722
rect 4037 3718 4038 3722
rect 1000 3703 1002 3707
rect 1006 3703 1009 3707
rect 1013 3703 1016 3707
rect 2024 3703 2026 3707
rect 2030 3703 2033 3707
rect 2037 3703 2040 3707
rect 3048 3703 3050 3707
rect 3054 3703 3057 3707
rect 3061 3703 3064 3707
rect 4080 3703 4082 3707
rect 4086 3703 4089 3707
rect 4093 3703 4096 3707
rect 518 3688 534 3691
rect 2362 3688 2363 3692
rect 50 3678 57 3681
rect 74 3678 89 3681
rect 1446 3672 1449 3681
rect 2396 3678 2398 3682
rect 2598 3678 2609 3681
rect 3062 3681 3065 3688
rect 3050 3678 3065 3681
rect 3966 3678 3977 3681
rect 3966 3677 3970 3678
rect 14 3668 41 3671
rect 94 3668 102 3671
rect 162 3668 170 3671
rect 598 3668 609 3671
rect 1542 3668 1570 3671
rect 2614 3668 2625 3671
rect 2906 3668 2913 3671
rect 3342 3668 3353 3671
rect 3406 3668 3414 3671
rect 3418 3668 3425 3671
rect 3470 3668 3481 3671
rect 3533 3668 3534 3672
rect 3582 3668 3610 3671
rect 3718 3668 3726 3671
rect 3758 3668 3769 3671
rect 3870 3668 3882 3671
rect 4222 3668 4233 3671
rect 4290 3668 4297 3671
rect 4350 3668 4361 3671
rect 4462 3668 4486 3671
rect 4566 3668 4574 3671
rect 366 3658 374 3661
rect 1134 3658 1153 3661
rect 1278 3658 1297 3661
rect 1422 3658 1441 3661
rect 1870 3658 1878 3661
rect 2638 3661 2641 3668
rect 2630 3658 2641 3661
rect 2726 3661 2729 3668
rect 2718 3658 2729 3661
rect 3834 3658 3841 3661
rect 3982 3658 4001 3661
rect 4222 3661 4225 3668
rect 4210 3658 4225 3661
rect 4246 3658 4254 3661
rect 4278 3658 4286 3661
rect 4350 3661 4353 3668
rect 4342 3658 4353 3661
rect 4510 3658 4518 3661
rect 4546 3658 4553 3661
rect 122 3649 124 3653
rect 2246 3648 2257 3651
rect 2430 3648 2441 3651
rect 2878 3648 2889 3651
rect 3038 3651 3041 3658
rect 2982 3648 2993 3651
rect 3030 3648 3041 3651
rect 3294 3648 3297 3658
rect 3302 3648 3321 3651
rect 3374 3648 3393 3651
rect 3398 3648 3409 3651
rect 4034 3648 4038 3652
rect 4342 3648 4345 3658
rect 3406 3642 3409 3648
rect 819 3638 822 3642
rect 2162 3638 2169 3641
rect 2194 3638 2217 3641
rect 2266 3638 2273 3641
rect 2526 3638 2534 3641
rect 2782 3638 2798 3641
rect 3074 3638 3097 3641
rect 3947 3638 3950 3642
rect 2214 3628 2217 3638
rect 3333 3618 3334 3622
rect 3749 3618 3750 3622
rect 4330 3618 4331 3622
rect 496 3603 498 3607
rect 502 3603 505 3607
rect 509 3603 512 3607
rect 1520 3603 1522 3607
rect 1526 3603 1529 3607
rect 1533 3603 1536 3607
rect 2544 3603 2546 3607
rect 2550 3603 2553 3607
rect 2557 3603 2560 3607
rect 3568 3603 3570 3607
rect 3574 3603 3577 3607
rect 3581 3603 3584 3607
rect 1890 3588 1891 3592
rect 1986 3588 1987 3592
rect 2021 3588 2022 3592
rect 2114 3588 2115 3592
rect 1922 3578 1923 3582
rect 2882 3568 2905 3571
rect 3382 3568 3393 3571
rect 3741 3568 3742 3572
rect 3390 3562 3393 3568
rect 3870 3566 3874 3568
rect 538 3558 545 3561
rect 1386 3558 1393 3561
rect 70 3548 94 3551
rect 22 3541 25 3548
rect 346 3548 353 3551
rect 462 3548 473 3551
rect 750 3548 774 3551
rect 830 3548 846 3551
rect 1286 3551 1290 3553
rect 1278 3548 1290 3551
rect 1430 3548 1438 3551
rect 1862 3551 1865 3558
rect 1854 3548 1865 3551
rect 1870 3548 1889 3551
rect 1934 3551 1937 3561
rect 2146 3558 2150 3562
rect 2158 3552 2161 3561
rect 2766 3558 2774 3561
rect 2830 3558 2841 3561
rect 2870 3558 2889 3561
rect 2926 3558 2937 3561
rect 2974 3558 2985 3561
rect 3374 3552 3377 3561
rect 3398 3552 3401 3561
rect 1934 3548 1953 3551
rect 2058 3548 2065 3551
rect 2130 3548 2145 3551
rect 14 3538 25 3541
rect 398 3538 406 3541
rect 430 3538 457 3541
rect 498 3538 521 3541
rect 958 3538 966 3541
rect 1030 3538 1038 3541
rect 1202 3538 1203 3542
rect 1250 3538 1257 3541
rect 1562 3538 1569 3541
rect 2090 3538 2105 3541
rect 2166 3541 2169 3548
rect 2794 3548 2801 3551
rect 2166 3538 2177 3541
rect 2554 3538 2569 3541
rect 2574 3538 2585 3541
rect 2614 3538 2625 3541
rect 2662 3538 2681 3541
rect 2710 3538 2721 3541
rect 2742 3538 2753 3541
rect 2798 3538 2801 3548
rect 3030 3538 3041 3541
rect 3050 3538 3073 3541
rect 3102 3538 3110 3541
rect 3150 3541 3153 3548
rect 4206 3548 4225 3551
rect 4542 3551 4545 3561
rect 4526 3548 4545 3551
rect 4558 3548 4566 3551
rect 3150 3538 3161 3541
rect 3178 3538 3185 3541
rect 3206 3538 3217 3541
rect 3262 3538 3273 3541
rect 3290 3538 3297 3541
rect 3442 3538 3449 3541
rect 3478 3538 3489 3541
rect 3750 3538 3761 3541
rect 4042 3538 4043 3542
rect 410 3528 417 3531
rect 1862 3528 1865 3538
rect 2050 3528 2057 3531
rect 2542 3528 2558 3531
rect 2566 3528 2569 3538
rect 2726 3528 2737 3531
rect 3046 3528 3062 3531
rect 3166 3528 3177 3531
rect 4190 3531 4194 3533
rect 4334 3532 4338 3533
rect 4190 3528 4201 3531
rect 30 3518 46 3521
rect 2301 3518 2302 3522
rect 2594 3518 2595 3522
rect 2762 3518 2763 3522
rect 2908 3518 2910 3522
rect 3197 3518 3198 3522
rect 4078 3518 4094 3521
rect 1000 3503 1002 3507
rect 1006 3503 1009 3507
rect 1013 3503 1016 3507
rect 2024 3503 2026 3507
rect 2030 3503 2033 3507
rect 2037 3503 2040 3507
rect 3048 3503 3050 3507
rect 3054 3503 3057 3507
rect 3061 3503 3064 3507
rect 4080 3503 4082 3507
rect 4086 3503 4089 3507
rect 4093 3503 4096 3507
rect 2580 3488 2582 3492
rect 3386 3488 3387 3492
rect 3429 3488 3430 3492
rect 3254 3478 3265 3481
rect 14 3468 22 3471
rect 154 3468 161 3471
rect 262 3468 286 3471
rect 382 3468 409 3471
rect 1262 3468 1270 3471
rect 1486 3468 1494 3471
rect 1898 3468 1905 3471
rect 2022 3468 2038 3471
rect 2298 3468 2305 3471
rect 2340 3468 2342 3472
rect 2426 3468 2433 3471
rect 3012 3468 3014 3472
rect 3030 3471 3034 3472
rect 3038 3471 3041 3478
rect 4286 3472 4290 3474
rect 3030 3468 3041 3471
rect 3058 3468 3073 3471
rect 3266 3468 3273 3471
rect 3466 3468 3473 3471
rect 3494 3468 3505 3471
rect 3542 3468 3577 3471
rect 3758 3468 3769 3471
rect 3894 3468 3905 3471
rect 4114 3468 4129 3471
rect 4398 3471 4401 3481
rect 4406 3478 4417 3481
rect 4478 3471 4481 3481
rect 4386 3468 4401 3471
rect 4462 3468 4473 3471
rect 4478 3468 4486 3471
rect 4566 3471 4569 3481
rect 4562 3468 4569 3471
rect 54 3458 78 3461
rect 206 3458 214 3461
rect 1270 3458 1282 3461
rect 1390 3458 1409 3461
rect 2002 3458 2009 3461
rect 2034 3458 2065 3461
rect 2142 3458 2150 3461
rect 2294 3458 2310 3461
rect 2454 3458 2470 3461
rect 2518 3458 2529 3461
rect 2626 3458 2633 3461
rect 3454 3458 3473 3461
rect 3578 3458 3585 3461
rect 3590 3458 3598 3461
rect 3782 3458 3790 3461
rect 4310 3458 4337 3461
rect 4354 3458 4361 3461
rect 4502 3461 4505 3468
rect 4494 3458 4505 3461
rect 4570 3458 4577 3461
rect 1278 3457 1282 3458
rect 478 3448 486 3451
rect 2174 3448 2182 3451
rect 2294 3448 2297 3458
rect 2454 3448 2457 3458
rect 2526 3452 2529 3458
rect 2534 3448 2561 3451
rect 3338 3448 3345 3451
rect 3418 3448 3425 3451
rect 3470 3448 3473 3458
rect 3726 3448 3729 3458
rect 3734 3448 3742 3451
rect 3882 3448 3886 3452
rect 450 3438 457 3441
rect 822 3438 830 3441
rect 1298 3438 1301 3442
rect 2678 3438 2686 3441
rect 2878 3441 2881 3448
rect 3534 3442 3538 3444
rect 2870 3438 2881 3441
rect 3002 3438 3009 3441
rect 3198 3438 3206 3441
rect 3522 3438 3529 3441
rect 2966 3428 2969 3438
rect 496 3403 498 3407
rect 502 3403 505 3407
rect 509 3403 512 3407
rect 1520 3403 1522 3407
rect 1526 3403 1529 3407
rect 1533 3403 1536 3407
rect 2544 3403 2546 3407
rect 2550 3403 2553 3407
rect 2557 3403 2560 3407
rect 3568 3403 3570 3407
rect 3574 3403 3577 3407
rect 3581 3403 3584 3407
rect 1941 3388 1942 3392
rect 2165 3388 2166 3392
rect 2194 3388 2195 3392
rect 2242 3388 2243 3392
rect 3038 3388 3046 3391
rect 2117 3378 2118 3382
rect 2782 3366 2786 3368
rect 2998 3366 3002 3368
rect 3358 3366 3362 3368
rect 3506 3368 3514 3371
rect 42 3357 44 3361
rect 1798 3358 1806 3361
rect 2058 3358 2073 3361
rect 2102 3352 2105 3361
rect 2650 3358 2657 3361
rect 2726 3358 2737 3361
rect 2862 3358 2873 3361
rect 3278 3358 3286 3361
rect 3478 3361 3481 3368
rect 3486 3366 3490 3368
rect 3510 3366 3514 3368
rect 3742 3366 3746 3368
rect 3462 3352 3465 3361
rect 3470 3358 3481 3361
rect 3530 3358 3537 3361
rect 3554 3358 3561 3361
rect 4574 3358 4590 3361
rect 4454 3352 4458 3353
rect 54 3348 62 3351
rect 574 3348 593 3351
rect 622 3348 641 3351
rect 670 3348 689 3351
rect 850 3348 857 3351
rect 946 3348 953 3351
rect 1350 3348 1369 3351
rect 1598 3348 1606 3351
rect 1654 3348 1662 3351
rect 1686 3348 1694 3351
rect 1942 3348 1950 3351
rect 2222 3348 2241 3351
rect 2470 3348 2481 3351
rect 2502 3348 2510 3351
rect 3330 3348 3337 3351
rect 2478 3342 2481 3348
rect 14 3338 22 3341
rect 326 3338 334 3341
rect 406 3338 414 3341
rect 1506 3338 1537 3341
rect 1594 3338 1617 3341
rect 2290 3338 2297 3341
rect 2322 3338 2329 3341
rect 2646 3338 2654 3341
rect 2670 3338 2678 3341
rect 2978 3338 2985 3341
rect 3022 3338 3030 3341
rect 3078 3338 3086 3341
rect 3206 3338 3225 3341
rect 3334 3338 3337 3348
rect 3434 3338 3441 3341
rect 3646 3341 3649 3348
rect 3866 3348 3873 3351
rect 3606 3338 3617 3341
rect 3646 3338 3657 3341
rect 3702 3338 3713 3341
rect 3854 3338 3865 3341
rect 4418 3338 4419 3342
rect 3830 3336 3834 3338
rect 4070 3336 4074 3338
rect 254 3332 258 3336
rect 1382 3331 1386 3333
rect 1814 3331 1818 3333
rect 4270 3332 4274 3336
rect 1374 3328 1386 3331
rect 1806 3328 1818 3331
rect 2714 3328 2721 3331
rect 3493 3318 3494 3322
rect 3517 3318 3518 3322
rect 3541 3318 3542 3322
rect 4498 3318 4499 3322
rect 4546 3318 4547 3322
rect 4570 3318 4571 3322
rect 1000 3303 1002 3307
rect 1006 3303 1009 3307
rect 1013 3303 1016 3307
rect 2024 3303 2026 3307
rect 2030 3303 2033 3307
rect 2037 3303 2040 3307
rect 3048 3303 3050 3307
rect 3054 3303 3057 3307
rect 3061 3303 3064 3307
rect 4080 3303 4082 3307
rect 4086 3303 4089 3307
rect 4093 3303 4096 3307
rect 293 3288 294 3292
rect 429 3288 430 3292
rect 1014 3288 1030 3291
rect 2389 3288 2390 3292
rect 2634 3288 2635 3292
rect 2658 3288 2659 3292
rect 2682 3288 2683 3292
rect 2701 3288 2702 3292
rect 2818 3288 2819 3292
rect 2909 3288 2910 3292
rect 3290 3288 3291 3292
rect 3314 3288 3315 3292
rect 3333 3288 3334 3292
rect 190 3278 201 3281
rect 330 3278 334 3282
rect 390 3278 401 3281
rect 190 3277 194 3278
rect 398 3272 401 3278
rect 222 3268 230 3271
rect 270 3268 286 3271
rect 306 3268 321 3271
rect 346 3268 353 3271
rect 462 3271 465 3278
rect 1478 3272 1481 3281
rect 1718 3278 1730 3281
rect 1726 3277 1730 3278
rect 2562 3278 2577 3281
rect 438 3268 457 3271
rect 462 3268 481 3271
rect 1494 3268 1502 3271
rect 1974 3268 1993 3271
rect 2062 3268 2065 3278
rect 3862 3277 3866 3278
rect 3958 3278 3969 3281
rect 4370 3278 4386 3281
rect 3958 3277 3962 3278
rect 4382 3274 4386 3278
rect 2454 3268 2465 3271
rect 2482 3268 2489 3271
rect 2506 3268 2513 3271
rect 2550 3268 2558 3271
rect 2582 3268 2593 3271
rect 206 3258 214 3261
rect 586 3258 593 3261
rect 682 3258 689 3261
rect 1358 3258 1366 3261
rect 1466 3258 1473 3261
rect 1942 3258 1961 3261
rect 1966 3258 1982 3261
rect 2006 3258 2014 3261
rect 2462 3262 2465 3268
rect 2614 3262 2617 3271
rect 2718 3268 2729 3271
rect 2770 3268 2785 3271
rect 3102 3268 3113 3271
rect 3178 3268 3185 3271
rect 3206 3268 3217 3271
rect 3270 3268 3278 3271
rect 3346 3268 3353 3271
rect 3374 3268 3385 3271
rect 3422 3268 3433 3271
rect 3566 3268 3593 3271
rect 3726 3268 3737 3271
rect 4094 3268 4102 3271
rect 4106 3268 4110 3271
rect 4542 3268 4553 3271
rect 2718 3262 2721 3268
rect 2422 3258 2438 3261
rect 2982 3258 2993 3261
rect 3166 3258 3185 3261
rect 3414 3258 3422 3261
rect 3558 3258 3566 3261
rect 3974 3258 3993 3261
rect 4018 3258 4025 3261
rect 4262 3258 4289 3261
rect 4554 3258 4561 3261
rect 734 3248 745 3251
rect 1426 3248 1433 3251
rect 1942 3248 1945 3258
rect 2422 3248 2425 3258
rect 2990 3252 2993 3258
rect 2526 3248 2534 3251
rect 2898 3248 2905 3251
rect 3102 3248 3110 3251
rect 3182 3248 3185 3258
rect 3322 3248 3329 3251
rect 4258 3248 4262 3252
rect 1710 3238 1718 3241
rect 2410 3238 2417 3241
rect 3939 3238 3942 3242
rect 4187 3238 4190 3242
rect 786 3228 787 3232
rect 410 3218 411 3222
rect 3557 3218 3558 3222
rect 496 3203 498 3207
rect 502 3203 505 3207
rect 509 3203 512 3207
rect 1520 3203 1522 3207
rect 1526 3203 1529 3207
rect 1533 3203 1536 3207
rect 2544 3203 2546 3207
rect 2550 3203 2553 3207
rect 2557 3203 2560 3207
rect 3568 3203 3570 3207
rect 3574 3203 3577 3207
rect 3581 3203 3584 3207
rect 2170 3188 2171 3192
rect 2218 3188 2219 3192
rect 2365 3188 2366 3192
rect 4069 3178 4070 3182
rect 1838 3168 1846 3171
rect 2070 3168 2078 3171
rect 3254 3168 3266 3171
rect 198 3161 201 3168
rect 3254 3162 3257 3168
rect 3262 3166 3266 3168
rect 190 3158 201 3161
rect 2082 3158 2089 3161
rect 10 3148 17 3151
rect 58 3148 65 3151
rect 414 3148 422 3151
rect 478 3148 489 3151
rect 486 3142 489 3148
rect 1170 3148 1177 3151
rect 110 3138 118 3141
rect 438 3138 465 3141
rect 498 3138 505 3141
rect 1034 3138 1049 3141
rect 1206 3138 1218 3141
rect 1342 3141 1345 3151
rect 1430 3148 1438 3151
rect 1470 3148 1478 3151
rect 1530 3148 1545 3151
rect 1654 3148 1662 3151
rect 1678 3148 1686 3151
rect 1710 3148 1718 3151
rect 1726 3148 1734 3151
rect 2098 3148 2105 3151
rect 2118 3151 2121 3161
rect 2250 3158 2254 3162
rect 2118 3148 2137 3151
rect 2198 3148 2217 3151
rect 2350 3151 2353 3161
rect 2938 3158 2945 3161
rect 3062 3158 3070 3161
rect 3278 3161 3281 3168
rect 3646 3166 3650 3168
rect 3278 3158 3289 3161
rect 2322 3148 2329 3151
rect 2334 3148 2353 3151
rect 2622 3151 2625 3158
rect 2622 3148 2641 3151
rect 3118 3148 3137 3151
rect 3334 3151 3337 3161
rect 3682 3158 3686 3162
rect 4046 3158 4057 3161
rect 4582 3158 4590 3161
rect 4046 3156 4050 3158
rect 4262 3156 4266 3158
rect 3318 3148 3337 3151
rect 1342 3138 1361 3141
rect 1442 3138 1457 3141
rect 1518 3138 1534 3141
rect 1586 3138 1593 3141
rect 1618 3138 1633 3141
rect 2378 3138 2385 3141
rect 2554 3138 2574 3141
rect 2854 3138 2862 3141
rect 2958 3138 2977 3141
rect 3134 3138 3137 3148
rect 3750 3148 3758 3151
rect 3278 3138 3286 3141
rect 3382 3138 3393 3141
rect 3694 3138 3705 3141
rect 3726 3138 3737 3141
rect 3854 3138 3866 3141
rect 4294 3138 4297 3148
rect 4538 3148 4545 3151
rect 4390 3138 4401 3141
rect 4486 3141 4489 3148
rect 4486 3138 4497 3141
rect 4542 3138 4545 3148
rect 166 3128 174 3131
rect 1742 3131 1746 3133
rect 1854 3131 1858 3133
rect 2678 3132 2681 3138
rect 4046 3136 4050 3138
rect 4390 3136 4394 3138
rect 1734 3128 1746 3131
rect 1846 3128 1858 3131
rect 2678 3128 2686 3132
rect 3062 3118 3070 3121
rect 3269 3118 3270 3122
rect 3293 3118 3294 3122
rect 3653 3118 3654 3122
rect 4578 3118 4579 3122
rect 1000 3103 1002 3107
rect 1006 3103 1009 3107
rect 1013 3103 1016 3107
rect 2024 3103 2026 3107
rect 2030 3103 2033 3107
rect 2037 3103 2040 3107
rect 3048 3103 3050 3107
rect 3054 3103 3057 3107
rect 3061 3103 3064 3107
rect 4080 3103 4082 3107
rect 4086 3103 4089 3107
rect 4093 3103 4096 3107
rect 365 3088 366 3092
rect 494 3088 510 3091
rect 634 3088 635 3092
rect 2498 3088 2499 3092
rect 2757 3088 2758 3092
rect 2893 3088 2894 3092
rect 3034 3088 3035 3092
rect 3098 3088 3099 3092
rect 4450 3088 4451 3092
rect 6 3072 9 3081
rect 30 3071 34 3072
rect 38 3071 41 3078
rect 246 3072 249 3081
rect 434 3078 441 3081
rect 30 3068 41 3071
rect 470 3071 473 3078
rect 1454 3072 1457 3081
rect 1502 3078 1518 3081
rect 1726 3072 1729 3078
rect 2678 3072 2681 3081
rect 4110 3081 4113 3088
rect 4094 3078 4113 3081
rect 4094 3077 4098 3078
rect 3998 3072 4002 3074
rect 374 3068 385 3071
rect 438 3068 465 3071
rect 470 3068 481 3071
rect 1334 3068 1350 3071
rect 1506 3068 1537 3071
rect 1726 3068 1730 3072
rect 2246 3068 2254 3071
rect 2374 3068 2382 3071
rect 2478 3068 2486 3071
rect 2514 3068 2521 3071
rect 2590 3068 2601 3071
rect 2686 3068 2697 3071
rect 2742 3068 2750 3071
rect 2798 3068 2809 3071
rect 2958 3068 2974 3071
rect 3042 3068 3057 3071
rect 3118 3068 3137 3071
rect 3278 3068 3297 3071
rect 3458 3068 3465 3071
rect 3550 3068 3561 3071
rect 3586 3068 3594 3071
rect 3702 3068 3710 3071
rect 3902 3068 3914 3071
rect 4270 3071 4274 3074
rect 4270 3068 4281 3071
rect 4354 3068 4361 3071
rect 4494 3068 4505 3071
rect 10 3058 17 3061
rect 254 3058 262 3061
rect 678 3058 697 3061
rect 710 3058 737 3061
rect 774 3061 777 3068
rect 774 3058 793 3061
rect 838 3058 846 3061
rect 1334 3058 1337 3068
rect 1430 3058 1449 3061
rect 1478 3058 1497 3061
rect 1582 3058 1590 3061
rect 2598 3062 2601 3068
rect 2110 3058 2129 3061
rect 2314 3058 2329 3061
rect 2342 3058 2361 3061
rect 2370 3058 2393 3061
rect 2418 3058 2425 3061
rect 2446 3058 2462 3061
rect 2542 3058 2574 3061
rect 2646 3058 2654 3061
rect 2718 3058 2737 3061
rect 3298 3058 3305 3061
rect 3486 3058 3494 3061
rect 3530 3058 3537 3061
rect 3866 3058 3873 3061
rect 4142 3058 4161 3061
rect 4166 3058 4174 3061
rect 4278 3062 4281 3068
rect 4310 3058 4329 3061
rect 4342 3058 4350 3061
rect 4438 3061 4441 3068
rect 4362 3058 4369 3061
rect 4430 3058 4441 3061
rect 326 3051 329 3058
rect 318 3048 329 3051
rect 354 3048 361 3051
rect 382 3048 390 3051
rect 702 3051 705 3058
rect 694 3048 705 3051
rect 766 3048 774 3051
rect 2126 3048 2129 3058
rect 2202 3048 2206 3052
rect 2298 3048 2302 3052
rect 2342 3048 2345 3058
rect 2446 3048 2449 3058
rect 2502 3048 2510 3051
rect 2542 3048 2545 3058
rect 2718 3048 2721 3058
rect 3102 3048 3110 3051
rect 3262 3048 3273 3051
rect 3510 3048 3529 3051
rect 4142 3048 4145 3058
rect 4282 3048 4289 3051
rect 4326 3048 4329 3058
rect 3270 3042 3273 3048
rect 674 3038 675 3042
rect 3787 3038 3790 3042
rect 3306 3018 3307 3022
rect 3485 3018 3486 3022
rect 496 3003 498 3007
rect 502 3003 505 3007
rect 509 3003 512 3007
rect 1520 3003 1522 3007
rect 1526 3003 1529 3007
rect 1533 3003 1536 3007
rect 2544 3003 2546 3007
rect 2550 3003 2553 3007
rect 2557 3003 2560 3007
rect 3568 3003 3570 3007
rect 3574 3003 3577 3007
rect 3581 3003 3584 3007
rect 2565 2988 2566 2992
rect 2733 2988 2734 2992
rect 2914 2988 2915 2992
rect 3229 2988 3230 2992
rect 4078 2988 4094 2991
rect 1874 2968 1877 2972
rect 1970 2968 1973 2972
rect 1014 2966 1018 2968
rect 2470 2966 2474 2968
rect 2614 2968 2622 2971
rect 2614 2966 2618 2968
rect 2638 2966 2642 2968
rect 2646 2966 2650 2968
rect 2694 2966 2698 2968
rect 2838 2966 2842 2968
rect 2878 2968 2886 2971
rect 2954 2968 2962 2971
rect 3058 2968 3074 2971
rect 2878 2966 2882 2968
rect 2958 2966 2962 2968
rect 3070 2966 3074 2968
rect 3094 2966 3098 2968
rect 3138 2968 3146 2971
rect 3118 2966 3122 2968
rect 3142 2966 3146 2968
rect 3182 2966 3186 2968
rect 3206 2966 3210 2968
rect 3262 2966 3266 2968
rect 3290 2968 3298 2971
rect 4562 2968 4577 2971
rect 3270 2966 3274 2968
rect 3294 2966 3298 2968
rect 518 2951 521 2961
rect 530 2958 534 2962
rect 558 2958 577 2961
rect 486 2948 521 2951
rect 742 2948 753 2951
rect 742 2941 745 2948
rect 1438 2948 1457 2951
rect 2470 2951 2473 2961
rect 2546 2958 2553 2961
rect 2666 2958 2673 2961
rect 2810 2958 2817 2961
rect 2458 2948 2465 2951
rect 2470 2948 2486 2951
rect 2494 2948 2510 2951
rect 2758 2948 2777 2951
rect 2782 2948 2790 2951
rect 2926 2951 2929 2961
rect 2978 2958 2985 2961
rect 3854 2952 3857 2961
rect 2926 2948 2945 2951
rect 2758 2942 2761 2948
rect 738 2938 745 2941
rect 754 2938 761 2941
rect 1042 2938 1049 2941
rect 1386 2938 1393 2941
rect 2058 2938 2065 2941
rect 2526 2938 2534 2941
rect 2574 2938 2585 2941
rect 2742 2938 2753 2941
rect 2790 2938 2801 2941
rect 2854 2938 2862 2941
rect 2894 2938 2905 2941
rect 2950 2938 2958 2941
rect 2982 2941 2985 2948
rect 3922 2948 3937 2951
rect 2982 2938 2993 2941
rect 3046 2938 3070 2941
rect 3110 2938 3118 2941
rect 3326 2938 3337 2941
rect 3670 2938 3681 2941
rect 3734 2938 3745 2941
rect 3966 2938 3978 2941
rect 4270 2941 4273 2948
rect 4490 2948 4497 2951
rect 4262 2938 4273 2941
rect 4310 2938 4318 2941
rect 4478 2938 4489 2941
rect 4542 2938 4550 2941
rect 1070 2931 1073 2938
rect 1010 2928 1041 2931
rect 1062 2928 1073 2931
rect 1598 2931 1602 2933
rect 2510 2932 2513 2938
rect 1590 2928 1602 2931
rect 2510 2928 2518 2932
rect 2806 2928 2809 2938
rect 3030 2932 3033 2938
rect 4262 2936 4266 2938
rect 3030 2928 3038 2932
rect 4062 2931 4066 2933
rect 4262 2931 4266 2933
rect 4462 2932 4466 2933
rect 4062 2928 4073 2931
rect 4262 2928 4273 2931
rect 2653 2918 2654 2922
rect 2845 2918 2846 2922
rect 2874 2918 2875 2922
rect 2965 2918 2966 2922
rect 3077 2918 3078 2922
rect 3101 2918 3102 2922
rect 3149 2918 3150 2922
rect 3277 2918 3278 2922
rect 3301 2918 3302 2922
rect 1000 2903 1002 2907
rect 1006 2903 1009 2907
rect 1013 2903 1016 2907
rect 2024 2903 2026 2907
rect 2030 2903 2033 2907
rect 2037 2903 2040 2907
rect 3048 2903 3050 2907
rect 3054 2903 3057 2907
rect 3061 2903 3064 2907
rect 4080 2903 4082 2907
rect 4086 2903 4089 2907
rect 4093 2903 4096 2907
rect 494 2888 510 2891
rect 974 2888 982 2891
rect 2541 2888 2542 2892
rect 2722 2888 2723 2892
rect 2906 2888 2907 2892
rect 3237 2888 3238 2892
rect 14 2878 22 2881
rect 70 2878 78 2881
rect 150 2878 158 2881
rect 310 2878 318 2881
rect 94 2868 102 2871
rect 302 2868 329 2871
rect 470 2871 473 2881
rect 830 2878 846 2881
rect 918 2872 921 2881
rect 1822 2872 1825 2881
rect 2630 2872 2633 2881
rect 3318 2872 3321 2881
rect 4142 2877 4146 2878
rect 470 2868 478 2871
rect 498 2868 529 2871
rect 854 2868 873 2871
rect 1133 2868 1134 2872
rect 1182 2868 1194 2871
rect 1830 2868 1838 2871
rect 2550 2868 2561 2871
rect 2570 2868 2585 2871
rect 2638 2868 2649 2871
rect 2682 2868 2689 2871
rect 2726 2868 2737 2871
rect 2754 2868 2761 2871
rect 2778 2868 2793 2871
rect 2830 2868 2838 2871
rect 2870 2868 2881 2871
rect 2890 2868 2897 2871
rect 2914 2868 2929 2871
rect 2974 2868 2993 2871
rect 3078 2868 3089 2871
rect 3158 2868 3169 2871
rect 3214 2868 3222 2871
rect 3302 2868 3313 2871
rect 3462 2868 3473 2871
rect 3534 2868 3545 2871
rect 3694 2868 3705 2871
rect 3714 2868 3721 2871
rect 394 2858 401 2861
rect 446 2858 457 2861
rect 606 2858 630 2861
rect 926 2858 937 2861
rect 1618 2858 1625 2861
rect 1798 2858 1817 2861
rect 2470 2858 2478 2861
rect 2558 2861 2561 2868
rect 2726 2862 2729 2868
rect 2558 2858 2574 2861
rect 3110 2858 3118 2861
rect 3194 2858 3201 2861
rect 3262 2858 3281 2861
rect 3686 2858 3694 2861
rect 3846 2862 3849 2871
rect 3870 2868 3881 2871
rect 3902 2868 3913 2871
rect 4414 2868 4422 2871
rect 4518 2871 4522 2874
rect 4518 2868 4529 2871
rect 4586 2868 4593 2871
rect 4482 2858 4489 2861
rect 4534 2858 4554 2861
rect 122 2849 124 2853
rect 282 2849 284 2853
rect 598 2848 609 2851
rect 2610 2848 2617 2851
rect 2750 2848 2758 2851
rect 3110 2848 3113 2858
rect 3278 2848 3281 2858
rect 4550 2856 4554 2858
rect 3482 2848 3489 2851
rect 3494 2848 3505 2851
rect 3502 2842 3505 2848
rect 2266 2838 2269 2842
rect 4011 2838 4014 2842
rect 3098 2818 3099 2822
rect 3178 2818 3179 2822
rect 3453 2818 3454 2822
rect 3685 2818 3686 2822
rect 3922 2818 3923 2822
rect 496 2803 498 2807
rect 502 2803 505 2807
rect 509 2803 512 2807
rect 1520 2803 1522 2807
rect 1526 2803 1529 2807
rect 1533 2803 1536 2807
rect 2544 2803 2546 2807
rect 2550 2803 2553 2807
rect 2557 2803 2560 2807
rect 3568 2803 3570 2807
rect 3574 2803 3577 2807
rect 3581 2803 3584 2807
rect 974 2788 990 2791
rect 3077 2788 3078 2792
rect 1930 2768 1933 2772
rect 2358 2766 2362 2768
rect 2382 2766 2386 2768
rect 2406 2766 2410 2768
rect 2430 2768 2438 2771
rect 2430 2766 2434 2768
rect 2734 2766 2738 2768
rect 2774 2766 2778 2768
rect 2814 2768 2822 2771
rect 2814 2766 2818 2768
rect 2838 2766 2842 2768
rect 2910 2768 2918 2771
rect 3723 2768 3726 2772
rect 4075 2768 4078 2772
rect 2910 2766 2914 2768
rect 350 2756 354 2758
rect 30 2748 38 2751
rect 70 2748 102 2751
rect 22 2741 25 2748
rect 294 2748 302 2751
rect 390 2748 398 2751
rect 1222 2748 1238 2751
rect 1630 2751 1634 2753
rect 1622 2748 1634 2751
rect 1682 2748 1689 2751
rect 1838 2748 1846 2751
rect 1854 2748 1873 2751
rect 2126 2748 2134 2751
rect 2302 2751 2305 2761
rect 3106 2758 3113 2761
rect 3646 2756 3650 2758
rect 2302 2748 2318 2751
rect 2946 2748 2953 2751
rect 2998 2748 3017 2751
rect 3038 2748 3046 2751
rect 3226 2748 3233 2751
rect 3238 2748 3246 2751
rect 3014 2742 3017 2748
rect 3766 2748 3785 2751
rect 3814 2748 3833 2751
rect 3950 2748 3961 2751
rect 4334 2748 4345 2751
rect 4466 2748 4473 2751
rect 14 2738 25 2741
rect 446 2738 457 2741
rect 1594 2738 1601 2741
rect 1730 2738 1737 2741
rect 1762 2738 1777 2741
rect 1810 2738 1817 2741
rect 2294 2738 2302 2741
rect 2446 2738 2457 2741
rect 2582 2738 2593 2741
rect 2630 2738 2641 2741
rect 2678 2738 2689 2741
rect 2746 2738 2753 2741
rect 2790 2738 2798 2741
rect 2870 2738 2881 2741
rect 2966 2738 2977 2741
rect 3086 2738 3097 2741
rect 3134 2738 3145 2741
rect 3166 2738 3177 2741
rect 3214 2738 3225 2741
rect 3374 2738 3385 2741
rect 3422 2738 3433 2741
rect 3974 2738 3982 2741
rect 4302 2741 4305 2748
rect 4294 2738 4305 2741
rect 4314 2738 4321 2741
rect 4366 2738 4385 2741
rect 4502 2738 4514 2741
rect 6 2728 9 2738
rect 446 2736 450 2738
rect 502 2736 506 2738
rect 150 2728 158 2731
rect 3974 2728 3977 2738
rect 470 2718 486 2721
rect 2354 2718 2355 2722
rect 2378 2718 2379 2722
rect 2402 2718 2403 2722
rect 2730 2718 2731 2722
rect 2810 2718 2811 2722
rect 2834 2718 2835 2722
rect 2906 2718 2907 2722
rect 3534 2718 3550 2721
rect 3989 2718 3990 2722
rect 1000 2703 1002 2707
rect 1006 2703 1009 2707
rect 1013 2703 1016 2707
rect 2024 2703 2026 2707
rect 2030 2703 2033 2707
rect 2037 2703 2040 2707
rect 3048 2703 3050 2707
rect 3054 2703 3057 2707
rect 3061 2703 3064 2707
rect 4080 2703 4082 2707
rect 4086 2703 4089 2707
rect 4093 2703 4096 2707
rect 1674 2688 1675 2692
rect 150 2678 158 2681
rect 638 2678 646 2681
rect 1654 2672 1657 2681
rect 1902 2678 1914 2681
rect 2754 2678 2770 2681
rect 1910 2677 1914 2678
rect 2766 2674 2770 2678
rect 3030 2672 3033 2681
rect 4422 2672 4426 2674
rect 30 2668 38 2671
rect 150 2668 177 2671
rect 1578 2668 1585 2671
rect 1686 2668 1694 2671
rect 2222 2668 2233 2671
rect 2270 2668 2281 2671
rect 2318 2668 2329 2671
rect 2574 2668 2582 2671
rect 2910 2668 2921 2671
rect 2954 2668 2969 2671
rect 3014 2668 3025 2671
rect 3062 2668 3089 2671
rect 150 2661 153 2668
rect 138 2658 153 2661
rect 674 2658 681 2661
rect 1310 2658 1326 2661
rect 1642 2658 1649 2661
rect 3198 2662 3201 2671
rect 3222 2668 3241 2671
rect 3386 2668 3393 2671
rect 3950 2668 3977 2671
rect 3990 2668 4009 2671
rect 4134 2668 4153 2671
rect 4502 2668 4514 2671
rect 3054 2658 3078 2661
rect 3374 2658 3382 2661
rect 3446 2658 3462 2661
rect 3638 2658 3657 2661
rect 3686 2658 3705 2661
rect 3914 2658 3921 2661
rect 4070 2658 4105 2661
rect 4214 2658 4217 2668
rect 4238 2658 4257 2661
rect 4270 2658 4278 2661
rect 4458 2658 4473 2661
rect 4542 2658 4558 2661
rect 2806 2652 2810 2657
rect 4054 2651 4057 2658
rect 4046 2648 4057 2651
rect 4070 2652 4073 2658
rect 4118 2648 4137 2651
rect 1539 2638 1542 2642
rect 3315 2638 3318 2642
rect 3394 2638 3401 2641
rect 2242 2628 2243 2632
rect 493 2618 494 2622
rect 2290 2618 2291 2622
rect 2901 2618 2902 2622
rect 3922 2618 3923 2622
rect 4106 2618 4107 2622
rect 4290 2618 4291 2622
rect 496 2603 498 2607
rect 502 2603 505 2607
rect 509 2603 512 2607
rect 1520 2603 1522 2607
rect 1526 2603 1529 2607
rect 1533 2603 1536 2607
rect 2544 2603 2546 2607
rect 2550 2603 2553 2607
rect 2557 2603 2560 2607
rect 3568 2603 3570 2607
rect 3574 2603 3577 2607
rect 3581 2603 3584 2607
rect 2237 2588 2238 2592
rect 3010 2588 3011 2592
rect 3154 2588 3155 2592
rect 4122 2588 4123 2592
rect 1902 2568 1910 2571
rect 1902 2566 1906 2568
rect 1926 2566 1930 2568
rect 1998 2568 2006 2571
rect 1998 2566 2002 2568
rect 2110 2566 2114 2568
rect 2166 2568 2174 2571
rect 2190 2568 2198 2571
rect 2286 2568 2294 2571
rect 2869 2568 2870 2572
rect 3586 2568 3593 2571
rect 2166 2566 2170 2568
rect 2190 2566 2194 2568
rect 2286 2566 2290 2568
rect 2950 2566 2954 2568
rect 3838 2566 3842 2568
rect 58 2557 60 2561
rect 22 2541 25 2548
rect 494 2548 502 2551
rect 550 2548 558 2551
rect 918 2548 926 2551
rect 1390 2548 1406 2551
rect 2222 2551 2225 2561
rect 2426 2558 2433 2561
rect 2206 2548 2225 2551
rect 2438 2551 2441 2561
rect 2438 2548 2446 2551
rect 2450 2548 2457 2551
rect 2462 2548 2470 2551
rect 2870 2548 2878 2551
rect 2990 2551 2993 2561
rect 3710 2558 3721 2561
rect 3830 2558 3841 2561
rect 2990 2548 3006 2551
rect 3302 2548 3310 2551
rect 14 2538 25 2541
rect 774 2538 782 2541
rect 1034 2538 1050 2541
rect 1282 2538 1289 2541
rect 1966 2538 1974 2541
rect 2018 2538 2025 2541
rect 2122 2538 2129 2541
rect 2246 2538 2257 2541
rect 2614 2538 2625 2541
rect 2646 2538 2657 2541
rect 2894 2538 2905 2541
rect 3334 2541 3337 2548
rect 3446 2548 3462 2551
rect 3478 2548 3486 2551
rect 3510 2548 3529 2551
rect 3558 2548 3566 2551
rect 3670 2548 3689 2551
rect 3726 2548 3742 2551
rect 3758 2548 3777 2551
rect 3846 2548 3854 2551
rect 4030 2548 4073 2551
rect 4126 2548 4134 2551
rect 4254 2551 4257 2561
rect 4358 2558 4369 2561
rect 4238 2548 4257 2551
rect 4282 2548 4289 2551
rect 4422 2548 4433 2551
rect 4502 2548 4521 2551
rect 3326 2538 3337 2541
rect 3630 2541 3633 2548
rect 3622 2538 3633 2541
rect 3786 2538 3793 2541
rect 3910 2541 3913 2548
rect 3902 2538 3913 2541
rect 3958 2538 3966 2541
rect 4090 2538 4113 2541
rect 4118 2538 4137 2541
rect 4158 2538 4177 2541
rect 4190 2538 4198 2541
rect 4278 2538 4297 2541
rect 4318 2538 4326 2541
rect 4398 2538 4414 2541
rect 4542 2538 4569 2541
rect 30 2528 38 2531
rect 150 2528 158 2531
rect 534 2531 538 2536
rect 534 2528 550 2531
rect 2342 2531 2346 2536
rect 2342 2528 2358 2531
rect 2494 2531 2498 2536
rect 2494 2528 2510 2531
rect 1898 2518 1899 2522
rect 1994 2518 1995 2522
rect 2106 2518 2107 2522
rect 2282 2518 2283 2522
rect 2586 2518 2593 2521
rect 2886 2518 2889 2531
rect 3062 2531 3066 2536
rect 3062 2528 3078 2531
rect 4110 2528 4113 2538
rect 4410 2528 4417 2531
rect 2946 2518 2947 2522
rect 4018 2518 4023 2522
rect 4530 2518 4531 2522
rect 1000 2503 1002 2507
rect 1006 2503 1009 2507
rect 1013 2503 1016 2507
rect 2024 2503 2026 2507
rect 2030 2503 2033 2507
rect 2037 2503 2040 2507
rect 3048 2503 3050 2507
rect 3054 2503 3057 2507
rect 3061 2503 3064 2507
rect 4080 2503 4082 2507
rect 4086 2503 4089 2507
rect 4093 2503 4096 2507
rect 2034 2488 2049 2491
rect 2749 2488 2750 2492
rect 3037 2488 3038 2492
rect 3202 2488 3203 2492
rect 3602 2488 3603 2492
rect 4098 2488 4105 2491
rect 70 2478 78 2481
rect 1522 2478 1538 2481
rect 2022 2478 2038 2481
rect 2230 2478 2241 2481
rect 3086 2478 3102 2481
rect 3806 2478 3825 2481
rect 1534 2474 1538 2478
rect 3086 2474 3090 2478
rect 14 2468 22 2471
rect 342 2468 369 2471
rect 470 2471 474 2474
rect 2726 2472 2730 2474
rect 2910 2472 2914 2474
rect 3078 2472 3082 2474
rect 470 2468 481 2471
rect 486 2468 529 2471
rect 946 2468 953 2471
rect 974 2468 982 2471
rect 1062 2468 1070 2471
rect 1958 2468 1969 2471
rect 2006 2468 2017 2471
rect 2174 2468 2182 2471
rect 2214 2468 2225 2471
rect 2806 2468 2817 2471
rect 2938 2468 2945 2471
rect 2982 2468 2993 2471
rect 3046 2468 3054 2471
rect 3278 2468 3286 2471
rect 3542 2468 3550 2471
rect 3678 2468 3694 2471
rect 3988 2468 3990 2472
rect 4266 2468 4281 2471
rect 478 2462 481 2468
rect 270 2458 281 2461
rect 334 2458 342 2461
rect 514 2458 537 2461
rect 938 2458 961 2461
rect 1130 2458 1137 2461
rect 1494 2458 1502 2461
rect 1690 2458 1705 2461
rect 2186 2458 2201 2461
rect 2470 2458 2489 2461
rect 2526 2458 2561 2461
rect 2598 2458 2617 2461
rect 2630 2458 2638 2461
rect 2758 2458 2769 2461
rect 2982 2462 2985 2468
rect 2970 2458 2977 2461
rect 3662 2461 3665 2468
rect 3654 2458 3665 2461
rect 3766 2461 3769 2468
rect 3758 2458 3769 2461
rect 3846 2458 3873 2461
rect 3942 2461 3945 2468
rect 3942 2458 3953 2461
rect 4046 2458 4062 2461
rect 4070 2458 4078 2461
rect 4202 2458 4209 2461
rect 4246 2458 4254 2461
rect 4354 2458 4369 2461
rect 4398 2458 4417 2461
rect 4510 2458 4529 2461
rect 4534 2458 4553 2461
rect 4566 2458 4593 2461
rect 270 2457 274 2458
rect 42 2449 44 2453
rect 2486 2448 2489 2458
rect 2558 2448 2561 2458
rect 2614 2448 2617 2458
rect 2758 2452 2761 2458
rect 3022 2448 3030 2451
rect 3346 2448 3353 2451
rect 3646 2451 3649 2458
rect 4414 2452 4417 2458
rect 3606 2448 3617 2451
rect 3638 2448 3649 2451
rect 3758 2448 3769 2451
rect 3774 2448 3782 2451
rect 3886 2448 3897 2451
rect 4382 2448 4401 2451
rect 4550 2448 4553 2458
rect 986 2438 993 2441
rect 3214 2438 3222 2441
rect 3322 2438 3329 2441
rect 4370 2438 4371 2442
rect 4470 2438 4497 2441
rect 1997 2418 1998 2422
rect 2154 2418 2155 2422
rect 4045 2418 4046 2422
rect 4429 2418 4430 2422
rect 4565 2418 4566 2422
rect 496 2403 498 2407
rect 502 2403 505 2407
rect 509 2403 512 2407
rect 1520 2403 1522 2407
rect 1526 2403 1529 2407
rect 1533 2403 1536 2407
rect 2544 2403 2546 2407
rect 2550 2403 2553 2407
rect 2557 2403 2560 2407
rect 3568 2403 3570 2407
rect 3574 2403 3577 2407
rect 3581 2403 3584 2407
rect 3546 2378 3547 2382
rect 1299 2368 1302 2372
rect 1395 2368 1398 2372
rect 2750 2368 2761 2371
rect 2758 2362 2761 2368
rect 4274 2368 4275 2372
rect 4286 2368 4297 2371
rect 4517 2368 4518 2372
rect 4546 2368 4547 2372
rect 1962 2358 1966 2362
rect 906 2348 913 2351
rect 990 2348 998 2351
rect 1598 2348 1606 2351
rect 1706 2348 1721 2351
rect 1966 2348 1974 2351
rect 2114 2348 2121 2351
rect 2226 2348 2233 2351
rect 2270 2348 2289 2351
rect 2390 2348 2398 2351
rect 2422 2351 2425 2361
rect 2406 2348 2425 2351
rect 2438 2348 2457 2351
rect 2646 2348 2654 2351
rect 102 2338 118 2341
rect 582 2338 609 2341
rect 750 2338 761 2341
rect 894 2338 905 2341
rect 1450 2338 1458 2341
rect 1554 2338 1570 2341
rect 1974 2338 1985 2341
rect 2134 2338 2145 2341
rect 2182 2338 2193 2341
rect 2214 2338 2225 2341
rect 2486 2338 2494 2341
rect 2498 2338 2510 2341
rect 2734 2341 2737 2348
rect 2726 2338 2737 2341
rect 2774 2341 2777 2361
rect 2918 2361 2921 2368
rect 2898 2358 2905 2361
rect 2910 2358 2921 2361
rect 3066 2358 3073 2361
rect 2782 2351 2785 2358
rect 2782 2348 2793 2351
rect 2886 2348 2894 2351
rect 2942 2348 2950 2351
rect 2998 2348 3025 2351
rect 3182 2351 3185 2361
rect 3194 2358 3198 2362
rect 3590 2358 3601 2361
rect 3678 2358 3689 2361
rect 4086 2358 4113 2361
rect 4362 2358 4366 2362
rect 3214 2351 3217 2358
rect 3166 2348 3185 2351
rect 3198 2348 3217 2351
rect 3470 2351 3474 2354
rect 3686 2352 3689 2358
rect 3422 2348 3441 2351
rect 3462 2348 3474 2351
rect 3518 2348 3526 2351
rect 3606 2348 3614 2351
rect 3698 2348 3705 2351
rect 3710 2348 3729 2351
rect 3974 2351 3977 2358
rect 3950 2348 3969 2351
rect 3974 2348 3985 2351
rect 4038 2348 4046 2351
rect 4434 2348 4441 2351
rect 4558 2351 4561 2361
rect 4558 2348 4577 2351
rect 2754 2338 2761 2341
rect 2774 2338 2785 2341
rect 3106 2338 3113 2341
rect 3302 2341 3305 2348
rect 3266 2338 3273 2341
rect 3278 2338 3289 2341
rect 3294 2338 3305 2341
rect 3618 2338 3625 2341
rect 3738 2338 3745 2341
rect 3826 2338 3833 2341
rect 3902 2338 3929 2341
rect 4054 2338 4073 2341
rect 4134 2338 4142 2341
rect 4478 2338 4489 2341
rect 158 2328 174 2331
rect 1870 2331 1874 2336
rect 2534 2333 2538 2338
rect 994 2328 1001 2331
rect 1870 2328 1886 2331
rect 2630 2331 2634 2336
rect 2630 2328 2646 2331
rect 2734 2328 2737 2338
rect 2782 2328 2785 2338
rect 3278 2332 3281 2338
rect 3622 2328 3625 2338
rect 2002 2318 2017 2321
rect 2333 2318 2334 2322
rect 4082 2318 4083 2322
rect 4202 2318 4203 2322
rect 1000 2303 1002 2307
rect 1006 2303 1009 2307
rect 1013 2303 1016 2307
rect 2024 2303 2026 2307
rect 2030 2303 2033 2307
rect 2037 2303 2040 2307
rect 3048 2303 3050 2307
rect 3054 2303 3057 2307
rect 3061 2303 3064 2307
rect 4080 2303 4082 2307
rect 4086 2303 4089 2307
rect 4093 2303 4096 2307
rect 2770 2288 2771 2292
rect 3861 2288 3862 2292
rect 4212 2288 4214 2292
rect 178 2278 185 2281
rect 190 2278 198 2281
rect 854 2278 865 2281
rect 966 2278 974 2281
rect 1002 2278 1025 2281
rect 2542 2278 2577 2281
rect 854 2277 858 2278
rect 134 2268 142 2271
rect 374 2268 382 2271
rect 550 2268 577 2271
rect 694 2268 702 2271
rect 910 2268 918 2271
rect 2038 2268 2066 2271
rect 22 2258 34 2261
rect 174 2258 190 2261
rect 1790 2258 1798 2261
rect 2334 2262 2337 2271
rect 2634 2268 2649 2271
rect 2822 2271 2825 2278
rect 2822 2268 2833 2271
rect 2990 2268 2998 2271
rect 3054 2268 3070 2271
rect 3086 2271 3089 2281
rect 3566 2278 3574 2281
rect 3074 2268 3089 2271
rect 3110 2268 3137 2271
rect 3206 2268 3225 2271
rect 3286 2268 3294 2271
rect 3398 2268 3417 2271
rect 3518 2268 3526 2271
rect 3678 2271 3681 2281
rect 3806 2278 3814 2281
rect 3662 2268 3681 2271
rect 3918 2271 3921 2281
rect 3766 2268 3785 2271
rect 3870 2268 3889 2271
rect 3902 2268 3921 2271
rect 3974 2268 3985 2271
rect 4238 2268 4246 2271
rect 4342 2268 4350 2271
rect 4574 2268 4582 2271
rect 2166 2258 2185 2261
rect 2270 2258 2289 2261
rect 2358 2258 2377 2261
rect 2550 2258 2574 2261
rect 2694 2258 2713 2261
rect 2726 2258 2745 2261
rect 2798 2258 2806 2261
rect 2826 2258 2841 2261
rect 2854 2258 2870 2261
rect 2890 2258 2905 2261
rect 2910 2258 2926 2261
rect 2934 2258 2950 2261
rect 3094 2258 3105 2261
rect 3526 2258 3534 2261
rect 3550 2261 3553 2268
rect 3974 2262 3977 2268
rect 3542 2258 3553 2261
rect 3622 2258 3641 2261
rect 3886 2258 3894 2261
rect 3914 2258 3921 2261
rect 3942 2258 3961 2261
rect 3990 2258 4001 2261
rect 4082 2258 4110 2261
rect 4266 2258 4273 2261
rect 4298 2258 4305 2261
rect 4350 2258 4361 2261
rect 4366 2258 4385 2261
rect 4442 2258 4449 2261
rect 4566 2258 4574 2261
rect 30 2257 34 2258
rect 678 2251 682 2254
rect 686 2251 689 2258
rect 678 2248 689 2251
rect 1062 2248 1070 2251
rect 2182 2248 2185 2258
rect 2242 2248 2249 2251
rect 2614 2251 2617 2258
rect 2614 2248 2625 2251
rect 2710 2248 2713 2258
rect 2786 2248 2793 2251
rect 2798 2248 2801 2258
rect 2854 2248 2857 2258
rect 2910 2248 2913 2258
rect 3102 2252 3105 2258
rect 3170 2248 3177 2251
rect 3246 2248 3254 2251
rect 3526 2248 3529 2258
rect 3558 2248 3566 2251
rect 3606 2251 3609 2258
rect 3598 2248 3609 2251
rect 3622 2248 3625 2258
rect 3710 2248 3721 2251
rect 3846 2248 3857 2251
rect 4254 2248 4262 2251
rect 4302 2248 4305 2258
rect 4350 2252 4353 2258
rect 4430 2248 4441 2251
rect 4506 2248 4513 2251
rect 2813 2238 2814 2242
rect 3358 2241 3361 2248
rect 3350 2238 3361 2241
rect 4518 2241 4521 2251
rect 4514 2238 4521 2241
rect 4565 2238 4566 2242
rect 1562 2218 1577 2221
rect 496 2203 498 2207
rect 502 2203 505 2207
rect 509 2203 512 2207
rect 1520 2203 1522 2207
rect 1526 2203 1529 2207
rect 1533 2203 1536 2207
rect 2544 2203 2546 2207
rect 2550 2203 2553 2207
rect 2557 2203 2560 2207
rect 3568 2203 3570 2207
rect 3574 2203 3577 2207
rect 3581 2203 3584 2207
rect 2757 2188 2758 2192
rect 3186 2188 3187 2192
rect 3234 2188 3235 2192
rect 3869 2188 3870 2192
rect 4301 2188 4302 2192
rect 4330 2188 4331 2192
rect 4477 2188 4478 2192
rect 4557 2188 4558 2192
rect 3518 2172 3521 2181
rect 4134 2172 4137 2181
rect 3350 2168 3361 2171
rect 4022 2168 4038 2171
rect 4253 2168 4254 2172
rect 4426 2168 4427 2172
rect 1158 2161 1161 2168
rect 1158 2158 1169 2161
rect 1438 2161 1441 2168
rect 1438 2158 1449 2161
rect 774 2153 778 2158
rect 526 2148 542 2151
rect 990 2148 998 2151
rect 1822 2148 1830 2151
rect 2206 2151 2209 2158
rect 2198 2148 2209 2151
rect 2214 2148 2222 2151
rect 2254 2151 2257 2161
rect 2238 2148 2257 2151
rect 2326 2151 2329 2158
rect 2374 2151 2377 2161
rect 2454 2161 2457 2168
rect 2446 2158 2457 2161
rect 3094 2158 3102 2161
rect 3470 2158 3481 2161
rect 3514 2158 3521 2161
rect 3702 2161 3705 2168
rect 3694 2158 3705 2161
rect 3794 2158 3798 2162
rect 2326 2148 2337 2151
rect 2358 2148 2377 2151
rect 2390 2148 2398 2151
rect 2710 2148 2729 2151
rect 2878 2148 2889 2151
rect 206 2138 218 2141
rect 542 2138 558 2141
rect 814 2138 830 2141
rect 918 2138 945 2141
rect 1466 2138 1473 2141
rect 1482 2138 1489 2141
rect 1594 2138 1601 2141
rect 2402 2138 2417 2141
rect 2654 2141 2657 2148
rect 2646 2138 2657 2141
rect 2830 2138 2857 2141
rect 2950 2141 2953 2151
rect 3010 2148 3017 2151
rect 3046 2148 3070 2151
rect 3354 2148 3361 2151
rect 3366 2148 3374 2151
rect 3390 2148 3409 2151
rect 3606 2148 3617 2151
rect 3722 2148 3729 2151
rect 3854 2148 3865 2151
rect 3910 2148 3918 2151
rect 4090 2148 4105 2151
rect 4190 2148 4198 2151
rect 4238 2151 4241 2161
rect 4534 2158 4545 2161
rect 4222 2148 4241 2151
rect 4290 2148 4297 2151
rect 4374 2148 4382 2151
rect 4558 2148 4577 2151
rect 2950 2138 2966 2141
rect 3066 2138 3073 2141
rect 3170 2138 3177 2141
rect 3318 2141 3321 2148
rect 3606 2142 3609 2148
rect 3294 2138 3321 2141
rect 3350 2138 3358 2141
rect 3646 2141 3649 2148
rect 3862 2142 3865 2148
rect 3646 2138 3657 2141
rect 3918 2138 3929 2141
rect 4054 2138 4066 2141
rect 4166 2138 4174 2141
rect 4366 2138 4390 2141
rect 4442 2138 4449 2141
rect 542 2128 545 2138
rect 670 2131 674 2133
rect 678 2131 681 2138
rect 1206 2132 1209 2138
rect 670 2128 681 2131
rect 950 2128 966 2131
rect 1138 2128 1150 2131
rect 1174 2128 1193 2131
rect 1206 2128 1214 2132
rect 1486 2128 1489 2138
rect 1806 2132 1810 2136
rect 1494 2128 1502 2131
rect 1998 2132 2002 2136
rect 3270 2132 3273 2138
rect 2942 2128 2950 2131
rect 3124 2128 3126 2132
rect 3142 2128 3161 2131
rect 3266 2128 3273 2132
rect 3578 2128 3590 2131
rect 3902 2131 3905 2138
rect 3882 2128 3889 2131
rect 3894 2128 3905 2131
rect 3918 2132 3921 2138
rect 4054 2132 4057 2138
rect 3950 2128 3961 2131
rect 4434 2128 4441 2131
rect 4522 2128 4529 2131
rect 4582 2128 4590 2131
rect 2482 2118 2484 2122
rect 1000 2103 1002 2107
rect 1006 2103 1009 2107
rect 1013 2103 1016 2107
rect 2024 2103 2026 2107
rect 2030 2103 2033 2107
rect 2037 2103 2040 2107
rect 3048 2103 3050 2107
rect 3054 2103 3057 2107
rect 3061 2103 3064 2107
rect 4080 2103 4082 2107
rect 4086 2103 4089 2107
rect 4093 2103 4096 2107
rect 2438 2088 2446 2091
rect 2964 2088 2966 2092
rect 3122 2088 3123 2092
rect 3293 2088 3294 2092
rect 3549 2088 3550 2092
rect 998 2078 1006 2081
rect 1214 2078 1233 2081
rect 1606 2078 1617 2081
rect 1966 2078 1982 2081
rect 346 2068 348 2072
rect 418 2068 425 2071
rect 670 2068 678 2071
rect 814 2071 817 2078
rect 804 2068 817 2071
rect 958 2068 977 2071
rect 1078 2071 1081 2078
rect 1966 2074 1970 2078
rect 1050 2068 1065 2071
rect 1070 2068 1081 2071
rect 46 2058 58 2061
rect 374 2058 393 2061
rect 406 2058 422 2061
rect 426 2058 433 2061
rect 1074 2058 1089 2061
rect 1126 2061 1129 2068
rect 1174 2062 1177 2071
rect 1366 2068 1377 2071
rect 1526 2068 1561 2071
rect 1666 2068 1678 2071
rect 2398 2071 2401 2081
rect 3654 2078 3665 2081
rect 3670 2078 3681 2081
rect 3722 2078 3729 2081
rect 4210 2078 4217 2081
rect 3678 2072 3681 2078
rect 2350 2068 2361 2071
rect 2382 2068 2401 2071
rect 2638 2068 2665 2071
rect 2710 2068 2721 2071
rect 2830 2068 2849 2071
rect 2878 2068 2889 2071
rect 2898 2068 2905 2071
rect 3014 2068 3033 2071
rect 3106 2068 3113 2071
rect 3364 2068 3377 2071
rect 3422 2068 3433 2071
rect 3470 2068 3481 2071
rect 3558 2068 3574 2071
rect 3630 2068 3638 2071
rect 3686 2068 3694 2071
rect 1118 2058 1129 2061
rect 1190 2058 1209 2061
rect 1242 2058 1254 2061
rect 1326 2061 1329 2068
rect 1366 2062 1369 2068
rect 1326 2058 1337 2061
rect 1526 2058 1529 2068
rect 1638 2061 1641 2068
rect 1578 2058 1585 2061
rect 1638 2058 1657 2061
rect 1702 2058 1713 2061
rect 2710 2062 2713 2068
rect 2878 2062 2881 2068
rect 3374 2062 3377 2068
rect 2226 2058 2233 2061
rect 2238 2058 2257 2061
rect 2270 2058 2289 2061
rect 2342 2058 2350 2061
rect 2358 2058 2377 2061
rect 2470 2058 2486 2061
rect 2542 2058 2569 2061
rect 2622 2058 2633 2061
rect 2818 2058 2825 2061
rect 2982 2058 3001 2061
rect 3070 2058 3089 2061
rect 3094 2058 3102 2061
rect 3142 2058 3161 2061
rect 3174 2058 3182 2061
rect 3218 2058 3225 2061
rect 3562 2058 3593 2061
rect 3654 2061 3657 2068
rect 3634 2058 3641 2061
rect 3646 2058 3657 2061
rect 3698 2058 3705 2061
rect 3710 2058 3718 2061
rect 3734 2058 3745 2061
rect 3818 2058 3825 2061
rect 3902 2061 3905 2071
rect 3938 2068 3945 2071
rect 4054 2068 4065 2071
rect 4134 2068 4142 2071
rect 4246 2071 4249 2081
rect 4486 2078 4497 2081
rect 4238 2068 4249 2071
rect 4322 2068 4329 2071
rect 4374 2068 4393 2071
rect 3902 2058 3913 2061
rect 3982 2058 3993 2061
rect 4166 2061 4169 2068
rect 4390 2062 4393 2068
rect 4158 2058 4169 2061
rect 4310 2058 4321 2061
rect 4494 2061 4497 2068
rect 4494 2058 4505 2061
rect 54 2057 58 2058
rect 326 2056 330 2058
rect 390 2048 393 2058
rect 494 2051 497 2058
rect 478 2048 497 2051
rect 526 2042 529 2051
rect 854 2048 865 2051
rect 982 2051 985 2058
rect 982 2048 993 2051
rect 1166 2048 1177 2051
rect 1342 2051 1345 2058
rect 1710 2052 1713 2058
rect 1342 2048 1353 2051
rect 2162 2048 2169 2051
rect 2204 2048 2206 2052
rect 2254 2048 2257 2058
rect 2630 2052 2633 2058
rect 2454 2048 2462 2051
rect 2858 2048 2862 2052
rect 2918 2051 2921 2058
rect 2918 2048 2929 2051
rect 3126 2048 3145 2051
rect 3174 2048 3177 2058
rect 3338 2048 3345 2051
rect 4350 2048 4358 2051
rect 755 2038 758 2042
rect 786 2038 793 2041
rect 1306 2038 1307 2042
rect 1827 2038 1830 2042
rect 2938 2038 2961 2041
rect 3346 2038 3361 2041
rect 2269 2028 2270 2032
rect 1138 2018 1139 2022
rect 2058 2018 2065 2021
rect 3794 2018 3795 2022
rect 4082 2018 4097 2021
rect 4565 2018 4566 2022
rect 496 2003 498 2007
rect 502 2003 505 2007
rect 509 2003 512 2007
rect 1520 2003 1522 2007
rect 1526 2003 1529 2007
rect 1533 2003 1536 2007
rect 2544 2003 2546 2007
rect 2550 2003 2553 2007
rect 2557 2003 2560 2007
rect 3568 2003 3570 2007
rect 3574 2003 3577 2007
rect 3581 2003 3584 2007
rect 2050 1988 2051 1992
rect 2530 1988 2531 1992
rect 2802 1988 2803 1992
rect 3786 1988 3787 1992
rect 4078 1988 4094 1991
rect 4330 1988 4331 1992
rect 397 1968 398 1972
rect 629 1968 630 1972
rect 1990 1968 1998 1971
rect 2085 1968 2086 1972
rect 3970 1968 3971 1972
rect 4294 1968 4305 1971
rect 4397 1968 4398 1972
rect 4498 1968 4499 1972
rect 270 1951 273 1961
rect 1614 1961 1617 1968
rect 4294 1962 4297 1968
rect 302 1952 306 1954
rect 270 1948 289 1951
rect 446 1948 454 1951
rect 510 1948 529 1951
rect 574 1948 582 1951
rect 510 1942 513 1948
rect 762 1948 769 1951
rect 1174 1951 1177 1958
rect 1166 1948 1177 1951
rect 1522 1948 1545 1951
rect 1558 1951 1561 1961
rect 1606 1958 1617 1961
rect 2126 1958 2145 1961
rect 2814 1958 2825 1961
rect 1554 1948 1561 1951
rect 1650 1948 1657 1951
rect 1662 1948 1689 1951
rect 1702 1948 1713 1951
rect 1806 1948 1814 1951
rect 2222 1948 2230 1951
rect 2290 1948 2297 1951
rect 2402 1948 2409 1951
rect 2574 1948 2585 1951
rect 2682 1948 2689 1951
rect 2734 1948 2742 1951
rect 2910 1948 2929 1951
rect 2950 1948 2961 1951
rect 3214 1948 3222 1951
rect 3310 1951 3313 1961
rect 3294 1948 3313 1951
rect 3330 1948 3345 1951
rect 3542 1948 3585 1951
rect 3606 1951 3609 1961
rect 3906 1958 3913 1961
rect 4342 1958 4353 1961
rect 3606 1948 3625 1951
rect 3790 1948 3806 1951
rect 3922 1948 3929 1951
rect 4006 1948 4033 1951
rect 4226 1948 4233 1951
rect 4278 1948 4289 1951
rect 4382 1951 4385 1961
rect 4378 1948 4385 1951
rect 4438 1951 4441 1961
rect 4510 1958 4521 1961
rect 4422 1948 4441 1951
rect 4542 1948 4550 1951
rect 350 1938 358 1941
rect 1118 1938 1142 1941
rect 1234 1938 1241 1941
rect 1262 1938 1281 1941
rect 1462 1941 1465 1948
rect 1454 1938 1465 1941
rect 1502 1938 1510 1941
rect 1578 1938 1593 1941
rect 1702 1938 1705 1948
rect 1946 1938 1953 1941
rect 2014 1938 2041 1941
rect 2094 1938 2105 1941
rect 2166 1938 2177 1941
rect 2334 1938 2353 1941
rect 2366 1938 2393 1941
rect 2430 1938 2441 1941
rect 2486 1938 2494 1941
rect 2590 1938 2609 1941
rect 3542 1942 3545 1948
rect 3582 1942 3585 1948
rect 2782 1938 2793 1941
rect 2870 1938 2886 1941
rect 2966 1938 2993 1941
rect 3046 1938 3089 1941
rect 3102 1938 3121 1941
rect 3142 1938 3150 1941
rect 3270 1938 3278 1941
rect 3282 1938 3286 1941
rect 3390 1938 3409 1941
rect 3474 1938 3481 1941
rect 3522 1938 3529 1941
rect 3630 1938 3641 1941
rect 3822 1938 3825 1948
rect 3846 1938 3849 1948
rect 4090 1938 4113 1941
rect 4134 1938 4150 1941
rect 4170 1938 4177 1941
rect 4270 1938 4278 1941
rect 4310 1938 4321 1941
rect 4454 1938 4473 1941
rect 4546 1938 4553 1941
rect 1278 1932 1281 1938
rect 2278 1932 2282 1933
rect 2430 1932 2433 1938
rect 1866 1928 1870 1932
rect 2474 1928 2481 1931
rect 2486 1928 2489 1938
rect 2750 1928 2761 1931
rect 2830 1928 2846 1931
rect 3006 1928 3025 1931
rect 3142 1928 3145 1938
rect 3406 1932 3409 1938
rect 3638 1932 3641 1938
rect 4310 1932 4313 1938
rect 4218 1928 4225 1931
rect 602 1918 603 1922
rect 654 1918 662 1921
rect 4162 1918 4163 1922
rect 4573 1918 4574 1922
rect 1000 1903 1002 1907
rect 1006 1903 1009 1907
rect 1013 1903 1016 1907
rect 2024 1903 2026 1907
rect 2030 1903 2033 1907
rect 2037 1903 2040 1907
rect 3048 1903 3050 1907
rect 3054 1903 3057 1907
rect 3061 1903 3064 1907
rect 4080 1903 4082 1907
rect 4086 1903 4089 1907
rect 4093 1903 4096 1907
rect 532 1888 534 1892
rect 1518 1888 1534 1891
rect 1933 1888 1934 1892
rect 2197 1888 2198 1892
rect 2986 1888 2987 1892
rect 4410 1888 4411 1892
rect 490 1868 505 1871
rect 646 1868 665 1871
rect 1150 1871 1153 1881
rect 1166 1878 1177 1881
rect 1310 1878 1321 1881
rect 1310 1872 1313 1878
rect 1150 1868 1169 1871
rect 1386 1868 1393 1871
rect 46 1858 58 1861
rect 646 1862 649 1868
rect 366 1858 382 1861
rect 538 1858 566 1861
rect 574 1858 593 1861
rect 962 1858 969 1861
rect 1126 1858 1137 1861
rect 1222 1858 1241 1861
rect 1302 1858 1313 1861
rect 1398 1858 1406 1861
rect 1642 1858 1660 1861
rect 54 1857 58 1858
rect 590 1848 593 1858
rect 1414 1848 1422 1851
rect 1734 1842 1737 1881
rect 1958 1878 1977 1881
rect 2106 1878 2113 1881
rect 2598 1878 2606 1881
rect 2742 1878 2758 1881
rect 2922 1878 2929 1881
rect 2742 1872 2745 1878
rect 1862 1868 1878 1871
rect 1978 1868 1985 1871
rect 2118 1868 2142 1871
rect 1874 1858 1897 1861
rect 2026 1858 2049 1861
rect 2082 1858 2089 1861
rect 2294 1861 2297 1871
rect 2326 1868 2345 1871
rect 2522 1868 2529 1871
rect 2294 1858 2305 1861
rect 2366 1858 2385 1861
rect 2518 1858 2521 1868
rect 2574 1858 2585 1861
rect 2638 1858 2649 1861
rect 2806 1861 2809 1871
rect 3006 1868 3014 1871
rect 3230 1868 3265 1871
rect 3286 1868 3294 1871
rect 3362 1868 3369 1871
rect 3478 1868 3486 1871
rect 3542 1868 3550 1871
rect 3686 1868 3697 1871
rect 3718 1871 3721 1878
rect 3838 1872 3841 1881
rect 3990 1878 4009 1881
rect 4062 1878 4073 1881
rect 4198 1872 4201 1881
rect 3718 1868 3729 1871
rect 4018 1868 4033 1871
rect 4038 1868 4046 1871
rect 4418 1868 4430 1871
rect 4454 1871 4457 1881
rect 4450 1868 4457 1871
rect 4502 1871 4505 1878
rect 4494 1868 4505 1871
rect 2790 1858 2809 1861
rect 2902 1861 2905 1868
rect 2826 1858 2841 1861
rect 2894 1858 2905 1861
rect 2934 1861 2937 1868
rect 2926 1858 2937 1861
rect 3222 1858 3230 1861
rect 3382 1858 3390 1861
rect 3418 1858 3433 1861
rect 3474 1858 3497 1861
rect 3646 1858 3665 1861
rect 3902 1858 3913 1861
rect 3958 1858 3966 1861
rect 4042 1858 4049 1861
rect 4190 1858 4206 1861
rect 4494 1858 4505 1861
rect 4546 1858 4561 1861
rect 1842 1849 1844 1853
rect 2294 1852 2297 1858
rect 2226 1848 2230 1852
rect 2542 1848 2550 1851
rect 2694 1848 2702 1851
rect 2842 1848 2846 1852
rect 2990 1848 3009 1851
rect 3030 1848 3041 1851
rect 3390 1848 3409 1851
rect 3446 1848 3454 1851
rect 3514 1848 3521 1851
rect 3662 1848 3665 1858
rect 3902 1852 3905 1858
rect 3786 1848 3793 1851
rect 3890 1848 3897 1851
rect 3958 1848 3961 1858
rect 4182 1848 4193 1851
rect 4326 1848 4337 1851
rect 4346 1848 4350 1852
rect 4562 1848 4566 1852
rect 437 1838 438 1842
rect 637 1838 638 1842
rect 1499 1838 1502 1842
rect 2286 1838 2294 1841
rect 2358 1841 2362 1844
rect 2350 1838 2362 1841
rect 2653 1838 2654 1842
rect 3469 1838 3470 1842
rect 4109 1838 4110 1842
rect 4390 1838 4398 1841
rect 1218 1828 1219 1832
rect 1274 1818 1275 1822
rect 2389 1818 2390 1822
rect 2469 1818 2470 1822
rect 2613 1818 2614 1822
rect 3189 1818 3190 1822
rect 3221 1818 3222 1822
rect 3306 1818 3307 1822
rect 3434 1818 3435 1822
rect 3498 1818 3499 1822
rect 3533 1818 3534 1822
rect 3677 1818 3678 1822
rect 3738 1818 3739 1822
rect 3770 1818 3771 1822
rect 3805 1818 3806 1822
rect 4053 1818 4054 1822
rect 4533 1818 4534 1822
rect 4594 1818 4595 1822
rect 496 1803 498 1807
rect 502 1803 505 1807
rect 509 1803 512 1807
rect 1520 1803 1522 1807
rect 1526 1803 1529 1807
rect 1533 1803 1536 1807
rect 2544 1803 2546 1807
rect 2550 1803 2553 1807
rect 2557 1803 2560 1807
rect 3568 1803 3570 1807
rect 3574 1803 3577 1807
rect 3581 1803 3584 1807
rect 204 1788 206 1792
rect 348 1788 350 1792
rect 1181 1788 1182 1792
rect 1550 1788 1566 1791
rect 1962 1788 1963 1792
rect 2810 1788 2811 1792
rect 702 1768 713 1771
rect 710 1761 713 1768
rect 1574 1768 1585 1771
rect 1898 1768 1905 1771
rect 2141 1768 2142 1772
rect 4394 1768 4395 1772
rect 4458 1768 4474 1771
rect 718 1761 721 1768
rect 1582 1762 1585 1768
rect 710 1758 721 1761
rect 278 1748 297 1751
rect 922 1748 929 1751
rect 250 1738 262 1741
rect 822 1738 830 1741
rect 982 1741 985 1751
rect 1018 1748 1041 1751
rect 1098 1748 1105 1751
rect 1134 1748 1153 1751
rect 1286 1751 1289 1761
rect 1910 1758 1926 1761
rect 1990 1758 2001 1761
rect 1270 1748 1289 1751
rect 982 1738 1001 1741
rect 1110 1741 1113 1748
rect 1862 1748 1873 1751
rect 1878 1748 1894 1751
rect 2054 1751 2057 1761
rect 1966 1748 1985 1751
rect 1998 1748 2017 1751
rect 2022 1748 2057 1751
rect 2062 1748 2078 1751
rect 2094 1748 2105 1751
rect 2166 1748 2177 1751
rect 2526 1748 2561 1751
rect 2826 1748 2833 1751
rect 3174 1751 3177 1761
rect 3310 1758 3318 1761
rect 3158 1748 3177 1751
rect 3210 1748 3217 1751
rect 3438 1751 3441 1761
rect 3478 1758 3497 1761
rect 3718 1758 3737 1761
rect 3742 1758 3750 1761
rect 3410 1748 3425 1751
rect 3438 1748 3457 1751
rect 3650 1748 3665 1751
rect 3866 1748 3873 1751
rect 3878 1748 3897 1751
rect 4170 1748 4177 1751
rect 4210 1748 4217 1751
rect 4406 1751 4409 1761
rect 4510 1758 4529 1761
rect 4406 1748 4425 1751
rect 4462 1751 4466 1754
rect 4462 1748 4481 1751
rect 2174 1742 2177 1748
rect 1110 1738 1121 1741
rect 1330 1738 1345 1741
rect 1678 1738 1686 1741
rect 1814 1738 1822 1741
rect 2202 1738 2209 1741
rect 2510 1738 2521 1741
rect 2566 1738 2590 1741
rect 2710 1738 2734 1741
rect 2794 1738 2809 1741
rect 2870 1738 2889 1741
rect 2946 1738 2953 1741
rect 3038 1738 3081 1741
rect 3086 1738 3105 1741
rect 3262 1738 3265 1748
rect 3302 1741 3305 1748
rect 3294 1738 3305 1741
rect 3350 1738 3361 1741
rect 3406 1738 3414 1741
rect 3462 1738 3470 1741
rect 3622 1738 3630 1741
rect 3638 1738 3657 1741
rect 3746 1738 3753 1741
rect 3878 1742 3881 1748
rect 3846 1738 3862 1741
rect 4122 1738 4129 1741
rect 4158 1738 4166 1741
rect 4378 1738 4385 1741
rect 4550 1738 4561 1741
rect 4570 1738 4585 1741
rect 1006 1728 1022 1731
rect 1062 1728 1073 1731
rect 1794 1728 1809 1731
rect 1814 1728 1817 1738
rect 2870 1732 2873 1738
rect 2242 1728 2249 1731
rect 2294 1728 2302 1731
rect 2790 1728 2798 1731
rect 4126 1728 4129 1738
rect 4134 1728 4153 1731
rect 242 1718 243 1722
rect 1354 1718 1355 1722
rect 1598 1718 1606 1721
rect 2453 1718 2454 1722
rect 3397 1718 3398 1722
rect 3821 1718 3822 1722
rect 4090 1718 4097 1721
rect 4330 1718 4331 1722
rect 1000 1703 1002 1707
rect 1006 1703 1009 1707
rect 1013 1703 1016 1707
rect 2024 1703 2026 1707
rect 2030 1703 2033 1707
rect 2037 1703 2040 1707
rect 3048 1703 3050 1707
rect 3054 1703 3057 1707
rect 3061 1703 3064 1707
rect 4080 1703 4082 1707
rect 4086 1703 4089 1707
rect 4093 1703 4096 1707
rect 2030 1688 2038 1691
rect 3005 1688 3006 1692
rect 162 1678 177 1681
rect 286 1678 297 1681
rect 1182 1678 1193 1681
rect 2142 1678 2150 1681
rect 286 1672 289 1678
rect 2182 1672 2185 1681
rect 2246 1678 2254 1682
rect 2422 1678 2430 1681
rect 2546 1678 2577 1681
rect 3038 1678 3057 1681
rect 3062 1678 3070 1681
rect 3258 1678 3265 1681
rect 4342 1678 4353 1681
rect 2246 1672 2249 1678
rect 334 1668 342 1671
rect 410 1668 417 1671
rect 526 1668 534 1671
rect 1686 1668 1694 1671
rect 1958 1668 1969 1671
rect 2102 1668 2113 1671
rect 470 1658 478 1661
rect 546 1658 553 1661
rect 1258 1658 1270 1661
rect 1542 1658 1550 1661
rect 1586 1658 1610 1661
rect 1690 1658 1697 1661
rect 1846 1661 1849 1668
rect 1822 1658 1841 1661
rect 1846 1658 1865 1661
rect 1998 1658 2017 1661
rect 2106 1658 2113 1661
rect 2190 1661 2193 1671
rect 2198 1668 2217 1671
rect 2406 1668 2417 1671
rect 2470 1668 2489 1671
rect 2606 1668 2625 1671
rect 2622 1662 2625 1668
rect 2642 1668 2649 1671
rect 2954 1668 2961 1671
rect 3478 1671 3481 1678
rect 3470 1668 3481 1671
rect 3486 1668 3497 1671
rect 3750 1668 3761 1671
rect 3806 1668 3814 1671
rect 4250 1668 4262 1671
rect 4322 1668 4329 1671
rect 4414 1671 4417 1678
rect 4446 1671 4449 1681
rect 4550 1678 4569 1681
rect 4374 1668 4385 1671
rect 4406 1668 4417 1671
rect 4422 1668 4449 1671
rect 2146 1658 2153 1661
rect 2174 1658 2193 1661
rect 2526 1658 2537 1661
rect 2594 1658 2601 1661
rect 2638 1658 2641 1668
rect 2942 1658 2953 1661
rect 3114 1658 3129 1661
rect 3206 1658 3226 1661
rect 3246 1658 3257 1661
rect 3274 1658 3289 1661
rect 3346 1658 3353 1661
rect 3382 1658 3390 1661
rect 3422 1658 3430 1661
rect 3486 1661 3489 1668
rect 4374 1662 4377 1668
rect 4526 1662 4529 1671
rect 3478 1658 3489 1661
rect 3566 1658 3574 1661
rect 3594 1658 3601 1661
rect 3638 1658 3646 1661
rect 3886 1658 3894 1661
rect 3906 1658 3913 1661
rect 3982 1658 4001 1661
rect 4018 1658 4033 1661
rect 4070 1658 4113 1661
rect 4150 1658 4170 1661
rect 4222 1658 4233 1661
rect 4386 1658 4393 1661
rect 4490 1658 4513 1661
rect 862 1656 866 1658
rect 1606 1656 1610 1658
rect 230 1648 241 1651
rect 178 1638 185 1641
rect 242 1638 257 1641
rect 325 1638 326 1642
rect 458 1638 461 1642
rect 678 1641 681 1651
rect 710 1648 718 1651
rect 1230 1648 1241 1651
rect 1510 1651 1514 1654
rect 1998 1652 2001 1658
rect 2534 1652 2537 1658
rect 3222 1656 3226 1658
rect 1510 1648 1518 1651
rect 1918 1648 1937 1651
rect 2030 1648 2065 1651
rect 2090 1648 2094 1652
rect 2366 1648 2385 1651
rect 2722 1648 2729 1651
rect 3098 1648 3102 1652
rect 3670 1651 3673 1658
rect 3662 1648 3673 1651
rect 3834 1648 3838 1652
rect 3946 1648 3950 1652
rect 3998 1648 4001 1658
rect 4030 1648 4033 1658
rect 4166 1656 4170 1658
rect 4278 1648 4289 1651
rect 670 1638 681 1641
rect 1658 1638 1660 1642
rect 1786 1638 1801 1641
rect 1986 1638 1993 1641
rect 2254 1638 2262 1641
rect 2426 1638 2433 1641
rect 2710 1638 2718 1641
rect 3858 1638 3865 1641
rect 1866 1618 1867 1622
rect 1949 1618 1950 1622
rect 2397 1618 2398 1622
rect 2586 1618 2587 1622
rect 2658 1618 2659 1622
rect 3154 1618 3155 1622
rect 3301 1618 3302 1622
rect 3370 1618 3371 1622
rect 3554 1618 3555 1622
rect 3741 1618 3742 1622
rect 4013 1618 4014 1622
rect 4125 1618 4126 1622
rect 4237 1618 4238 1622
rect 496 1603 498 1607
rect 502 1603 505 1607
rect 509 1603 512 1607
rect 1520 1603 1522 1607
rect 1526 1603 1529 1607
rect 1533 1603 1536 1607
rect 2544 1603 2546 1607
rect 2550 1603 2553 1607
rect 2557 1603 2560 1607
rect 3568 1603 3570 1607
rect 3574 1603 3577 1607
rect 3581 1603 3584 1607
rect 253 1588 254 1592
rect 557 1588 558 1592
rect 2818 1588 2819 1592
rect 3045 1588 3046 1592
rect 3093 1588 3094 1592
rect 522 1578 529 1581
rect 589 1578 590 1582
rect 618 1578 619 1582
rect 3445 1578 3446 1582
rect 4070 1581 4073 1588
rect 4062 1578 4073 1581
rect 963 1568 966 1572
rect 1822 1568 1849 1571
rect 1957 1568 1958 1572
rect 2526 1568 2537 1571
rect 3846 1568 3858 1571
rect 4242 1568 4243 1572
rect 230 1566 234 1568
rect 630 1552 633 1561
rect 758 1558 766 1561
rect 1158 1558 1169 1561
rect 1438 1558 1449 1561
rect 1578 1558 1580 1562
rect 2278 1561 2281 1568
rect 2526 1562 2529 1568
rect 3854 1566 3858 1568
rect 4374 1566 4378 1568
rect 1158 1552 1161 1558
rect 142 1548 150 1551
rect 190 1548 225 1551
rect 274 1548 281 1551
rect 286 1548 294 1551
rect 406 1548 433 1551
rect 594 1548 617 1551
rect 190 1538 193 1548
rect 1118 1548 1129 1551
rect 1310 1548 1342 1551
rect 1358 1548 1366 1551
rect 1406 1548 1425 1551
rect 1550 1548 1558 1551
rect 1642 1548 1649 1551
rect 1118 1542 1121 1548
rect 210 1538 217 1541
rect 390 1538 401 1541
rect 478 1538 497 1541
rect 602 1538 609 1541
rect 1058 1538 1065 1541
rect 1094 1538 1105 1541
rect 1190 1538 1198 1541
rect 1554 1538 1561 1541
rect 1782 1538 1790 1541
rect 1998 1541 2001 1551
rect 2026 1548 2057 1551
rect 2062 1548 2078 1551
rect 2142 1551 2145 1561
rect 2126 1548 2145 1551
rect 2206 1551 2209 1561
rect 2278 1558 2289 1561
rect 2202 1548 2209 1551
rect 2226 1548 2233 1551
rect 2270 1548 2278 1551
rect 2394 1548 2401 1551
rect 2510 1551 2513 1561
rect 2498 1548 2513 1551
rect 2534 1548 2569 1551
rect 2718 1548 2726 1551
rect 2918 1551 2921 1561
rect 3178 1558 3182 1562
rect 2142 1542 2145 1548
rect 1998 1538 2017 1541
rect 2094 1538 2102 1541
rect 2114 1538 2121 1541
rect 2158 1538 2166 1541
rect 2170 1538 2177 1541
rect 2294 1541 2297 1548
rect 2254 1538 2273 1541
rect 2294 1538 2305 1541
rect 2322 1538 2329 1541
rect 2414 1538 2425 1541
rect 2566 1538 2569 1548
rect 2654 1538 2665 1541
rect 2698 1538 2705 1541
rect 2746 1538 2761 1541
rect 2894 1541 2897 1551
rect 2902 1548 2921 1551
rect 3198 1551 3201 1561
rect 3206 1558 3225 1561
rect 3426 1558 3433 1561
rect 3170 1548 3177 1551
rect 3182 1548 3201 1551
rect 3226 1548 3233 1551
rect 3450 1548 3465 1551
rect 3598 1551 3601 1561
rect 3566 1548 3601 1551
rect 3654 1548 3662 1551
rect 3782 1548 3790 1551
rect 3822 1551 3825 1561
rect 4358 1558 4377 1561
rect 4474 1558 4478 1562
rect 4486 1558 4505 1561
rect 3822 1548 3841 1551
rect 3846 1548 3854 1551
rect 3894 1551 3897 1558
rect 3894 1548 3905 1551
rect 4034 1548 4041 1551
rect 4082 1548 4089 1551
rect 4446 1548 4462 1551
rect 2794 1538 2809 1541
rect 2878 1538 2897 1541
rect 2914 1538 2929 1541
rect 2934 1538 2945 1541
rect 2966 1538 2985 1541
rect 3338 1538 3345 1541
rect 3462 1541 3465 1548
rect 3462 1538 3473 1541
rect 3654 1538 3657 1548
rect 3666 1538 3681 1541
rect 3714 1538 3726 1541
rect 3966 1538 3974 1541
rect 3998 1541 4001 1548
rect 3990 1538 4001 1541
rect 4030 1538 4038 1541
rect 4118 1538 4134 1541
rect 4290 1538 4297 1541
rect 4318 1538 4337 1541
rect 4422 1538 4433 1541
rect 4514 1538 4521 1541
rect 398 1532 401 1538
rect 186 1528 193 1531
rect 1190 1528 1193 1538
rect 1202 1528 1206 1532
rect 1382 1528 1398 1531
rect 1454 1528 1462 1531
rect 1542 1528 1550 1531
rect 1726 1528 1737 1531
rect 2010 1528 2017 1531
rect 2022 1528 2030 1531
rect 2094 1528 2097 1538
rect 2254 1528 2257 1538
rect 226 1518 227 1522
rect 1114 1518 1115 1522
rect 1501 1518 1502 1522
rect 1773 1518 1774 1522
rect 2149 1518 2150 1522
rect 2178 1518 2179 1522
rect 2341 1518 2342 1522
rect 2734 1518 2742 1521
rect 3861 1518 3862 1522
rect 4381 1518 4382 1522
rect 1000 1503 1002 1507
rect 1006 1503 1009 1507
rect 1013 1503 1016 1507
rect 2024 1503 2026 1507
rect 2030 1503 2033 1507
rect 2037 1503 2040 1507
rect 3048 1503 3050 1507
rect 3054 1503 3057 1507
rect 3061 1503 3064 1507
rect 4080 1503 4082 1507
rect 4086 1503 4089 1507
rect 4093 1503 4096 1507
rect 277 1488 278 1492
rect 442 1488 443 1492
rect 1124 1488 1126 1492
rect 1890 1488 1892 1492
rect 2030 1488 2046 1491
rect 2702 1488 2710 1491
rect 2885 1488 2886 1492
rect 2970 1488 2971 1492
rect 3501 1488 3502 1492
rect 3842 1488 3855 1491
rect 4130 1488 4131 1492
rect 4196 1488 4198 1492
rect 174 1478 182 1481
rect 198 1471 201 1481
rect 226 1478 233 1481
rect 998 1478 1006 1482
rect 1270 1478 1278 1482
rect 1538 1478 1542 1482
rect 1670 1478 1689 1481
rect 2654 1481 2657 1488
rect 2646 1478 2657 1481
rect 2686 1478 2700 1481
rect 998 1472 1001 1478
rect 1270 1472 1273 1478
rect 2750 1472 2753 1481
rect 2942 1478 2950 1481
rect 3098 1478 3105 1481
rect 3878 1478 3886 1481
rect 166 1468 193 1471
rect 198 1468 217 1471
rect 238 1468 249 1471
rect 402 1468 409 1471
rect 622 1468 634 1471
rect 210 1458 217 1461
rect 222 1458 230 1461
rect 290 1458 297 1461
rect 366 1458 377 1461
rect 622 1462 625 1468
rect 862 1461 865 1471
rect 1486 1468 1497 1471
rect 1522 1468 1537 1471
rect 1614 1468 1622 1471
rect 1750 1468 1761 1471
rect 1798 1468 1809 1471
rect 1486 1462 1489 1468
rect 1918 1462 1921 1471
rect 1998 1468 2006 1471
rect 2162 1468 2169 1471
rect 2310 1468 2321 1471
rect 2318 1462 2321 1468
rect 862 1458 878 1461
rect 1142 1458 1153 1461
rect 1202 1458 1209 1461
rect 1298 1458 1305 1461
rect 1622 1458 1630 1461
rect 1690 1458 1702 1461
rect 1830 1458 1849 1461
rect 1958 1458 1966 1461
rect 1990 1458 2014 1461
rect 2058 1458 2065 1461
rect 2118 1458 2137 1461
rect 2502 1461 2505 1471
rect 2590 1468 2598 1471
rect 2902 1468 2913 1471
rect 2954 1468 2961 1471
rect 3038 1468 3054 1471
rect 2902 1462 2905 1468
rect 3198 1462 3201 1471
rect 3758 1468 3777 1471
rect 4054 1471 4057 1481
rect 4054 1468 4065 1471
rect 4138 1468 4145 1471
rect 4318 1471 4321 1481
rect 4318 1468 4326 1471
rect 4462 1471 4465 1478
rect 4454 1468 4465 1471
rect 4582 1468 4590 1471
rect 2494 1458 2505 1461
rect 2526 1458 2545 1461
rect 2950 1458 2958 1461
rect 3006 1458 3025 1461
rect 3122 1458 3129 1461
rect 3222 1458 3230 1461
rect 3422 1458 3438 1461
rect 3446 1458 3454 1461
rect 3478 1458 3497 1461
rect 3542 1461 3545 1468
rect 3774 1462 3777 1468
rect 4062 1462 4065 1468
rect 3542 1458 3553 1461
rect 3586 1458 3601 1461
rect 3682 1458 3689 1461
rect 4046 1458 4054 1461
rect 4222 1458 4230 1461
rect 4350 1458 4369 1461
rect 366 1452 369 1458
rect 1150 1452 1153 1458
rect 290 1438 297 1441
rect 726 1441 729 1451
rect 978 1448 982 1452
rect 1186 1448 1190 1452
rect 1230 1448 1241 1451
rect 1446 1448 1457 1451
rect 1830 1448 1833 1458
rect 2134 1448 2137 1458
rect 2146 1448 2150 1452
rect 2238 1448 2249 1451
rect 2338 1448 2342 1452
rect 2526 1448 2529 1458
rect 3006 1448 3009 1458
rect 3218 1448 3222 1452
rect 3422 1448 3425 1458
rect 3494 1448 3497 1458
rect 4350 1448 4353 1458
rect 4506 1448 4513 1451
rect 3494 1442 3498 1444
rect 718 1438 729 1441
rect 1050 1438 1057 1441
rect 1574 1438 1582 1441
rect 1866 1438 1873 1441
rect 2226 1438 2227 1442
rect 2677 1438 2678 1442
rect 2746 1438 2753 1441
rect 2994 1438 2995 1442
rect 3966 1438 3982 1441
rect 4221 1438 4222 1442
rect 1645 1428 1646 1432
rect 466 1418 473 1421
rect 909 1418 910 1422
rect 1402 1418 1404 1422
rect 1770 1418 1771 1422
rect 1818 1418 1819 1422
rect 1989 1418 1990 1422
rect 2445 1418 2446 1422
rect 2514 1418 2515 1422
rect 2797 1418 2798 1422
rect 3130 1418 3131 1422
rect 3410 1418 3411 1422
rect 3533 1418 3534 1422
rect 3557 1418 3558 1422
rect 3810 1418 3811 1422
rect 3941 1418 3942 1422
rect 496 1403 498 1407
rect 502 1403 505 1407
rect 509 1403 512 1407
rect 1520 1403 1522 1407
rect 1526 1403 1529 1407
rect 1533 1403 1536 1407
rect 2544 1403 2546 1407
rect 2550 1403 2553 1407
rect 2557 1403 2560 1407
rect 3568 1403 3570 1407
rect 3574 1403 3577 1407
rect 3581 1403 3584 1407
rect 562 1388 563 1392
rect 1330 1388 1331 1392
rect 1898 1388 1899 1392
rect 1978 1388 1979 1392
rect 2805 1388 2806 1392
rect 3509 1388 3510 1392
rect 3725 1388 3726 1392
rect 4078 1388 4086 1391
rect 4234 1388 4235 1392
rect 4333 1388 4334 1392
rect 4530 1388 4531 1392
rect 597 1378 598 1382
rect 1166 1368 1174 1371
rect 1918 1368 1929 1371
rect 2610 1368 2611 1372
rect 1918 1362 1921 1368
rect 330 1348 337 1351
rect 342 1348 369 1351
rect 382 1351 385 1361
rect 1254 1358 1265 1361
rect 1694 1358 1713 1361
rect 1254 1352 1257 1358
rect 382 1348 401 1351
rect 482 1348 497 1351
rect 546 1348 561 1351
rect 1130 1348 1145 1351
rect 1186 1348 1193 1351
rect 1334 1348 1353 1351
rect 1434 1348 1457 1351
rect 1468 1348 1494 1351
rect 1910 1351 1913 1361
rect 1910 1348 1918 1351
rect 2134 1348 2142 1351
rect 2230 1351 2233 1361
rect 2434 1358 2438 1362
rect 3570 1358 3585 1361
rect 2230 1348 2238 1351
rect 406 1338 414 1341
rect 746 1338 753 1341
rect 910 1338 921 1341
rect 1206 1338 1225 1341
rect 1926 1338 1945 1341
rect 2014 1341 2017 1348
rect 2014 1338 2041 1341
rect 2078 1338 2089 1341
rect 2270 1341 2273 1351
rect 2398 1348 2406 1351
rect 2806 1348 2833 1351
rect 3262 1348 3273 1351
rect 3378 1348 3385 1351
rect 3390 1348 3409 1351
rect 3598 1348 3614 1351
rect 3798 1348 3809 1351
rect 4206 1348 4214 1351
rect 4542 1348 4566 1351
rect 3262 1342 3265 1348
rect 3390 1342 3393 1348
rect 2270 1338 2305 1341
rect 2374 1338 2393 1341
rect 2460 1338 2473 1341
rect 2870 1338 2886 1341
rect 2978 1338 2985 1341
rect 3302 1338 3329 1341
rect 3562 1338 3585 1341
rect 3810 1338 3817 1341
rect 3966 1341 3969 1348
rect 3958 1338 3969 1341
rect 4110 1338 4129 1341
rect 4454 1341 4457 1348
rect 4414 1338 4425 1341
rect 4454 1338 4465 1341
rect 1114 1328 1121 1331
rect 1174 1328 1185 1331
rect 1422 1328 1441 1331
rect 1566 1328 1577 1331
rect 1614 1328 1625 1331
rect 1778 1328 1785 1331
rect 2006 1328 2014 1331
rect 2302 1328 2305 1338
rect 2390 1332 2393 1338
rect 2470 1332 2473 1338
rect 3222 1328 3241 1331
rect 1301 1318 1302 1322
rect 1397 1318 1398 1322
rect 1805 1318 1806 1322
rect 2194 1318 2195 1322
rect 2834 1318 2835 1322
rect 3062 1318 3070 1321
rect 3162 1318 3163 1322
rect 3754 1318 3755 1322
rect 1000 1303 1002 1307
rect 1006 1303 1009 1307
rect 1013 1303 1016 1307
rect 2024 1303 2026 1307
rect 2030 1303 2033 1307
rect 2037 1303 2040 1307
rect 3048 1303 3050 1307
rect 3054 1303 3057 1307
rect 3061 1303 3064 1307
rect 4080 1303 4082 1307
rect 4086 1303 4089 1307
rect 4093 1303 4096 1307
rect 162 1288 163 1292
rect 1189 1288 1190 1292
rect 1260 1288 1262 1292
rect 2477 1288 2478 1292
rect 2525 1288 2526 1292
rect 3130 1288 3131 1292
rect 3194 1288 3215 1291
rect 3485 1288 3486 1292
rect 262 1268 286 1271
rect 358 1268 369 1271
rect 406 1268 417 1271
rect 462 1268 473 1271
rect 926 1268 937 1271
rect 998 1268 1022 1271
rect 1038 1271 1041 1281
rect 2038 1278 2065 1281
rect 2134 1278 2145 1281
rect 2220 1278 2222 1282
rect 2398 1278 2406 1281
rect 3390 1278 3398 1281
rect 1038 1268 1054 1271
rect 1082 1268 1089 1271
rect 1278 1268 1286 1271
rect 1350 1268 1358 1271
rect 1598 1268 1614 1271
rect 46 1258 58 1261
rect 214 1258 222 1261
rect 238 1258 254 1261
rect 326 1261 329 1268
rect 318 1258 329 1261
rect 366 1262 369 1268
rect 470 1262 473 1268
rect 374 1258 393 1261
rect 1214 1258 1230 1261
rect 1430 1258 1441 1261
rect 1470 1258 1486 1261
rect 1566 1258 1574 1261
rect 1670 1261 1673 1271
rect 1702 1268 1710 1271
rect 1766 1268 1774 1271
rect 1846 1268 1857 1271
rect 1950 1268 1969 1271
rect 1854 1262 1857 1268
rect 1670 1258 1681 1261
rect 1726 1258 1734 1261
rect 1770 1258 1785 1261
rect 1918 1261 1921 1268
rect 2162 1268 2177 1271
rect 1890 1258 1897 1261
rect 1910 1258 1921 1261
rect 1998 1258 2017 1261
rect 2190 1261 2193 1268
rect 2286 1271 2289 1278
rect 2278 1268 2289 1271
rect 2294 1268 2313 1271
rect 2362 1268 2369 1271
rect 2438 1268 2465 1271
rect 2534 1268 2542 1271
rect 2670 1268 2686 1271
rect 2734 1268 2750 1271
rect 2830 1268 2849 1271
rect 2974 1268 2990 1271
rect 3062 1268 3070 1271
rect 3174 1268 3185 1271
rect 3326 1268 3334 1271
rect 3450 1268 3457 1271
rect 3518 1271 3521 1281
rect 3518 1268 3526 1271
rect 3726 1268 3734 1271
rect 3750 1268 3758 1271
rect 3174 1262 3177 1268
rect 2182 1258 2193 1261
rect 2358 1258 2366 1261
rect 2398 1258 2409 1261
rect 2414 1258 2433 1261
rect 2502 1258 2521 1261
rect 2682 1258 2697 1261
rect 2810 1258 2817 1261
rect 2910 1258 2918 1261
rect 2942 1258 2950 1261
rect 3054 1258 3062 1261
rect 3302 1258 3321 1261
rect 3414 1258 3422 1261
rect 3530 1258 3537 1261
rect 3550 1258 3585 1261
rect 3830 1261 3833 1271
rect 3882 1268 3889 1271
rect 4062 1268 4073 1271
rect 4098 1268 4105 1271
rect 4062 1262 4065 1268
rect 3814 1258 3833 1261
rect 3846 1258 3865 1261
rect 3914 1258 3921 1261
rect 3978 1258 3985 1261
rect 4134 1261 4137 1271
rect 4286 1268 4305 1271
rect 4330 1268 4342 1271
rect 4438 1268 4449 1271
rect 4534 1268 4542 1271
rect 4126 1258 4137 1261
rect 4282 1258 4289 1261
rect 4302 1258 4305 1268
rect 4438 1262 4441 1268
rect 4526 1258 4534 1261
rect 54 1257 58 1258
rect 1302 1256 1306 1258
rect 1438 1252 1441 1258
rect 554 1248 561 1251
rect 1294 1248 1305 1251
rect 1494 1248 1505 1251
rect 1546 1248 1553 1251
rect 1798 1248 1806 1251
rect 1910 1248 1913 1258
rect 1934 1248 1953 1251
rect 2090 1248 2094 1252
rect 2370 1248 2377 1251
rect 2518 1248 2521 1258
rect 2938 1248 2942 1252
rect 3550 1248 3553 1258
rect 3846 1248 3849 1258
rect 4350 1248 4369 1251
rect 534 1238 542 1241
rect 1156 1238 1158 1242
rect 1446 1238 1454 1241
rect 1590 1238 1598 1241
rect 1898 1238 1899 1242
rect 2998 1238 3006 1241
rect 4493 1238 4494 1242
rect 522 1228 529 1231
rect 3621 1228 3622 1232
rect 1010 1218 1025 1221
rect 1378 1218 1379 1222
rect 1565 1218 1566 1222
rect 1757 1218 1758 1222
rect 1786 1218 1787 1222
rect 2322 1218 2323 1222
rect 3053 1218 3054 1222
rect 3381 1218 3382 1222
rect 3682 1218 3683 1222
rect 3789 1218 3790 1222
rect 3954 1218 3955 1222
rect 4045 1218 4046 1222
rect 4146 1218 4147 1222
rect 496 1203 498 1207
rect 502 1203 505 1207
rect 509 1203 512 1207
rect 1520 1203 1522 1207
rect 1526 1203 1529 1207
rect 1533 1203 1536 1207
rect 2544 1203 2546 1207
rect 2550 1203 2553 1207
rect 2557 1203 2560 1207
rect 3568 1203 3570 1207
rect 3574 1203 3577 1207
rect 3581 1203 3584 1207
rect 546 1188 547 1192
rect 1141 1188 1142 1192
rect 2122 1188 2123 1192
rect 2285 1188 2286 1192
rect 3658 1188 3659 1192
rect 4514 1188 4515 1192
rect 274 1168 281 1171
rect 1338 1168 1345 1171
rect 2474 1168 2481 1171
rect 3946 1168 3953 1171
rect 482 1158 486 1162
rect 494 1158 521 1161
rect 590 1151 593 1161
rect 1018 1158 1041 1161
rect 1082 1158 1086 1162
rect 1118 1161 1121 1168
rect 1110 1158 1121 1161
rect 1558 1158 1566 1161
rect 1782 1158 1801 1161
rect 2258 1158 2265 1161
rect 2922 1158 2926 1162
rect 3046 1158 3054 1161
rect 590 1148 609 1151
rect 614 1148 633 1151
rect 670 1151 673 1158
rect 3396 1157 3398 1161
rect 702 1152 706 1154
rect 670 1148 689 1151
rect 614 1142 617 1148
rect 1042 1148 1049 1151
rect 1298 1148 1305 1151
rect 1326 1148 1337 1151
rect 1362 1148 1369 1151
rect 1842 1148 1857 1151
rect 1898 1148 1905 1151
rect 2014 1151 2018 1154
rect 3454 1152 3457 1161
rect 3562 1158 3566 1162
rect 3582 1161 3585 1168
rect 3582 1158 3601 1161
rect 3698 1158 3705 1161
rect 3906 1158 3910 1162
rect 4062 1158 4070 1161
rect 1998 1148 2018 1151
rect 2058 1148 2073 1151
rect 1334 1142 1337 1148
rect 310 1138 318 1141
rect 530 1138 537 1141
rect 674 1138 681 1141
rect 770 1138 777 1141
rect 1014 1138 1030 1141
rect 1218 1138 1225 1141
rect 1394 1138 1409 1141
rect 1766 1141 1769 1148
rect 1758 1138 1769 1141
rect 1822 1138 1833 1141
rect 2078 1141 2081 1151
rect 2818 1148 2833 1151
rect 2938 1148 2945 1151
rect 3638 1148 3657 1151
rect 3898 1148 3905 1151
rect 4086 1151 4089 1161
rect 4022 1148 4049 1151
rect 4054 1148 4089 1151
rect 4270 1148 4278 1151
rect 4494 1148 4513 1151
rect 4530 1148 4537 1151
rect 4558 1151 4561 1161
rect 4554 1148 4561 1151
rect 2078 1138 2097 1141
rect 2162 1138 2169 1141
rect 2214 1141 2217 1148
rect 2214 1138 2225 1141
rect 2246 1138 2265 1141
rect 2294 1138 2302 1141
rect 2406 1141 2409 1148
rect 2398 1138 2409 1141
rect 2530 1138 2561 1141
rect 2670 1138 2689 1141
rect 2854 1138 2865 1141
rect 3078 1138 3089 1141
rect 3118 1138 3126 1141
rect 3186 1138 3193 1141
rect 3202 1138 3217 1141
rect 3370 1138 3377 1141
rect 3418 1138 3425 1141
rect 3614 1138 3630 1141
rect 3758 1141 3761 1148
rect 4494 1142 4497 1148
rect 3758 1138 3769 1141
rect 3814 1138 3833 1141
rect 3878 1138 3897 1141
rect 4082 1138 4089 1141
rect 4246 1138 4257 1141
rect 4310 1138 4318 1141
rect 4410 1138 4417 1141
rect 4470 1138 4478 1141
rect 1366 1128 1377 1131
rect 1406 1128 1409 1138
rect 1614 1128 1633 1131
rect 2022 1131 2025 1138
rect 2022 1128 2033 1131
rect 2166 1128 2169 1138
rect 3678 1132 3681 1138
rect 2210 1128 2214 1132
rect 2498 1128 2505 1131
rect 2574 1128 2593 1131
rect 2946 1128 2953 1131
rect 3678 1128 3686 1132
rect 301 1118 302 1122
rect 1554 1118 1555 1122
rect 2154 1118 2155 1122
rect 3010 1118 3011 1122
rect 3858 1118 3859 1122
rect 3933 1118 3934 1122
rect 4397 1118 4398 1122
rect 4485 1118 4486 1122
rect 1000 1103 1002 1107
rect 1006 1103 1009 1107
rect 1013 1103 1016 1107
rect 2024 1103 2026 1107
rect 2030 1103 2033 1107
rect 2037 1103 2040 1107
rect 3048 1103 3050 1107
rect 3054 1103 3057 1107
rect 3061 1103 3064 1107
rect 4080 1103 4082 1107
rect 4086 1103 4089 1107
rect 4093 1103 4096 1107
rect 413 1088 414 1092
rect 470 1088 478 1091
rect 1053 1088 1054 1092
rect 1629 1088 1630 1092
rect 2517 1088 2518 1092
rect 2550 1088 2558 1091
rect 2586 1088 2587 1092
rect 3685 1088 3686 1092
rect 4125 1088 4126 1092
rect 1494 1078 1505 1081
rect 1510 1078 1526 1081
rect 1806 1078 1817 1081
rect 1910 1078 1921 1081
rect 1958 1078 1969 1081
rect 270 1058 278 1061
rect 310 1061 313 1071
rect 490 1068 498 1071
rect 1002 1068 1017 1071
rect 1398 1068 1406 1071
rect 1446 1071 1449 1078
rect 1446 1068 1460 1071
rect 1566 1068 1582 1071
rect 1750 1071 1753 1078
rect 1718 1068 1737 1071
rect 1742 1068 1753 1071
rect 1990 1068 2009 1071
rect 306 1058 313 1061
rect 326 1058 345 1061
rect 950 1058 958 1061
rect 1166 1058 1177 1061
rect 1394 1058 1417 1061
rect 1514 1058 1537 1061
rect 1566 1058 1569 1068
rect 1938 1058 1945 1061
rect 1990 1058 1993 1068
rect 2014 1062 2017 1081
rect 2034 1078 2046 1081
rect 2742 1078 2753 1081
rect 2826 1078 2833 1081
rect 4050 1078 4057 1081
rect 4410 1078 4417 1081
rect 2198 1068 2214 1071
rect 2310 1068 2329 1071
rect 2342 1068 2350 1071
rect 2366 1068 2385 1071
rect 2526 1068 2534 1071
rect 2570 1068 2577 1071
rect 2594 1068 2601 1071
rect 2622 1068 2633 1071
rect 2894 1068 2902 1071
rect 3058 1068 3065 1071
rect 2374 1058 2382 1061
rect 2802 1058 2817 1061
rect 2846 1058 2857 1061
rect 3066 1058 3073 1061
rect 3122 1058 3129 1061
rect 3226 1058 3233 1061
rect 3310 1061 3313 1068
rect 3578 1068 3585 1071
rect 3742 1068 3753 1071
rect 3742 1062 3745 1068
rect 3270 1058 3289 1061
rect 3294 1058 3313 1061
rect 3430 1058 3438 1061
rect 3598 1058 3625 1061
rect 3630 1058 3646 1061
rect 3706 1058 3713 1061
rect 3754 1058 3761 1061
rect 3870 1061 3874 1064
rect 3854 1058 3874 1061
rect 3958 1061 3961 1071
rect 3998 1068 4017 1071
rect 4038 1068 4046 1071
rect 4422 1068 4433 1071
rect 3942 1058 3961 1061
rect 3974 1058 3982 1061
rect 4018 1058 4025 1061
rect 4062 1061 4065 1068
rect 4422 1062 4425 1068
rect 4062 1058 4089 1061
rect 4110 1058 4118 1061
rect 4446 1058 4454 1061
rect 4534 1058 4542 1061
rect 290 1048 294 1052
rect 342 1048 345 1058
rect 686 1056 690 1058
rect 1174 1052 1177 1058
rect 1246 1048 1257 1051
rect 1366 1048 1377 1051
rect 1434 1048 1441 1051
rect 2058 1048 2065 1051
rect 2266 1048 2270 1052
rect 2438 1048 2446 1051
rect 2798 1048 2801 1058
rect 3270 1052 3273 1058
rect 2978 1048 2985 1051
rect 3130 1048 3134 1052
rect 3794 1048 3798 1052
rect 3806 1048 3817 1051
rect 4214 1048 4233 1051
rect 787 1038 790 1042
rect 1389 1038 1390 1042
rect 2942 1038 2950 1041
rect 3101 1038 3102 1042
rect 3326 1038 3334 1041
rect 3426 1038 3427 1042
rect 3517 1038 3518 1042
rect 3762 1038 3763 1042
rect 4198 1038 4214 1041
rect 357 1028 358 1032
rect 694 1028 697 1038
rect 1202 1018 1203 1022
rect 1234 1018 1235 1022
rect 1418 1018 1419 1022
rect 1669 1018 1670 1022
rect 1781 1018 1782 1022
rect 2077 1018 2078 1022
rect 2426 1018 2427 1022
rect 2842 1018 2843 1022
rect 3202 1018 3203 1022
rect 3650 1018 3651 1022
rect 4498 1018 4499 1022
rect 496 1003 498 1007
rect 502 1003 505 1007
rect 509 1003 512 1007
rect 1520 1003 1522 1007
rect 1526 1003 1529 1007
rect 1533 1003 1536 1007
rect 2544 1003 2546 1007
rect 2550 1003 2553 1007
rect 2557 1003 2560 1007
rect 3568 1003 3570 1007
rect 3574 1003 3577 1007
rect 3581 1003 3584 1007
rect 157 988 158 992
rect 914 988 915 992
rect 1773 988 1774 992
rect 2205 988 2206 992
rect 2637 988 2638 992
rect 2794 988 2795 992
rect 2949 988 2950 992
rect 3341 988 3342 992
rect 3666 988 3667 992
rect 3754 988 3755 992
rect 4005 988 4006 992
rect 250 978 251 982
rect 458 968 459 972
rect 595 968 598 972
rect 678 968 689 971
rect 851 968 854 972
rect 2230 968 2238 971
rect 2253 968 2254 972
rect 3013 968 3014 972
rect 3157 968 3158 972
rect 3402 968 3403 972
rect 3722 968 3723 972
rect 262 958 273 961
rect 678 958 681 968
rect 702 953 706 958
rect 1322 957 1324 961
rect 30 951 34 953
rect 22 948 34 951
rect 134 948 153 951
rect 198 948 206 951
rect 226 948 249 951
rect 374 948 382 951
rect 450 948 457 951
rect 614 951 618 953
rect 234 938 241 941
rect 406 941 409 948
rect 614 948 633 951
rect 942 948 950 951
rect 1150 948 1166 951
rect 1334 948 1358 951
rect 1574 951 1577 961
rect 1662 958 1673 961
rect 1750 958 1761 961
rect 2290 958 2294 962
rect 2918 958 2937 961
rect 3574 958 3590 961
rect 3634 958 3638 962
rect 3914 958 3918 962
rect 1670 952 1673 958
rect 1558 948 1577 951
rect 1678 948 1686 951
rect 2242 948 2249 951
rect 2386 948 2393 951
rect 2466 948 2473 951
rect 2542 948 2566 951
rect 2638 948 2646 951
rect 406 938 425 941
rect 484 938 497 941
rect 774 938 786 941
rect 1046 938 1057 941
rect 1222 941 1225 948
rect 1222 938 1233 941
rect 1254 938 1265 941
rect 1410 938 1417 941
rect 1526 938 1550 941
rect 1598 938 1609 941
rect 1718 938 1726 941
rect 2126 941 2129 948
rect 2798 942 2801 951
rect 2814 948 2825 951
rect 3014 948 3033 951
rect 3142 951 3145 958
rect 3134 948 3145 951
rect 3158 948 3166 951
rect 3342 948 3350 951
rect 3446 948 3454 951
rect 3566 948 3601 951
rect 3926 951 3929 961
rect 3926 948 3945 951
rect 4018 948 4025 951
rect 4074 948 4105 951
rect 4110 948 4126 951
rect 4310 948 4337 951
rect 4482 948 4489 951
rect 4518 948 4537 951
rect 2822 942 2825 948
rect 3102 946 3106 948
rect 2126 938 2137 941
rect 2158 938 2166 941
rect 2238 938 2246 941
rect 2374 938 2382 941
rect 2494 938 2502 941
rect 2726 938 2750 941
rect 2890 938 2897 941
rect 3022 938 3030 941
rect 3114 938 3121 941
rect 3174 938 3177 948
rect 3214 938 3222 941
rect 3246 938 3265 941
rect 3294 938 3302 941
rect 3362 938 3369 941
rect 3798 938 3801 948
rect 3822 938 3830 941
rect 4014 938 4022 941
rect 4030 938 4049 941
rect 4070 938 4086 941
rect 4110 938 4113 948
rect 4154 938 4161 941
rect 4286 941 4289 948
rect 4262 938 4273 941
rect 4278 938 4289 941
rect 4342 941 4345 948
rect 4342 938 4353 941
rect 494 932 497 938
rect 170 928 177 931
rect 890 928 905 931
rect 966 928 974 931
rect 1294 928 1310 931
rect 1338 928 1345 931
rect 1390 928 1401 931
rect 2126 928 2137 931
rect 2374 928 2377 938
rect 2494 928 2497 938
rect 2662 928 2670 931
rect 3510 928 3521 931
rect 3594 928 3609 931
rect 3862 928 3873 931
rect 890 918 891 922
rect 1014 918 1030 921
rect 1274 918 1275 922
rect 1517 918 1518 922
rect 1909 918 1910 922
rect 1000 903 1002 907
rect 1006 903 1009 907
rect 1013 903 1016 907
rect 2024 903 2026 907
rect 2030 903 2033 907
rect 2037 903 2040 907
rect 3048 903 3050 907
rect 3054 903 3057 907
rect 3061 903 3064 907
rect 4080 903 4082 907
rect 4086 903 4089 907
rect 4093 903 4096 907
rect 234 888 235 892
rect 1030 888 1046 891
rect 1122 888 1123 892
rect 1250 888 1251 892
rect 2098 888 2099 892
rect 2970 888 2971 892
rect 3062 888 3070 891
rect 3405 888 3406 892
rect 1146 878 1153 881
rect 4350 878 4361 881
rect 4382 878 4393 881
rect 93 868 94 872
rect 242 868 254 871
rect 534 868 550 871
rect 1154 868 1161 871
rect 1482 868 1489 871
rect 1650 868 1657 871
rect 1686 868 1697 871
rect 1774 868 1793 871
rect 1982 868 2001 871
rect 2050 868 2057 871
rect 46 858 58 861
rect 1334 858 1350 861
rect 1470 858 1478 861
rect 1934 861 1937 868
rect 1926 858 1937 861
rect 1982 858 1985 868
rect 2158 868 2174 871
rect 2234 868 2241 871
rect 2258 868 2265 871
rect 2282 868 2289 871
rect 2310 862 2313 871
rect 2374 862 2377 871
rect 2386 868 2393 871
rect 2402 868 2409 871
rect 2434 868 2441 871
rect 2654 868 2673 871
rect 3082 868 3089 871
rect 3734 871 3737 878
rect 3726 868 3737 871
rect 3874 868 3881 871
rect 3926 868 3937 871
rect 3934 862 3937 868
rect 2106 858 2121 861
rect 2314 858 2329 861
rect 2414 858 2433 861
rect 2542 858 2577 861
rect 3102 858 3110 861
rect 3318 858 3337 861
rect 3570 858 3601 861
rect 3694 858 3713 861
rect 3730 858 3737 861
rect 3902 858 3921 861
rect 4006 861 4009 871
rect 4118 868 4126 871
rect 4310 868 4326 871
rect 4506 868 4529 871
rect 4562 868 4569 871
rect 4006 858 4022 861
rect 4062 858 4086 861
rect 4218 858 4225 861
rect 4430 858 4438 861
rect 4538 858 4545 861
rect 54 857 58 858
rect 718 856 722 858
rect 546 848 558 851
rect 554 838 569 841
rect 686 841 689 851
rect 1126 848 1137 851
rect 1254 848 1262 851
rect 1862 848 1873 851
rect 2622 848 2630 851
rect 2798 848 2817 851
rect 3158 848 3166 851
rect 3334 848 3337 858
rect 3694 852 3697 858
rect 3378 848 3382 852
rect 3558 848 3574 851
rect 3890 848 3894 852
rect 3902 848 3905 858
rect 3982 851 3985 858
rect 3974 848 3985 851
rect 4082 848 4097 851
rect 4478 848 4489 851
rect 678 838 689 841
rect 3221 838 3222 842
rect 566 828 569 838
rect 726 828 729 838
rect 3437 828 3438 832
rect 1370 818 1372 822
rect 1421 818 1422 822
rect 1453 818 1454 822
rect 1506 818 1508 822
rect 1706 818 1707 822
rect 2122 818 2123 822
rect 2330 818 2331 822
rect 2786 818 2787 822
rect 3133 818 3134 822
rect 4290 818 4291 822
rect 496 803 498 807
rect 502 803 505 807
rect 509 803 512 807
rect 1520 803 1522 807
rect 1526 803 1529 807
rect 1533 803 1536 807
rect 2544 803 2546 807
rect 2550 803 2553 807
rect 2557 803 2560 807
rect 3568 803 3570 807
rect 3574 803 3577 807
rect 3581 803 3584 807
rect 1242 788 1243 792
rect 1698 788 1699 792
rect 1813 788 1814 792
rect 2106 788 2107 792
rect 2138 788 2139 792
rect 2202 788 2203 792
rect 2834 788 2835 792
rect 3418 788 3419 792
rect 3549 788 3550 792
rect 3717 788 3718 792
rect 4429 788 4430 792
rect 301 768 302 772
rect 550 768 561 771
rect 558 762 561 768
rect 1958 768 1969 771
rect 1998 768 2006 771
rect 2933 768 2934 772
rect 3990 768 3998 771
rect 4114 768 4115 772
rect 4206 768 4222 771
rect 4261 768 4262 772
rect 4334 768 4350 771
rect 110 758 121 761
rect 130 758 134 762
rect 186 748 209 751
rect 246 748 254 751
rect 286 751 289 761
rect 270 748 289 751
rect 374 751 377 761
rect 374 748 393 751
rect 398 748 414 751
rect 438 748 446 751
rect 682 748 689 751
rect 806 751 810 753
rect 798 748 810 751
rect 222 738 225 748
rect 238 738 257 741
rect 498 738 529 741
rect 578 738 593 741
rect 606 738 617 741
rect 734 741 737 748
rect 934 748 950 751
rect 1086 751 1089 761
rect 1044 748 1073 751
rect 1086 748 1113 751
rect 1190 751 1193 761
rect 1350 761 1353 768
rect 1350 758 1361 761
rect 1466 758 1470 762
rect 1518 758 1545 761
rect 2150 758 2161 761
rect 2570 758 2577 761
rect 2758 758 2769 761
rect 2802 758 2809 761
rect 2914 758 2921 761
rect 3106 758 3110 762
rect 3118 758 3137 761
rect 1190 748 1206 751
rect 1214 748 1230 751
rect 1678 748 1694 751
rect 1850 748 1865 751
rect 1926 748 1945 751
rect 1950 748 1958 751
rect 2194 748 2201 751
rect 2350 748 2361 751
rect 2630 748 2641 751
rect 2698 748 2705 751
rect 2938 748 2953 751
rect 718 738 737 741
rect 894 738 906 741
rect 1070 738 1073 748
rect 1926 746 1930 748
rect 2950 742 2953 748
rect 2990 748 3001 751
rect 3194 748 3209 751
rect 3214 748 3222 751
rect 3346 748 3353 751
rect 3502 751 3505 761
rect 3502 748 3521 751
rect 3550 748 3585 751
rect 3766 751 3769 761
rect 4126 758 4137 761
rect 4174 758 4185 761
rect 3750 748 3769 751
rect 4078 748 4105 751
rect 4502 748 4513 751
rect 2990 742 2993 748
rect 1318 738 1326 741
rect 1346 738 1353 741
rect 1426 738 1441 741
rect 1494 738 1505 741
rect 1558 738 1574 741
rect 1830 738 1841 741
rect 2298 738 2305 741
rect 2350 738 2358 741
rect 2406 738 2425 741
rect 2706 738 2713 741
rect 3026 738 3041 741
rect 3046 738 3062 741
rect 3334 738 3342 741
rect 3462 738 3470 741
rect 3626 738 3633 741
rect 4102 742 4105 748
rect 3910 738 3918 741
rect 4038 738 4065 741
rect 4286 741 4289 748
rect 4270 738 4281 741
rect 4286 738 4297 741
rect 4366 738 4374 741
rect 4470 738 4473 748
rect 4514 738 4521 741
rect 4546 738 4553 741
rect 1086 732 1089 738
rect 1830 732 1833 738
rect 1082 728 1089 732
rect 1586 728 1596 731
rect 1670 728 1678 731
rect 2446 728 2457 731
rect 3066 728 3081 731
rect 4286 728 4297 731
rect 746 718 747 722
rect 770 718 771 722
rect 1124 718 1126 722
rect 1514 718 1515 722
rect 2066 718 2067 722
rect 2541 718 2542 722
rect 2690 718 2691 722
rect 2754 718 2755 722
rect 3162 718 3163 722
rect 3181 718 3182 722
rect 3389 718 3390 722
rect 4570 718 4572 722
rect 1000 703 1002 707
rect 1006 703 1009 707
rect 1013 703 1016 707
rect 2024 703 2026 707
rect 2030 703 2033 707
rect 2037 703 2040 707
rect 3048 703 3050 707
rect 3054 703 3057 707
rect 3061 703 3064 707
rect 4080 703 4082 707
rect 4086 703 4089 707
rect 4093 703 4096 707
rect 1292 688 1294 692
rect 2450 688 2451 692
rect 2501 688 2502 692
rect 2597 688 2598 692
rect 3178 688 3179 692
rect 3202 688 3203 692
rect 3341 688 3342 692
rect 3501 688 3502 692
rect 3557 688 3558 692
rect 3829 688 3830 692
rect 790 678 806 681
rect 790 674 794 678
rect 246 668 257 671
rect 482 668 489 671
rect 694 668 702 671
rect 862 668 874 671
rect 1014 668 1022 671
rect 62 658 70 661
rect 142 661 145 668
rect 246 662 249 668
rect 142 658 153 661
rect 502 658 518 661
rect 1126 662 1129 671
rect 1182 671 1185 681
rect 1190 678 1198 681
rect 1230 678 1249 681
rect 1178 668 1185 671
rect 1190 668 1209 671
rect 1254 671 1257 681
rect 1378 678 1393 681
rect 2038 678 2065 681
rect 2630 678 2649 681
rect 3902 678 3913 681
rect 4310 678 4318 681
rect 1254 668 1262 671
rect 1342 671 1345 678
rect 1326 668 1345 671
rect 1902 668 1921 671
rect 1998 668 2025 671
rect 922 658 929 661
rect 1206 658 1209 668
rect 2094 662 2097 671
rect 2186 668 2193 671
rect 2250 668 2257 671
rect 2326 668 2337 671
rect 2606 668 2614 671
rect 2658 668 2673 671
rect 2838 668 2846 671
rect 3126 668 3137 671
rect 3566 668 3590 671
rect 3766 668 3777 671
rect 3954 668 3961 671
rect 3966 668 3982 671
rect 4102 668 4110 671
rect 1338 658 1345 661
rect 1434 658 1460 661
rect 1822 658 1841 661
rect 2206 661 2210 664
rect 3134 662 3137 668
rect 3766 662 3769 668
rect 2190 658 2210 661
rect 2286 658 2305 661
rect 2346 658 2353 661
rect 2386 658 2398 661
rect 2534 658 2558 661
rect 2578 658 2593 661
rect 2610 658 2617 661
rect 2634 658 2641 661
rect 3302 658 3321 661
rect 3390 658 3409 661
rect 3446 658 3465 661
rect 3534 658 3553 661
rect 3670 658 3689 661
rect 3790 658 3798 661
rect 3926 658 3934 661
rect 3942 658 3950 661
rect 4142 658 4150 661
rect 4378 658 4385 661
rect 4438 661 4441 671
rect 4438 658 4457 661
rect 4502 661 4505 671
rect 4494 658 4505 661
rect 766 641 769 651
rect 1822 648 1825 658
rect 1886 648 1894 651
rect 2302 648 2305 658
rect 2406 648 2417 651
rect 2546 648 2561 651
rect 2590 648 2593 658
rect 2826 648 2830 652
rect 3302 648 3305 658
rect 3406 648 3409 658
rect 3462 648 3465 658
rect 3550 652 3553 658
rect 3514 648 3521 651
rect 3686 648 3689 658
rect 4494 656 4498 658
rect 4178 648 4182 652
rect 4450 648 4457 651
rect 766 638 777 641
rect 1694 638 1706 641
rect 1717 638 1718 642
rect 1922 638 1929 641
rect 3646 638 3654 641
rect 1950 628 1953 638
rect 1349 618 1350 622
rect 1506 618 1507 622
rect 2530 618 2531 622
rect 2573 618 2574 622
rect 2954 618 2955 622
rect 3741 618 3742 622
rect 4061 618 4062 622
rect 4130 618 4131 622
rect 4574 618 4582 621
rect 496 603 498 607
rect 502 603 505 607
rect 509 603 512 607
rect 1520 603 1522 607
rect 1526 603 1529 607
rect 1533 603 1536 607
rect 2544 603 2546 607
rect 2550 603 2553 607
rect 2557 603 2560 607
rect 3568 603 3570 607
rect 3574 603 3577 607
rect 3581 603 3584 607
rect 530 588 532 592
rect 1866 588 1867 592
rect 1978 588 1979 592
rect 2058 588 2059 592
rect 2253 588 2254 592
rect 2442 588 2443 592
rect 2618 588 2619 592
rect 2874 588 2875 592
rect 3317 588 3318 592
rect 3397 588 3398 592
rect 3453 588 3454 592
rect 3546 588 3547 592
rect 4013 588 4014 592
rect 4245 588 4246 592
rect 4541 588 4542 592
rect 4573 588 4574 592
rect 74 568 77 572
rect 238 568 249 571
rect 246 561 249 568
rect 797 568 798 572
rect 866 568 881 571
rect 886 568 902 571
rect 1444 568 1446 572
rect 1490 568 1506 571
rect 1782 568 1793 571
rect 1894 568 1929 571
rect 2341 568 2342 572
rect 2750 568 2761 571
rect 3846 568 3857 571
rect 4394 568 4395 572
rect 254 561 257 568
rect 1502 566 1506 568
rect 1790 562 1793 568
rect 2758 562 2761 568
rect 3854 562 3857 568
rect 246 558 257 561
rect 54 551 58 553
rect 782 552 785 561
rect 46 548 58 551
rect 722 548 729 551
rect 1018 548 1025 551
rect 142 538 154 541
rect 774 541 777 548
rect 1574 551 1577 561
rect 1574 548 1593 551
rect 1670 551 1673 561
rect 1654 548 1673 551
rect 1702 551 1705 558
rect 1694 548 1705 551
rect 1774 551 1777 561
rect 1762 548 1777 551
rect 1794 548 1809 551
rect 1934 551 1937 561
rect 2070 558 2078 561
rect 2370 558 2374 562
rect 2486 558 2494 561
rect 2514 558 2521 561
rect 2886 558 2905 561
rect 3042 558 3046 562
rect 3054 558 3089 561
rect 3178 558 3182 562
rect 1934 548 1953 551
rect 1958 548 1969 551
rect 2002 548 2009 551
rect 2070 548 2089 551
rect 2162 548 2169 551
rect 2254 548 2262 551
rect 2342 548 2358 551
rect 2422 548 2433 551
rect 2454 551 2457 558
rect 2454 548 2465 551
rect 2478 548 2486 551
rect 2514 548 2529 551
rect 2670 548 2686 551
rect 2998 551 3002 554
rect 2998 548 3017 551
rect 3158 548 3166 551
rect 3254 548 3262 551
rect 3374 551 3377 561
rect 3374 548 3382 551
rect 3398 548 3406 551
rect 3438 551 3441 561
rect 3510 558 3518 561
rect 3422 548 3441 551
rect 3502 548 3510 551
rect 3558 551 3561 561
rect 3630 551 3633 561
rect 4430 558 4438 561
rect 3558 548 3593 551
rect 3614 548 3633 551
rect 3866 548 3873 551
rect 3966 548 3990 551
rect 702 538 721 541
rect 766 538 777 541
rect 1350 541 1353 548
rect 1350 538 1361 541
rect 1606 538 1617 541
rect 1694 538 1697 548
rect 1790 538 1793 548
rect 1966 542 1969 548
rect 2390 546 2394 548
rect 2430 538 2433 548
rect 2462 538 2465 548
rect 2590 538 2606 541
rect 2654 541 2657 548
rect 2646 538 2657 541
rect 2694 538 2713 541
rect 2758 538 2766 541
rect 2846 538 2854 541
rect 3074 538 3081 541
rect 3326 538 3337 541
rect 3462 538 3470 541
rect 3526 538 3537 541
rect 3738 538 3745 541
rect 3750 538 3777 541
rect 3834 538 3849 541
rect 3886 538 3918 541
rect 4110 541 4113 548
rect 4086 538 4113 541
rect 4158 538 4166 541
rect 4190 541 4193 551
rect 4310 548 4318 551
rect 4386 548 4393 551
rect 4422 548 4430 551
rect 4466 548 4473 551
rect 4530 548 4537 551
rect 4190 538 4198 541
rect 4334 538 4353 541
rect 4378 538 4385 541
rect 4474 538 4481 541
rect 2574 531 2577 538
rect 2546 528 2561 531
rect 2566 528 2577 531
rect 3734 528 3737 538
rect 4114 528 4121 531
rect 4350 528 4353 538
rect 4510 531 4513 538
rect 4510 528 4521 531
rect 4526 528 4534 531
rect 285 518 286 522
rect 850 518 852 522
rect 1509 518 1510 522
rect 1709 518 1710 522
rect 2925 518 2926 522
rect 1000 503 1002 507
rect 1006 503 1009 507
rect 1013 503 1016 507
rect 2024 503 2026 507
rect 2030 503 2033 507
rect 2037 503 2040 507
rect 3048 503 3050 507
rect 3054 503 3057 507
rect 3061 503 3064 507
rect 4080 503 4082 507
rect 4086 503 4089 507
rect 4093 503 4096 507
rect 717 488 718 492
rect 1434 488 1435 492
rect 1658 488 1659 492
rect 2082 488 2083 492
rect 2205 488 2206 492
rect 2837 488 2838 492
rect 3221 488 3222 492
rect 3277 488 3278 492
rect 3381 488 3382 492
rect 3901 488 3902 492
rect 4005 488 4006 492
rect 4314 488 4315 492
rect 4397 488 4398 492
rect 4445 488 4446 492
rect 4549 488 4550 492
rect 626 478 630 482
rect 3046 478 3062 481
rect 318 468 329 471
rect 550 468 558 471
rect 726 468 734 471
rect 2098 468 2105 471
rect 2150 468 2158 471
rect 2310 468 2329 471
rect 2350 468 2369 471
rect 2390 468 2398 471
rect 2426 468 2438 471
rect 2662 468 2670 471
rect 2722 468 2729 471
rect 3086 471 3089 481
rect 3858 478 3865 481
rect 4122 478 4129 481
rect 4254 478 4262 482
rect 4254 472 4257 478
rect 3086 468 3094 471
rect 3526 468 3542 471
rect 3606 468 3617 471
rect 3622 468 3641 471
rect 3726 468 3737 471
rect 3990 468 4001 471
rect 4182 468 4190 471
rect 4294 471 4297 481
rect 4294 468 4302 471
rect 4462 471 4465 478
rect 4454 468 4465 471
rect 4470 468 4497 471
rect 4558 468 4569 471
rect 318 462 321 468
rect 526 458 545 461
rect 742 458 761 461
rect 486 448 513 451
rect 878 448 881 458
rect 966 448 982 451
rect 1438 448 1441 468
rect 1450 458 1457 461
rect 1530 458 1572 461
rect 1638 458 1646 461
rect 1682 458 1689 461
rect 1826 458 1833 461
rect 1838 458 1857 461
rect 1910 458 1929 461
rect 1966 458 1985 461
rect 2130 458 2137 461
rect 2150 458 2169 461
rect 2246 458 2254 461
rect 2430 458 2449 461
rect 2538 458 2577 461
rect 2666 458 2673 461
rect 2798 458 2806 461
rect 2814 458 2830 461
rect 2854 461 2858 464
rect 3622 462 3625 468
rect 3998 462 4001 468
rect 2838 458 2858 461
rect 3150 458 3169 461
rect 3414 458 3430 461
rect 3530 458 3545 461
rect 3570 458 3593 461
rect 3634 458 3641 461
rect 3686 458 3705 461
rect 4078 458 4113 461
rect 4218 458 4225 461
rect 4286 458 4294 461
rect 4518 461 4521 468
rect 4518 458 4529 461
rect 4558 458 4569 461
rect 1810 448 1814 452
rect 1854 448 1857 458
rect 1910 448 1913 458
rect 1966 448 1969 458
rect 2062 448 2070 451
rect 2086 448 2105 451
rect 2150 448 2153 458
rect 2190 448 2201 451
rect 2970 448 2974 452
rect 3150 448 3153 458
rect 3542 448 3545 458
rect 3550 448 3585 451
rect 3702 448 3705 458
rect 3994 448 4001 451
rect 4202 448 4206 452
rect 4222 448 4225 458
rect 4558 452 4561 458
rect 470 438 478 441
rect 893 438 894 442
rect 930 438 945 441
rect 1155 438 1158 442
rect 2730 438 2737 441
rect 269 428 270 432
rect 694 428 697 438
rect 1402 418 1403 422
rect 1698 418 1699 422
rect 1757 418 1758 422
rect 2610 418 2611 422
rect 2653 418 2654 422
rect 3717 418 3718 422
rect 4037 418 4038 422
rect 4173 418 4174 422
rect 4237 418 4238 422
rect 496 403 498 407
rect 502 403 505 407
rect 509 403 512 407
rect 1520 403 1522 407
rect 1526 403 1529 407
rect 1533 403 1536 407
rect 2544 403 2546 407
rect 2550 403 2553 407
rect 2557 403 2560 407
rect 3568 403 3570 407
rect 3574 403 3577 407
rect 3581 403 3584 407
rect 730 388 731 392
rect 1526 388 1534 391
rect 1789 388 1790 392
rect 1821 388 1822 392
rect 1850 388 1851 392
rect 2029 388 2030 392
rect 2077 388 2078 392
rect 2133 388 2134 392
rect 2349 388 2350 392
rect 2426 388 2427 392
rect 2650 388 2651 392
rect 2765 388 2766 392
rect 2890 388 2891 392
rect 2946 388 2947 392
rect 2994 388 2995 392
rect 3029 388 3030 392
rect 3077 388 3078 392
rect 3114 388 3115 392
rect 3266 388 3267 392
rect 3306 388 3307 392
rect 3365 388 3366 392
rect 3418 388 3419 392
rect 3453 388 3454 392
rect 3610 388 3611 392
rect 3669 388 3670 392
rect 3933 388 3934 392
rect 4042 388 4043 392
rect 4341 388 4342 392
rect 4562 388 4563 392
rect 77 378 78 382
rect 1666 378 1668 382
rect 294 368 310 371
rect 330 368 331 372
rect 2238 368 2250 371
rect 2261 368 2262 372
rect 3798 368 3825 371
rect 54 358 65 361
rect 306 358 313 361
rect 1610 358 1612 362
rect 1766 358 1777 361
rect 34 348 41 351
rect 82 348 105 351
rect 226 348 233 351
rect 494 348 529 351
rect 534 348 550 351
rect 566 348 577 351
rect 650 348 665 351
rect 746 348 761 351
rect 86 338 94 341
rect 126 341 129 348
rect 126 338 137 341
rect 142 338 153 341
rect 190 338 201 341
rect 494 338 497 348
rect 566 342 569 348
rect 1034 348 1041 351
rect 1426 348 1433 351
rect 1558 348 1569 351
rect 1830 348 1846 351
rect 1894 348 1905 351
rect 1922 348 1929 351
rect 1946 348 1961 351
rect 2030 348 2046 351
rect 2398 348 2425 351
rect 2450 348 2457 351
rect 2502 351 2505 361
rect 2502 348 2553 351
rect 2606 348 2614 351
rect 2662 348 2673 351
rect 2702 348 2710 351
rect 2902 351 2905 361
rect 2902 348 2921 351
rect 2938 348 2945 351
rect 2974 348 2993 351
rect 3082 348 3086 351
rect 3090 348 3097 351
rect 3126 348 3134 351
rect 3326 351 3329 361
rect 3334 358 3353 361
rect 3742 352 3745 361
rect 3310 348 3329 351
rect 3454 348 3462 351
rect 3574 348 3609 351
rect 3670 348 3678 351
rect 3726 348 3742 351
rect 3918 351 3921 361
rect 1566 342 1569 348
rect 710 338 721 341
rect 770 338 777 341
rect 958 338 986 341
rect 1418 338 1425 341
rect 1830 338 1833 348
rect 2662 342 2665 348
rect 1942 338 1950 341
rect 2038 338 2054 341
rect 2270 338 2278 341
rect 2302 338 2310 341
rect 2374 338 2382 341
rect 2614 338 2625 341
rect 2774 338 2782 341
rect 2926 338 2934 341
rect 3474 338 3481 341
rect 3594 338 3601 341
rect 3838 338 3841 348
rect 3894 341 3897 351
rect 3902 348 3921 351
rect 3934 348 3942 351
rect 4270 348 4281 351
rect 4346 348 4369 351
rect 4406 348 4414 351
rect 4486 348 4497 351
rect 4510 348 4521 351
rect 4542 348 4561 351
rect 4270 342 4273 348
rect 4494 342 4497 348
rect 4542 346 4546 348
rect 3878 338 3897 341
rect 4378 338 4385 341
rect 4438 338 4457 341
rect 22 332 25 338
rect 198 332 201 338
rect 18 328 25 332
rect 158 328 166 331
rect 1422 328 1425 338
rect 4006 332 4009 338
rect 1558 328 1569 331
rect 3394 328 3398 332
rect 4006 328 4014 332
rect 2573 318 2574 322
rect 3514 318 3515 322
rect 3533 318 3534 322
rect 1000 303 1002 307
rect 1006 303 1009 307
rect 1013 303 1016 307
rect 2024 303 2026 307
rect 2030 303 2033 307
rect 2037 303 2040 307
rect 3048 303 3050 307
rect 3054 303 3057 307
rect 3061 303 3064 307
rect 4080 303 4082 307
rect 4086 303 4089 307
rect 4093 303 4096 307
rect 330 288 331 292
rect 756 288 758 292
rect 1690 288 1692 292
rect 1914 288 1915 292
rect 2101 288 2102 292
rect 2165 288 2166 292
rect 2226 288 2227 292
rect 2845 288 2846 292
rect 2954 288 2955 292
rect 3054 288 3070 291
rect 3085 288 3086 292
rect 3109 288 3110 292
rect 3266 288 3267 292
rect 3482 288 3483 292
rect 3570 288 3571 292
rect 3981 288 3982 292
rect 4402 288 4409 291
rect 506 278 529 281
rect 622 278 630 282
rect 1834 278 1838 282
rect 2058 278 2065 281
rect 2342 278 2350 281
rect 622 272 625 278
rect 1494 276 1498 278
rect 3758 272 3761 281
rect 266 268 276 271
rect 666 268 673 271
rect 1084 268 1086 272
rect 1758 268 1769 271
rect 1814 268 1822 271
rect 1850 268 1873 271
rect 1982 268 1990 271
rect 2074 268 2081 271
rect 2274 268 2281 271
rect 2426 268 2433 271
rect 2962 268 2977 271
rect 3118 268 3126 271
rect 3374 268 3382 271
rect 3762 268 3769 271
rect 3858 268 3865 271
rect 3902 268 3921 271
rect 4294 268 4313 271
rect 4322 268 4337 271
rect 4358 268 4369 271
rect 174 258 193 261
rect 414 258 433 261
rect 446 258 473 261
rect 490 258 497 261
rect 562 258 569 261
rect 574 258 601 261
rect 646 258 657 261
rect 686 258 694 261
rect 862 258 881 261
rect 190 248 193 258
rect 238 241 241 248
rect 254 241 257 251
rect 310 248 313 258
rect 398 248 406 251
rect 430 248 433 258
rect 558 248 561 258
rect 646 252 649 258
rect 694 248 713 251
rect 878 248 881 258
rect 922 248 926 252
rect 958 242 961 261
rect 990 258 1006 261
rect 1718 261 1721 268
rect 1718 258 1729 261
rect 1898 258 1905 261
rect 2010 258 2017 261
rect 2050 258 2057 261
rect 2138 258 2153 261
rect 2234 258 2249 261
rect 2458 258 2473 261
rect 2514 258 2521 261
rect 2590 258 2606 261
rect 3166 258 3190 261
rect 3218 258 3225 261
rect 3278 258 3297 261
rect 3434 258 3441 261
rect 3486 258 3505 261
rect 3626 258 3641 261
rect 3646 258 3662 261
rect 3738 258 3745 261
rect 3782 258 3809 261
rect 3918 258 3921 268
rect 4358 262 4361 268
rect 3926 258 3934 261
rect 4074 258 4097 261
rect 4246 258 4265 261
rect 4442 258 4454 261
rect 4546 258 4553 261
rect 1102 256 1106 258
rect 1786 248 1788 252
rect 2014 248 2017 258
rect 3294 252 3297 258
rect 2690 248 2697 251
rect 2874 248 2878 252
rect 3058 248 3081 251
rect 3438 248 3441 258
rect 3486 252 3489 258
rect 4246 252 4249 258
rect 3574 248 3590 251
rect 3622 248 3630 251
rect 3642 248 3646 252
rect 4266 248 4270 252
rect 238 238 257 241
rect 797 238 798 242
rect 893 238 894 242
rect 205 228 206 232
rect 298 218 299 222
rect 386 218 387 222
rect 496 203 498 207
rect 502 203 505 207
rect 509 203 512 207
rect 1520 203 1522 207
rect 1526 203 1529 207
rect 1533 203 1536 207
rect 2544 203 2546 207
rect 2550 203 2553 207
rect 2557 203 2560 207
rect 3568 203 3570 207
rect 3574 203 3577 207
rect 3581 203 3584 207
rect 658 188 659 192
rect 2442 188 2443 192
rect 2538 188 2539 192
rect 2637 188 2638 192
rect 2677 188 2678 192
rect 2842 188 2843 192
rect 2962 188 2963 192
rect 3045 188 3046 192
rect 3090 188 3091 192
rect 3125 188 3126 192
rect 3298 188 3299 192
rect 3365 188 3366 192
rect 3677 188 3678 192
rect 3770 188 3771 192
rect 4106 188 4107 192
rect 4242 188 4243 192
rect 4314 188 4315 192
rect 4341 188 4342 192
rect 4458 188 4459 192
rect 4498 188 4499 192
rect 238 172 241 181
rect 570 178 571 182
rect 3941 178 3942 182
rect 2773 168 2774 172
rect 3170 168 3177 171
rect 3470 168 3490 171
rect 3810 168 3817 171
rect 4062 168 4086 171
rect 4370 168 4371 172
rect 230 152 234 154
rect 358 152 362 154
rect 542 148 561 151
rect 670 151 673 161
rect 838 152 842 154
rect 958 152 962 154
rect 670 148 689 151
rect 558 142 561 148
rect 718 141 721 148
rect 906 148 913 151
rect 1034 148 1041 151
rect 1142 148 1169 151
rect 1190 151 1193 161
rect 1226 158 1233 161
rect 1190 148 1209 151
rect 718 138 729 141
rect 886 138 905 141
rect 1166 138 1169 148
rect 1298 148 1305 151
rect 1434 148 1449 151
rect 2022 151 2025 161
rect 2174 158 2193 161
rect 2202 158 2206 162
rect 2286 158 2305 161
rect 2022 148 2057 151
rect 2066 148 2073 151
rect 2270 148 2289 151
rect 2378 148 2393 151
rect 2502 151 2505 161
rect 2550 158 2558 161
rect 2854 158 2873 161
rect 3266 158 3270 162
rect 2498 148 2505 151
rect 2510 148 2529 151
rect 2554 148 2585 151
rect 2710 148 2718 151
rect 2742 148 2750 151
rect 3046 148 3054 151
rect 3310 151 3313 161
rect 3454 158 3465 161
rect 3290 148 3297 151
rect 3310 148 3329 151
rect 3386 148 3393 151
rect 3490 148 3497 151
rect 3502 148 3518 151
rect 3582 148 3590 151
rect 1218 138 1225 141
rect 1478 138 1506 141
rect 1990 138 2001 141
rect 2214 138 2225 141
rect 2326 138 2345 141
rect 2526 138 2529 148
rect 2722 138 2729 141
rect 2822 138 2833 141
rect 2950 138 2953 148
rect 3054 138 3062 141
rect 3158 138 3166 141
rect 3462 141 3465 148
rect 3446 138 3465 141
rect 3646 141 3649 151
rect 3990 151 3993 161
rect 3986 148 3993 151
rect 4082 148 4105 151
rect 4122 148 4129 151
rect 4166 151 4169 161
rect 4162 148 4169 151
rect 4182 148 4190 151
rect 4382 151 4385 158
rect 4362 148 4369 151
rect 4382 148 4393 151
rect 4430 148 4438 151
rect 4474 148 4497 151
rect 3646 138 3665 141
rect 3742 138 3750 141
rect 3802 138 3809 141
rect 4130 138 4137 141
rect 4290 138 4313 141
rect 4482 138 4489 141
rect 546 128 561 131
rect 742 131 746 133
rect 706 128 713 131
rect 718 128 729 131
rect 734 128 746 131
rect 3006 128 3017 131
rect 3565 128 3566 132
rect 3754 128 3761 131
rect 978 118 985 121
rect 2141 118 2142 122
rect 1000 103 1002 107
rect 1006 103 1009 107
rect 1013 103 1016 107
rect 2024 103 2026 107
rect 2030 103 2033 107
rect 2037 103 2040 107
rect 3048 103 3050 107
rect 3054 103 3057 107
rect 3061 103 3064 107
rect 4080 103 4082 107
rect 4086 103 4089 107
rect 4093 103 4096 107
rect 522 88 529 91
rect 1518 88 1526 91
rect 1930 88 1931 92
rect 2205 88 2206 92
rect 2613 88 2614 92
rect 3445 88 3446 92
rect 3574 88 3590 91
rect 3669 88 3670 92
rect 1650 78 1666 81
rect 1958 78 1969 81
rect 182 68 185 78
rect 1662 74 1666 78
rect 1838 68 1849 71
rect 238 58 250 61
rect 502 58 518 61
rect 578 58 585 61
rect 1230 58 1241 61
rect 1294 58 1310 61
rect 1350 58 1361 61
rect 1530 58 1545 61
rect 1870 62 1873 71
rect 1878 68 1897 71
rect 2166 71 2169 81
rect 3142 78 3153 81
rect 3258 78 3265 81
rect 3482 78 3489 81
rect 3630 78 3641 81
rect 3646 78 3654 81
rect 3698 78 3705 82
rect 4346 78 4353 81
rect 4358 78 4366 81
rect 4374 78 4385 81
rect 3142 72 3145 78
rect 3702 72 3705 78
rect 4374 72 4377 78
rect 2150 68 2169 71
rect 2342 68 2353 71
rect 2406 68 2414 71
rect 2538 68 2561 71
rect 2742 68 2753 71
rect 2838 68 2846 71
rect 2934 68 2945 71
rect 3198 68 3206 71
rect 3238 68 3254 71
rect 3322 68 3329 71
rect 3554 68 3561 71
rect 3630 68 3641 71
rect 3682 68 3689 71
rect 4330 68 4337 71
rect 4494 68 4513 71
rect 1774 58 1790 61
rect 1934 58 1942 61
rect 1982 61 1985 68
rect 1966 58 1985 61
rect 2082 58 2089 61
rect 2150 58 2158 61
rect 2190 58 2209 61
rect 2278 58 2286 61
rect 2290 58 2297 61
rect 2446 58 2454 61
rect 2538 58 2558 61
rect 2802 58 2809 61
rect 2846 61 2849 68
rect 3638 62 3641 68
rect 2846 58 2865 61
rect 2946 58 2953 61
rect 3074 58 3081 61
rect 3246 58 3257 61
rect 3370 58 3377 61
rect 3426 58 3433 61
rect 3658 58 3665 61
rect 3838 58 3846 61
rect 3938 58 3945 61
rect 4478 61 4481 68
rect 4422 58 4441 61
rect 4462 58 4481 61
rect 4494 62 4497 68
rect 4562 58 4569 61
rect 246 57 250 58
rect 1230 57 1234 58
rect 1350 57 1354 58
rect 1774 57 1778 58
rect 1934 48 1937 58
rect 2294 48 2297 58
rect 2302 48 2321 51
rect 2494 48 2513 51
rect 2522 48 2526 52
rect 2602 48 2609 51
rect 2654 48 2673 51
rect 2774 48 2793 51
rect 2878 48 2897 51
rect 2954 48 2958 52
rect 3030 48 3038 51
rect 3070 51 3073 58
rect 3246 52 3249 58
rect 3054 48 3073 51
rect 3374 48 3377 58
rect 3402 48 3409 51
rect 3662 48 3665 58
rect 4070 51 4073 58
rect 4070 48 4081 51
rect 4422 48 4425 58
rect 2022 38 2030 41
rect 2333 38 2334 42
rect 3802 38 3803 42
rect 4570 38 4571 42
rect 4490 28 4491 32
rect 3085 18 3086 22
rect 4053 18 4054 22
rect 496 3 498 7
rect 502 3 505 7
rect 509 3 512 7
rect 1520 3 1522 7
rect 1526 3 1529 7
rect 1533 3 1536 7
rect 2544 3 2546 7
rect 2550 3 2553 7
rect 2557 3 2560 7
rect 3568 3 3570 7
rect 3574 3 3577 7
rect 3581 3 3584 7
<< m2contact >>
rect 498 4403 502 4407
rect 505 4403 509 4407
rect 1522 4403 1526 4407
rect 1529 4403 1533 4407
rect 2546 4403 2550 4407
rect 2553 4403 2557 4407
rect 3570 4403 3574 4407
rect 3577 4403 3581 4407
rect 2270 4388 2274 4392
rect 2742 4388 2746 4392
rect 2766 4388 2770 4392
rect 3126 4388 3130 4392
rect 3150 4388 3154 4392
rect 3190 4388 3194 4392
rect 3214 4388 3218 4392
rect 3294 4388 3298 4392
rect 3318 4388 3322 4392
rect 3374 4388 3378 4392
rect 3398 4388 3402 4392
rect 3454 4388 3458 4392
rect 3526 4388 3530 4392
rect 2030 4378 2034 4382
rect 3862 4378 3866 4382
rect 4046 4378 4050 4382
rect 1918 4368 1922 4372
rect 3014 4368 3018 4372
rect 3134 4368 3138 4372
rect 3182 4368 3186 4372
rect 3206 4368 3210 4372
rect 3438 4368 3442 4372
rect 3494 4368 3498 4372
rect 3598 4368 3602 4372
rect 3622 4368 3626 4372
rect 4198 4368 4202 4372
rect 38 4357 42 4361
rect 630 4358 634 4362
rect 654 4358 658 4362
rect 774 4358 778 4362
rect 790 4358 794 4362
rect 926 4358 930 4362
rect 1510 4358 1514 4362
rect 1542 4358 1546 4362
rect 1742 4358 1746 4362
rect 1774 4358 1778 4362
rect 2150 4358 2154 4362
rect 2190 4358 2194 4362
rect 2246 4358 2250 4362
rect 2342 4358 2346 4362
rect 2414 4358 2418 4362
rect 2454 4358 2458 4362
rect 2526 4358 2530 4362
rect 2606 4358 2610 4362
rect 2678 4358 2682 4362
rect 2702 4358 2706 4362
rect 2966 4358 2970 4362
rect 3246 4358 3250 4362
rect 3302 4358 3306 4362
rect 3342 4358 3346 4362
rect 3422 4358 3426 4362
rect 3478 4358 3482 4362
rect 3558 4358 3562 4362
rect 70 4348 74 4352
rect 118 4348 122 4352
rect 190 4347 194 4351
rect 286 4347 290 4351
rect 550 4347 554 4351
rect 694 4348 698 4352
rect 726 4348 730 4352
rect 734 4348 738 4352
rect 774 4348 778 4352
rect 790 4348 794 4352
rect 854 4348 858 4352
rect 926 4348 930 4352
rect 942 4348 946 4352
rect 982 4348 986 4352
rect 1070 4347 1074 4351
rect 1158 4348 1162 4352
rect 1222 4347 1226 4351
rect 1318 4347 1322 4351
rect 1422 4348 1426 4352
rect 1518 4348 1522 4352
rect 1638 4348 1642 4352
rect 1686 4348 1690 4352
rect 1702 4348 1706 4352
rect 1726 4348 1730 4352
rect 1742 4348 1746 4352
rect 1758 4348 1762 4352
rect 1886 4347 1890 4351
rect 1982 4347 1986 4351
rect 2094 4347 2098 4351
rect 2166 4348 2170 4352
rect 2254 4348 2258 4352
rect 2302 4348 2306 4352
rect 2310 4348 2314 4352
rect 2422 4348 2426 4352
rect 2758 4348 2762 4352
rect 2782 4348 2786 4352
rect 2822 4348 2826 4352
rect 2990 4348 2994 4352
rect 3086 4348 3090 4352
rect 3142 4348 3146 4352
rect 3174 4348 3178 4352
rect 3198 4348 3202 4352
rect 3254 4348 3258 4352
rect 3262 4348 3266 4352
rect 3270 4348 3274 4352
rect 3334 4348 3338 4352
rect 3358 4348 3362 4352
rect 3390 4348 3394 4352
rect 3414 4348 3418 4352
rect 3430 4348 3434 4352
rect 3446 4348 3450 4352
rect 3470 4348 3474 4352
rect 3486 4348 3490 4352
rect 3502 4348 3506 4352
rect 3510 4348 3514 4352
rect 3542 4348 3546 4352
rect 3710 4358 3714 4362
rect 3918 4358 3922 4362
rect 3942 4358 3946 4362
rect 3958 4358 3962 4362
rect 3974 4358 3978 4362
rect 3990 4358 3994 4362
rect 4022 4358 4026 4362
rect 3598 4348 3602 4352
rect 3638 4348 3642 4352
rect 3654 4348 3658 4352
rect 3670 4348 3674 4352
rect 3702 4348 3706 4352
rect 3734 4348 3738 4352
rect 3750 4348 3754 4352
rect 3766 4348 3770 4352
rect 3782 4348 3786 4352
rect 3806 4348 3810 4352
rect 3814 4348 3818 4352
rect 3830 4348 3834 4352
rect 3846 4348 3850 4352
rect 3894 4348 3898 4352
rect 3926 4348 3930 4352
rect 3942 4348 3946 4352
rect 3974 4348 3978 4352
rect 4006 4348 4010 4352
rect 4062 4358 4066 4362
rect 4158 4358 4162 4362
rect 4214 4358 4218 4362
rect 4278 4358 4282 4362
rect 4366 4358 4370 4362
rect 4438 4358 4442 4362
rect 4566 4358 4570 4362
rect 4046 4348 4050 4352
rect 4118 4348 4122 4352
rect 4150 4348 4154 4352
rect 4174 4348 4178 4352
rect 4198 4348 4202 4352
rect 4214 4348 4218 4352
rect 4246 4348 4250 4352
rect 4262 4348 4266 4352
rect 4278 4348 4282 4352
rect 4294 4348 4298 4352
rect 4302 4348 4306 4352
rect 4326 4348 4330 4352
rect 4342 4348 4346 4352
rect 4358 4348 4362 4352
rect 4382 4348 4386 4352
rect 4398 4348 4402 4352
rect 4414 4348 4418 4352
rect 4430 4348 4434 4352
rect 4454 4348 4458 4352
rect 4470 4348 4474 4352
rect 4494 4348 4498 4352
rect 4518 4348 4522 4352
rect 4542 4348 4546 4352
rect 4582 4348 4586 4352
rect 22 4338 26 4342
rect 62 4338 66 4342
rect 110 4338 114 4342
rect 270 4338 274 4342
rect 358 4338 362 4342
rect 406 4338 410 4342
rect 414 4338 418 4342
rect 462 4338 466 4342
rect 542 4338 546 4342
rect 590 4338 594 4342
rect 614 4338 618 4342
rect 638 4338 642 4342
rect 670 4338 674 4342
rect 694 4338 698 4342
rect 710 4338 714 4342
rect 742 4338 746 4342
rect 766 4338 770 4342
rect 846 4338 850 4342
rect 950 4338 954 4342
rect 974 4338 978 4342
rect 1086 4338 1090 4342
rect 6 4328 10 4332
rect 78 4328 82 4332
rect 126 4328 130 4332
rect 158 4328 162 4332
rect 190 4328 194 4332
rect 582 4328 586 4332
rect 702 4328 706 4332
rect 758 4328 762 4332
rect 806 4328 810 4332
rect 870 4328 874 4332
rect 1494 4338 1498 4342
rect 1510 4338 1514 4342
rect 1566 4338 1570 4342
rect 1710 4338 1714 4342
rect 1766 4338 1770 4342
rect 1798 4338 1802 4342
rect 1966 4338 1970 4342
rect 2078 4338 2082 4342
rect 2174 4338 2178 4342
rect 2214 4338 2218 4342
rect 2446 4338 2450 4342
rect 2646 4338 2650 4342
rect 2662 4338 2666 4342
rect 2686 4338 2690 4342
rect 2718 4338 2722 4342
rect 2950 4338 2954 4342
rect 3078 4338 3082 4342
rect 3238 4338 3242 4342
rect 3270 4338 3274 4342
rect 3366 4338 3370 4342
rect 3534 4338 3538 4342
rect 3630 4338 3634 4342
rect 3662 4338 3666 4342
rect 3678 4338 3682 4342
rect 3694 4338 3698 4342
rect 3726 4338 3730 4342
rect 3758 4338 3762 4342
rect 3774 4338 3778 4342
rect 3790 4338 3794 4342
rect 3822 4338 3826 4342
rect 3838 4338 3842 4342
rect 3878 4338 3882 4342
rect 3894 4338 3898 4342
rect 3918 4338 3922 4342
rect 3934 4338 3938 4342
rect 3966 4338 3970 4342
rect 3998 4338 4002 4342
rect 4054 4338 4058 4342
rect 4078 4338 4082 4342
rect 4126 4338 4130 4342
rect 4142 4338 4146 4342
rect 4182 4338 4186 4342
rect 4190 4338 4194 4342
rect 4238 4338 4242 4342
rect 4270 4338 4274 4342
rect 4334 4338 4338 4342
rect 4350 4338 4354 4342
rect 4390 4338 4394 4342
rect 4406 4338 4410 4342
rect 4422 4338 4426 4342
rect 4462 4338 4466 4342
rect 4518 4338 4522 4342
rect 4590 4338 4594 4342
rect 958 4328 962 4332
rect 1134 4328 1138 4332
rect 1166 4328 1170 4332
rect 1270 4328 1274 4332
rect 1318 4328 1322 4332
rect 1414 4328 1418 4332
rect 1582 4328 1586 4332
rect 1614 4328 1618 4332
rect 1726 4328 1730 4332
rect 1886 4328 1890 4332
rect 2126 4328 2130 4332
rect 2134 4328 2138 4332
rect 2198 4328 2202 4332
rect 2598 4328 2602 4332
rect 2710 4328 2714 4332
rect 2750 4327 2754 4331
rect 2774 4327 2778 4331
rect 2814 4328 2818 4332
rect 2886 4328 2890 4332
rect 2926 4328 2930 4332
rect 2974 4328 2978 4332
rect 2990 4328 2994 4332
rect 3302 4328 3306 4332
rect 3622 4328 3626 4332
rect 3806 4328 3810 4332
rect 3870 4328 3874 4332
rect 4094 4328 4098 4332
rect 4110 4328 4114 4332
rect 4230 4328 4234 4332
rect 4318 4328 4322 4332
rect 4486 4328 4490 4332
rect 4510 4328 4514 4332
rect 4534 4328 4538 4332
rect 254 4318 258 4322
rect 350 4318 354 4322
rect 374 4318 378 4322
rect 446 4318 450 4322
rect 606 4318 610 4322
rect 622 4318 626 4322
rect 678 4318 682 4322
rect 750 4318 754 4322
rect 926 4318 930 4322
rect 966 4318 970 4322
rect 990 4318 994 4322
rect 1102 4318 1106 4322
rect 1382 4318 1386 4322
rect 2182 4318 2186 4322
rect 2206 4318 2210 4322
rect 2246 4318 2250 4322
rect 2286 4318 2290 4322
rect 2326 4318 2330 4322
rect 2350 4318 2354 4322
rect 2406 4318 2410 4322
rect 2462 4318 2466 4322
rect 2518 4318 2522 4322
rect 2542 4318 2546 4322
rect 2614 4318 2618 4322
rect 2678 4318 2682 4322
rect 2702 4318 2706 4322
rect 2910 4318 2914 4322
rect 2934 4318 2938 4322
rect 2982 4318 2986 4322
rect 3006 4318 3010 4322
rect 3230 4318 3234 4322
rect 3638 4318 3642 4322
rect 3686 4318 3690 4322
rect 3886 4318 3890 4322
rect 4070 4318 4074 4322
rect 4134 4318 4138 4322
rect 4246 4318 4250 4322
rect 4438 4318 4442 4322
rect 4478 4318 4482 4322
rect 4526 4318 4530 4322
rect 1002 4303 1006 4307
rect 1009 4303 1013 4307
rect 2026 4303 2030 4307
rect 2033 4303 2037 4307
rect 3050 4303 3054 4307
rect 3057 4303 3061 4307
rect 4082 4303 4086 4307
rect 4089 4303 4093 4307
rect 334 4288 338 4292
rect 406 4288 410 4292
rect 686 4288 690 4292
rect 790 4288 794 4292
rect 934 4288 938 4292
rect 1286 4288 1290 4292
rect 1694 4288 1698 4292
rect 1718 4288 1722 4292
rect 1846 4288 1850 4292
rect 2078 4288 2082 4292
rect 2102 4288 2106 4292
rect 2254 4288 2258 4292
rect 2966 4288 2970 4292
rect 3142 4288 3146 4292
rect 3246 4288 3250 4292
rect 3446 4288 3450 4292
rect 3486 4288 3490 4292
rect 3518 4288 3522 4292
rect 3590 4288 3594 4292
rect 3622 4288 3626 4292
rect 3710 4288 3714 4292
rect 3990 4288 3994 4292
rect 4046 4288 4050 4292
rect 4118 4288 4122 4292
rect 4302 4288 4306 4292
rect 4366 4288 4370 4292
rect 6 4278 10 4282
rect 78 4278 82 4282
rect 358 4278 362 4282
rect 438 4278 442 4282
rect 462 4278 466 4282
rect 542 4278 546 4282
rect 638 4278 642 4282
rect 862 4278 866 4282
rect 1038 4278 1042 4282
rect 1254 4278 1258 4282
rect 1982 4278 1986 4282
rect 2022 4278 2026 4282
rect 2094 4278 2098 4282
rect 2230 4278 2234 4282
rect 2414 4278 2418 4282
rect 2438 4278 2442 4282
rect 2454 4278 2458 4282
rect 2502 4278 2506 4282
rect 2726 4278 2730 4282
rect 3006 4278 3010 4282
rect 3014 4278 3018 4282
rect 3094 4278 3098 4282
rect 3102 4278 3106 4282
rect 3134 4278 3138 4282
rect 3262 4278 3266 4282
rect 3334 4278 3338 4282
rect 3478 4278 3482 4282
rect 3614 4278 3618 4282
rect 3646 4278 3650 4282
rect 3702 4278 3706 4282
rect 3830 4278 3834 4282
rect 3982 4278 3986 4282
rect 4054 4278 4058 4282
rect 4062 4278 4066 4282
rect 4238 4278 4242 4282
rect 4422 4278 4426 4282
rect 22 4268 26 4272
rect 46 4268 50 4272
rect 62 4268 66 4272
rect 190 4268 194 4272
rect 302 4268 306 4272
rect 350 4268 354 4272
rect 382 4268 386 4272
rect 430 4268 434 4272
rect 574 4268 578 4272
rect 622 4268 626 4272
rect 646 4268 650 4272
rect 662 4268 666 4272
rect 670 4268 674 4272
rect 734 4268 738 4272
rect 806 4268 810 4272
rect 846 4268 850 4272
rect 886 4268 890 4272
rect 918 4268 922 4272
rect 974 4268 978 4272
rect 1046 4268 1050 4272
rect 1062 4268 1066 4272
rect 54 4258 58 4262
rect 70 4258 74 4262
rect 110 4259 114 4263
rect 142 4258 146 4262
rect 206 4259 210 4263
rect 302 4258 306 4262
rect 374 4258 378 4262
rect 454 4258 458 4262
rect 510 4258 514 4262
rect 542 4259 546 4263
rect 598 4258 602 4262
rect 630 4258 634 4262
rect 718 4259 722 4263
rect 822 4258 826 4262
rect 862 4258 866 4262
rect 878 4258 882 4262
rect 894 4258 898 4262
rect 910 4258 914 4262
rect 950 4258 954 4262
rect 982 4258 986 4262
rect 1038 4258 1042 4262
rect 1094 4268 1098 4272
rect 1110 4268 1114 4272
rect 1126 4268 1130 4272
rect 1158 4268 1162 4272
rect 1214 4268 1218 4272
rect 1230 4268 1234 4272
rect 1246 4268 1250 4272
rect 1270 4268 1274 4272
rect 1318 4268 1322 4272
rect 1342 4268 1346 4272
rect 1414 4268 1418 4272
rect 1478 4268 1482 4272
rect 1494 4268 1498 4272
rect 1510 4268 1514 4272
rect 1574 4268 1578 4272
rect 1590 4268 1594 4272
rect 1614 4268 1618 4272
rect 1702 4268 1706 4272
rect 1814 4268 1818 4272
rect 1950 4268 1954 4272
rect 1966 4268 1970 4272
rect 2038 4268 2042 4272
rect 2862 4268 2866 4272
rect 2982 4268 2986 4272
rect 3038 4268 3042 4272
rect 3054 4268 3058 4272
rect 3254 4268 3258 4272
rect 3366 4268 3370 4272
rect 3422 4268 3426 4272
rect 3430 4268 3434 4272
rect 3462 4268 3466 4272
rect 3502 4268 3506 4272
rect 3526 4268 3530 4272
rect 3534 4268 3538 4272
rect 3630 4268 3634 4272
rect 3662 4268 3666 4272
rect 3670 4268 3674 4272
rect 3734 4268 3738 4272
rect 3758 4268 3762 4272
rect 3790 4268 3794 4272
rect 3846 4268 3850 4272
rect 3870 4268 3874 4272
rect 3886 4268 3890 4272
rect 3902 4268 3906 4272
rect 3918 4268 3922 4272
rect 3974 4268 3978 4272
rect 3998 4268 4002 4272
rect 4038 4268 4042 4272
rect 4094 4268 4098 4272
rect 4126 4268 4130 4272
rect 4142 4268 4146 4272
rect 4166 4268 4170 4272
rect 1102 4258 1106 4262
rect 1118 4258 1122 4262
rect 1142 4258 1146 4262
rect 1166 4258 1170 4262
rect 1206 4258 1210 4262
rect 1222 4258 1226 4262
rect 1238 4258 1242 4262
rect 1278 4258 1282 4262
rect 1350 4259 1354 4263
rect 1406 4259 1410 4263
rect 1606 4259 1610 4263
rect 1678 4258 1682 4262
rect 1710 4258 1714 4262
rect 1750 4258 1754 4262
rect 1782 4259 1786 4263
rect 1822 4258 1826 4262
rect 1878 4258 1882 4262
rect 1910 4259 1914 4263
rect 2006 4258 2010 4262
rect 2134 4258 2138 4262
rect 2166 4259 2170 4263
rect 2214 4258 2218 4262
rect 2254 4258 2258 4262
rect 2286 4258 2290 4262
rect 2302 4258 2306 4262
rect 2326 4258 2330 4262
rect 2350 4258 2354 4262
rect 2374 4258 2378 4262
rect 2390 4258 2394 4262
rect 2438 4258 2442 4262
rect 2478 4258 2482 4262
rect 2526 4258 2530 4262
rect 2558 4258 2562 4262
rect 2574 4258 2578 4262
rect 2614 4258 2618 4262
rect 2638 4258 2642 4262
rect 2670 4258 2674 4262
rect 2686 4258 2690 4262
rect 2710 4258 2714 4262
rect 2750 4258 2754 4262
rect 2766 4258 2770 4262
rect 2790 4258 2794 4262
rect 2814 4258 2818 4262
rect 2830 4258 2834 4262
rect 2846 4258 2850 4262
rect 2886 4258 2890 4262
rect 2910 4258 2914 4262
rect 2950 4258 2954 4262
rect 2990 4258 2994 4262
rect 3174 4258 3178 4262
rect 3198 4258 3202 4262
rect 3286 4258 3290 4262
rect 3318 4258 3322 4262
rect 3358 4258 3362 4262
rect 3374 4258 3378 4262
rect 3414 4258 3418 4262
rect 3454 4258 3458 4262
rect 3542 4258 3546 4262
rect 3606 4258 3610 4262
rect 3638 4258 3642 4262
rect 3654 4258 3658 4262
rect 3670 4258 3674 4262
rect 3678 4258 3682 4262
rect 3694 4258 3698 4262
rect 3726 4258 3730 4262
rect 3766 4258 3770 4262
rect 3782 4258 3786 4262
rect 3814 4258 3818 4262
rect 3854 4258 3858 4262
rect 3862 4258 3866 4262
rect 3918 4258 3922 4262
rect 3958 4258 3962 4262
rect 3974 4258 3978 4262
rect 4006 4258 4010 4262
rect 4038 4258 4042 4262
rect 4086 4258 4090 4262
rect 4102 4258 4106 4262
rect 4118 4258 4122 4262
rect 4134 4258 4138 4262
rect 4198 4268 4202 4272
rect 4254 4268 4258 4272
rect 4270 4268 4274 4272
rect 4326 4268 4330 4272
rect 4358 4268 4362 4272
rect 4390 4268 4394 4272
rect 4406 4268 4410 4272
rect 4470 4268 4474 4272
rect 4486 4268 4490 4272
rect 4502 4268 4506 4272
rect 4518 4268 4522 4272
rect 4550 4268 4554 4272
rect 4558 4268 4562 4272
rect 4198 4258 4202 4262
rect 4230 4258 4234 4262
rect 4262 4258 4266 4262
rect 4278 4258 4282 4262
rect 4294 4258 4298 4262
rect 4318 4258 4322 4262
rect 4350 4258 4354 4262
rect 4390 4258 4394 4262
rect 4398 4258 4402 4262
rect 4430 4258 4434 4262
rect 4462 4258 4466 4262
rect 4478 4258 4482 4262
rect 4494 4258 4498 4262
rect 4542 4258 4546 4262
rect 4566 4258 4570 4262
rect 590 4248 594 4252
rect 686 4248 690 4252
rect 790 4248 794 4252
rect 814 4248 818 4252
rect 910 4248 914 4252
rect 934 4248 938 4252
rect 942 4248 946 4252
rect 998 4248 1002 4252
rect 1046 4248 1050 4252
rect 1062 4248 1066 4252
rect 1118 4248 1122 4252
rect 1150 4248 1154 4252
rect 1182 4248 1186 4252
rect 1838 4248 1842 4252
rect 1942 4248 1946 4252
rect 2022 4248 2026 4252
rect 2078 4248 2082 4252
rect 2230 4248 2234 4252
rect 2278 4248 2282 4252
rect 2342 4248 2346 4252
rect 2454 4248 2458 4252
rect 2590 4248 2594 4252
rect 2630 4248 2634 4252
rect 2662 4248 2666 4252
rect 2718 4248 2722 4252
rect 2798 4248 2802 4252
rect 2806 4248 2810 4252
rect 2838 4248 2842 4252
rect 2894 4248 2898 4252
rect 2958 4248 2962 4252
rect 2966 4248 2970 4252
rect 3038 4248 3042 4252
rect 3238 4248 3242 4252
rect 3302 4248 3306 4252
rect 3310 4248 3314 4252
rect 3342 4248 3346 4252
rect 3358 4248 3362 4252
rect 3382 4248 3386 4252
rect 3398 4248 3402 4252
rect 3446 4248 3450 4252
rect 3486 4248 3490 4252
rect 3510 4248 3514 4252
rect 3558 4248 3562 4252
rect 3710 4248 3714 4252
rect 3742 4248 3746 4252
rect 3798 4248 3802 4252
rect 3910 4248 3914 4252
rect 3942 4248 3946 4252
rect 4014 4248 4018 4252
rect 4158 4248 4162 4252
rect 4174 4248 4178 4252
rect 4206 4248 4210 4252
rect 4294 4248 4298 4252
rect 4334 4248 4338 4252
rect 4366 4248 4370 4252
rect 4454 4248 4458 4252
rect 4518 4248 4522 4252
rect 4582 4248 4586 4252
rect 254 4238 258 4242
rect 374 4238 378 4242
rect 814 4238 818 4242
rect 958 4238 962 4242
rect 1206 4238 1210 4242
rect 1254 4238 1258 4242
rect 1470 4238 1474 4242
rect 1998 4238 2002 4242
rect 2206 4238 2210 4242
rect 2262 4238 2266 4242
rect 2294 4238 2298 4242
rect 2318 4238 2322 4242
rect 2358 4238 2362 4242
rect 2382 4238 2386 4242
rect 2486 4238 2490 4242
rect 2534 4238 2538 4242
rect 2574 4238 2578 4242
rect 2606 4238 2610 4242
rect 2622 4238 2626 4242
rect 2678 4238 2682 4242
rect 2702 4238 2706 4242
rect 2742 4238 2746 4242
rect 2782 4238 2786 4242
rect 2790 4238 2794 4242
rect 2854 4238 2858 4242
rect 2878 4238 2882 4242
rect 2918 4238 2922 4242
rect 2942 4238 2946 4242
rect 3294 4238 3298 4242
rect 3326 4238 3330 4242
rect 4302 4238 4306 4242
rect 470 4228 474 4232
rect 2494 4228 2498 4232
rect 2950 4228 2954 4232
rect 3478 4228 3482 4232
rect 174 4218 178 4222
rect 270 4218 274 4222
rect 622 4218 626 4222
rect 782 4218 786 4222
rect 822 4218 826 4222
rect 854 4218 858 4222
rect 966 4218 970 4222
rect 1078 4218 1082 4222
rect 1822 4218 1826 4222
rect 2006 4218 2010 4222
rect 2086 4218 2090 4222
rect 2102 4218 2106 4222
rect 2214 4218 2218 4222
rect 2254 4218 2258 4222
rect 2326 4218 2330 4222
rect 2350 4218 2354 4222
rect 2582 4218 2586 4222
rect 2614 4218 2618 4222
rect 2654 4218 2658 4222
rect 2710 4218 2714 4222
rect 2790 4218 2794 4222
rect 2886 4218 2890 4222
rect 2926 4218 2930 4222
rect 2990 4218 2994 4222
rect 3118 4218 3122 4222
rect 3870 4218 3874 4222
rect 498 4203 502 4207
rect 505 4203 509 4207
rect 1522 4203 1526 4207
rect 1529 4203 1533 4207
rect 2546 4203 2550 4207
rect 2553 4203 2557 4207
rect 3570 4203 3574 4207
rect 3577 4203 3581 4207
rect 30 4188 34 4192
rect 446 4188 450 4192
rect 478 4188 482 4192
rect 630 4188 634 4192
rect 942 4188 946 4192
rect 1094 4188 1098 4192
rect 1662 4188 1666 4192
rect 1790 4188 1794 4192
rect 1822 4188 1826 4192
rect 1974 4188 1978 4192
rect 2030 4188 2034 4192
rect 2134 4188 2138 4192
rect 2334 4188 2338 4192
rect 2590 4188 2594 4192
rect 2662 4188 2666 4192
rect 2782 4188 2786 4192
rect 2918 4188 2922 4192
rect 2934 4188 2938 4192
rect 3246 4188 3250 4192
rect 3278 4188 3282 4192
rect 3374 4188 3378 4192
rect 3470 4188 3474 4192
rect 3502 4188 3506 4192
rect 3510 4188 3514 4192
rect 3894 4188 3898 4192
rect 3926 4188 3930 4192
rect 4014 4188 4018 4192
rect 4078 4188 4082 4192
rect 4550 4188 4554 4192
rect 694 4178 698 4182
rect 2246 4178 2250 4182
rect 2390 4178 2394 4182
rect 558 4168 562 4172
rect 870 4168 874 4172
rect 878 4168 882 4172
rect 1142 4168 1146 4172
rect 1286 4168 1290 4172
rect 1334 4168 1338 4172
rect 1806 4168 1810 4172
rect 1838 4168 1842 4172
rect 1902 4168 1906 4172
rect 1926 4168 1930 4172
rect 2014 4168 2018 4172
rect 2054 4168 2058 4172
rect 2174 4168 2178 4172
rect 2326 4168 2330 4172
rect 2446 4168 2450 4172
rect 2478 4168 2482 4172
rect 2502 4168 2506 4172
rect 2686 4168 2690 4172
rect 2942 4168 2946 4172
rect 2974 4168 2978 4172
rect 2998 4168 3002 4172
rect 3238 4168 3242 4172
rect 3270 4168 3274 4172
rect 3302 4168 3306 4172
rect 3310 4168 3314 4172
rect 3350 4168 3354 4172
rect 3966 4168 3970 4172
rect 118 4158 122 4162
rect 254 4158 258 4162
rect 574 4158 578 4162
rect 598 4158 602 4162
rect 798 4158 802 4162
rect 814 4158 818 4162
rect 854 4158 858 4162
rect 894 4158 898 4162
rect 1078 4158 1082 4162
rect 1262 4158 1266 4162
rect 1446 4158 1450 4162
rect 1494 4158 1498 4162
rect 1710 4158 1714 4162
rect 1742 4158 1746 4162
rect 54 4148 58 4152
rect 174 4148 178 4152
rect 214 4148 218 4152
rect 230 4148 234 4152
rect 262 4148 266 4152
rect 286 4148 290 4152
rect 318 4148 322 4152
rect 350 4148 354 4152
rect 382 4147 386 4151
rect 726 4148 730 4152
rect 742 4148 746 4152
rect 806 4148 810 4152
rect 878 4148 882 4152
rect 1942 4158 1946 4162
rect 2110 4158 2114 4162
rect 2206 4158 2210 4162
rect 2222 4158 2226 4162
rect 2278 4158 2282 4162
rect 2398 4158 2402 4162
rect 2422 4158 2426 4162
rect 2430 4158 2434 4162
rect 2462 4158 2466 4162
rect 2518 4158 2522 4162
rect 2526 4158 2530 4162
rect 2614 4158 2618 4162
rect 2926 4158 2930 4162
rect 3142 4157 3146 4161
rect 3254 4158 3258 4162
rect 3286 4158 3290 4162
rect 3318 4158 3322 4162
rect 3358 4158 3362 4162
rect 3454 4158 3458 4162
rect 3766 4158 3770 4162
rect 3798 4158 3802 4162
rect 3910 4158 3914 4162
rect 3950 4158 3954 4162
rect 3974 4158 3978 4162
rect 4134 4158 4138 4162
rect 4150 4158 4154 4162
rect 4198 4158 4202 4162
rect 926 4148 930 4152
rect 942 4148 946 4152
rect 974 4148 978 4152
rect 1006 4148 1010 4152
rect 1118 4148 1122 4152
rect 1134 4148 1138 4152
rect 22 4138 26 4142
rect 62 4138 66 4142
rect 86 4138 90 4142
rect 134 4138 138 4142
rect 182 4138 186 4142
rect 206 4138 210 4142
rect 238 4138 242 4142
rect 254 4138 258 4142
rect 294 4138 298 4142
rect 326 4138 330 4142
rect 342 4138 346 4142
rect 366 4138 370 4142
rect 454 4138 458 4142
rect 534 4138 538 4142
rect 558 4138 562 4142
rect 598 4138 602 4142
rect 606 4138 610 4142
rect 638 4138 642 4142
rect 678 4138 682 4142
rect 686 4138 690 4142
rect 702 4138 706 4142
rect 718 4138 722 4142
rect 734 4138 738 4142
rect 774 4138 778 4142
rect 798 4138 802 4142
rect 830 4138 834 4142
rect 838 4138 842 4142
rect 854 4138 858 4142
rect 1206 4147 1210 4151
rect 1238 4148 1242 4152
rect 1278 4148 1282 4152
rect 1318 4148 1322 4152
rect 1398 4147 1402 4151
rect 1622 4147 1626 4151
rect 1678 4148 1682 4152
rect 1694 4148 1698 4152
rect 1710 4148 1714 4152
rect 1726 4148 1730 4152
rect 1750 4148 1754 4152
rect 1774 4148 1778 4152
rect 1822 4148 1826 4152
rect 1846 4148 1850 4152
rect 1886 4148 1890 4152
rect 1894 4148 1898 4152
rect 1910 4148 1914 4152
rect 2006 4148 2010 4152
rect 2062 4148 2066 4152
rect 2094 4148 2098 4152
rect 2166 4148 2170 4152
rect 2222 4148 2226 4152
rect 2334 4148 2338 4152
rect 2438 4148 2442 4152
rect 2470 4148 2474 4152
rect 2486 4148 2490 4152
rect 2510 4148 2514 4152
rect 2678 4148 2682 4152
rect 918 4138 922 4142
rect 1046 4138 1050 4142
rect 1062 4138 1066 4142
rect 1110 4138 1114 4142
rect 1126 4138 1130 4142
rect 1222 4138 1226 4142
rect 1246 4138 1250 4142
rect 1262 4138 1266 4142
rect 1270 4138 1274 4142
rect 1302 4138 1306 4142
rect 1414 4138 1418 4142
rect 1438 4138 1442 4142
rect 1470 4138 1474 4142
rect 1518 4138 1522 4142
rect 1614 4138 1618 4142
rect 1686 4138 1690 4142
rect 2750 4147 2754 4151
rect 2798 4148 2802 4152
rect 2830 4148 2834 4152
rect 2846 4148 2850 4152
rect 2862 4148 2866 4152
rect 2894 4148 2898 4152
rect 2966 4148 2970 4152
rect 2974 4148 2978 4152
rect 3038 4148 3042 4152
rect 3126 4148 3130 4152
rect 3158 4148 3162 4152
rect 3246 4148 3250 4152
rect 3278 4148 3282 4152
rect 3310 4148 3314 4152
rect 3334 4148 3338 4152
rect 3374 4148 3378 4152
rect 3446 4148 3450 4152
rect 3486 4148 3490 4152
rect 3502 4148 3506 4152
rect 3566 4148 3570 4152
rect 3582 4148 3586 4152
rect 3678 4148 3682 4152
rect 3782 4148 3786 4152
rect 3814 4148 3818 4152
rect 3830 4148 3834 4152
rect 3894 4148 3898 4152
rect 3950 4148 3954 4152
rect 3990 4148 3994 4152
rect 4038 4148 4042 4152
rect 4054 4148 4058 4152
rect 4062 4148 4066 4152
rect 4110 4148 4114 4152
rect 4150 4148 4154 4152
rect 4174 4148 4178 4152
rect 4238 4158 4242 4162
rect 4254 4158 4258 4162
rect 4270 4158 4274 4162
rect 4286 4158 4290 4162
rect 4358 4158 4362 4162
rect 4390 4158 4394 4162
rect 4438 4158 4442 4162
rect 4446 4158 4450 4162
rect 4518 4158 4522 4162
rect 4222 4148 4226 4152
rect 4254 4148 4258 4152
rect 4294 4148 4298 4152
rect 4302 4148 4306 4152
rect 4334 4148 4338 4152
rect 4366 4148 4370 4152
rect 4430 4148 4434 4152
rect 4454 4148 4458 4152
rect 4462 4148 4466 4152
rect 4486 4148 4490 4152
rect 4502 4148 4506 4152
rect 4518 4148 4522 4152
rect 4534 4148 4538 4152
rect 4566 4148 4570 4152
rect 4582 4148 4586 4152
rect 4598 4148 4602 4152
rect 1718 4138 1722 4142
rect 1750 4138 1754 4142
rect 1782 4138 1786 4142
rect 1814 4138 1818 4142
rect 1862 4138 1866 4142
rect 1870 4138 1874 4142
rect 1958 4138 1962 4142
rect 2206 4138 2210 4142
rect 2398 4138 2402 4142
rect 2766 4138 2770 4142
rect 2806 4138 2810 4142
rect 2838 4138 2842 4142
rect 2870 4138 2874 4142
rect 2878 4138 2882 4142
rect 2894 4138 2898 4142
rect 2942 4138 2946 4142
rect 3078 4138 3082 4142
rect 3094 4138 3098 4142
rect 3102 4138 3106 4142
rect 3166 4138 3170 4142
rect 3222 4138 3226 4142
rect 3310 4138 3314 4142
rect 3390 4138 3394 4142
rect 3430 4138 3434 4142
rect 3478 4138 3482 4142
rect 3574 4138 3578 4142
rect 3726 4138 3730 4142
rect 3774 4138 3778 4142
rect 3822 4138 3826 4142
rect 3934 4138 3938 4142
rect 4006 4138 4010 4142
rect 4118 4138 4122 4142
rect 4134 4138 4138 4142
rect 4174 4138 4178 4142
rect 4182 4138 4186 4142
rect 4206 4138 4210 4142
rect 4230 4138 4234 4142
rect 4262 4138 4266 4142
rect 4294 4138 4298 4142
rect 4310 4138 4314 4142
rect 4366 4138 4370 4142
rect 4406 4138 4410 4142
rect 4414 4138 4418 4142
rect 4438 4138 4442 4142
rect 4478 4138 4482 4142
rect 4510 4138 4514 4142
rect 4542 4138 4546 4142
rect 4574 4138 4578 4142
rect 4590 4138 4594 4142
rect 6 4128 10 4132
rect 78 4128 82 4132
rect 190 4128 194 4132
rect 214 4128 218 4132
rect 254 4128 258 4132
rect 310 4128 314 4132
rect 486 4128 490 4132
rect 646 4128 650 4132
rect 766 4128 770 4132
rect 958 4128 962 4132
rect 1030 4128 1034 4132
rect 1038 4128 1042 4132
rect 1086 4128 1090 4132
rect 1318 4128 1322 4132
rect 1430 4128 1434 4132
rect 1486 4128 1490 4132
rect 1966 4128 1970 4132
rect 1982 4128 1986 4132
rect 2086 4128 2090 4132
rect 2126 4128 2130 4132
rect 2142 4128 2146 4132
rect 2190 4128 2194 4132
rect 2262 4128 2266 4132
rect 2310 4128 2314 4132
rect 2358 4128 2362 4132
rect 2366 4128 2370 4132
rect 2574 4128 2578 4132
rect 2582 4128 2586 4132
rect 2598 4128 2602 4132
rect 2646 4128 2650 4132
rect 2878 4128 2882 4132
rect 3086 4128 3090 4132
rect 3190 4128 3194 4132
rect 3222 4128 3226 4132
rect 3430 4128 3434 4132
rect 3486 4128 3490 4132
rect 3526 4128 3530 4132
rect 3590 4128 3594 4132
rect 3638 4128 3642 4132
rect 3678 4128 3682 4132
rect 3718 4128 3722 4132
rect 3814 4128 3818 4132
rect 3870 4128 3874 4132
rect 4038 4128 4042 4132
rect 4326 4128 4330 4132
rect 4486 4128 4490 4132
rect 4558 4128 4562 4132
rect 182 4118 186 4122
rect 286 4118 290 4122
rect 302 4118 306 4122
rect 334 4118 338 4122
rect 526 4118 530 4122
rect 574 4118 578 4122
rect 614 4118 618 4122
rect 670 4118 674 4122
rect 710 4118 714 4122
rect 822 4118 826 4122
rect 1326 4118 1330 4122
rect 1662 4118 1666 4122
rect 1742 4118 1746 4122
rect 1950 4118 1954 4122
rect 2062 4118 2066 4122
rect 2182 4118 2186 4122
rect 2222 4118 2226 4122
rect 2270 4118 2274 4122
rect 2278 4118 2282 4122
rect 2422 4118 2426 4122
rect 2454 4118 2458 4122
rect 2510 4118 2514 4122
rect 2526 4118 2530 4122
rect 2606 4118 2610 4122
rect 2614 4118 2618 4122
rect 2814 4118 2818 4122
rect 3430 4118 3434 4122
rect 3574 4118 3578 4122
rect 3630 4118 3634 4122
rect 3686 4118 3690 4122
rect 3846 4118 3850 4122
rect 3926 4118 3930 4122
rect 4046 4118 4050 4122
rect 1002 4103 1006 4107
rect 1009 4103 1013 4107
rect 2026 4103 2030 4107
rect 2033 4103 2037 4107
rect 3050 4103 3054 4107
rect 3057 4103 3061 4107
rect 4082 4103 4086 4107
rect 4089 4103 4093 4107
rect 110 4088 114 4092
rect 590 4088 594 4092
rect 966 4088 970 4092
rect 1038 4088 1042 4092
rect 1190 4088 1194 4092
rect 1286 4088 1290 4092
rect 1550 4088 1554 4092
rect 1646 4088 1650 4092
rect 1742 4088 1746 4092
rect 2302 4088 2306 4092
rect 2686 4088 2690 4092
rect 2942 4088 2946 4092
rect 3078 4088 3082 4092
rect 3246 4088 3250 4092
rect 3310 4088 3314 4092
rect 3350 4088 3354 4092
rect 3398 4088 3402 4092
rect 3454 4088 3458 4092
rect 3518 4088 3522 4092
rect 3558 4088 3562 4092
rect 3678 4088 3682 4092
rect 3766 4088 3770 4092
rect 4206 4088 4210 4092
rect 4318 4088 4322 4092
rect 4446 4088 4450 4092
rect 174 4078 178 4082
rect 310 4078 314 4082
rect 718 4078 722 4082
rect 734 4078 738 4082
rect 774 4078 778 4082
rect 902 4078 906 4082
rect 974 4078 978 4082
rect 982 4078 986 4082
rect 990 4078 994 4082
rect 1006 4078 1010 4082
rect 1022 4078 1026 4082
rect 1222 4078 1226 4082
rect 1614 4078 1618 4082
rect 1774 4078 1778 4082
rect 1990 4078 1994 4082
rect 2054 4078 2058 4082
rect 2246 4078 2250 4082
rect 2334 4078 2338 4082
rect 2382 4078 2386 4082
rect 2446 4078 2450 4082
rect 2470 4078 2474 4082
rect 2558 4078 2562 4082
rect 2638 4078 2642 4082
rect 2654 4078 2658 4082
rect 3070 4078 3074 4082
rect 3174 4078 3178 4082
rect 3198 4078 3202 4082
rect 3238 4078 3242 4082
rect 3278 4078 3282 4082
rect 3358 4078 3362 4082
rect 3366 4078 3370 4082
rect 3454 4078 3458 4082
rect 3518 4078 3522 4082
rect 3646 4078 3650 4082
rect 3686 4078 3690 4082
rect 4054 4078 4058 4082
rect 4166 4078 4170 4082
rect 4190 4078 4194 4082
rect 4198 4078 4202 4082
rect 4518 4078 4522 4082
rect 4526 4078 4530 4082
rect 30 4068 34 4072
rect 166 4068 170 4072
rect 174 4068 178 4072
rect 190 4068 194 4072
rect 222 4068 226 4072
rect 230 4068 234 4072
rect 254 4068 258 4072
rect 270 4068 274 4072
rect 302 4068 306 4072
rect 350 4068 354 4072
rect 446 4068 450 4072
rect 510 4068 514 4072
rect 654 4068 658 4072
rect 726 4068 730 4072
rect 750 4068 754 4072
rect 798 4068 802 4072
rect 822 4068 826 4072
rect 830 4068 834 4072
rect 886 4068 890 4072
rect 910 4068 914 4072
rect 958 4068 962 4072
rect 1030 4068 1034 4072
rect 1062 4068 1066 4072
rect 1094 4068 1098 4072
rect 1230 4068 1234 4072
rect 1390 4068 1394 4072
rect 1414 4068 1418 4072
rect 1462 4068 1466 4072
rect 1494 4068 1498 4072
rect 1518 4068 1522 4072
rect 1766 4068 1770 4072
rect 1790 4068 1794 4072
rect 1814 4068 1818 4072
rect 1846 4068 1850 4072
rect 1854 4068 1858 4072
rect 1886 4068 1890 4072
rect 2598 4068 2602 4072
rect 2654 4068 2658 4072
rect 2734 4068 2738 4072
rect 2758 4068 2762 4072
rect 2774 4068 2778 4072
rect 2998 4068 3002 4072
rect 3174 4068 3178 4072
rect 3318 4068 3322 4072
rect 3326 4068 3330 4072
rect 3406 4068 3410 4072
rect 3454 4068 3458 4072
rect 3550 4068 3554 4072
rect 3598 4068 3602 4072
rect 3654 4068 3658 4072
rect 3742 4068 3746 4072
rect 3774 4068 3778 4072
rect 3806 4068 3810 4072
rect 3862 4068 3866 4072
rect 3870 4068 3874 4072
rect 3894 4068 3898 4072
rect 3990 4068 3994 4072
rect 4054 4068 4058 4072
rect 4078 4068 4082 4072
rect 4086 4068 4090 4072
rect 4134 4068 4138 4072
rect 4142 4068 4146 4072
rect 4174 4068 4178 4072
rect 4214 4068 4218 4072
rect 4230 4068 4234 4072
rect 4262 4068 4266 4072
rect 4294 4068 4298 4072
rect 4326 4068 4330 4072
rect 4358 4068 4362 4072
rect 4390 4068 4394 4072
rect 4422 4068 4426 4072
rect 4478 4068 4482 4072
rect 4510 4068 4514 4072
rect 4542 4068 4546 4072
rect 4558 4068 4562 4072
rect 4574 4068 4578 4072
rect 38 4058 42 4062
rect 198 4058 202 4062
rect 214 4058 218 4062
rect 230 4058 234 4062
rect 246 4058 250 4062
rect 270 4058 274 4062
rect 310 4058 314 4062
rect 326 4058 330 4062
rect 342 4058 346 4062
rect 358 4058 362 4062
rect 374 4058 378 4062
rect 470 4058 474 4062
rect 526 4059 530 4063
rect 614 4058 618 4062
rect 630 4058 634 4062
rect 686 4058 690 4062
rect 758 4058 762 4062
rect 782 4058 786 4062
rect 806 4058 810 4062
rect 862 4058 866 4062
rect 886 4058 890 4062
rect 918 4058 922 4062
rect 934 4058 938 4062
rect 950 4058 954 4062
rect 990 4058 994 4062
rect 1046 4058 1050 4062
rect 1086 4058 1090 4062
rect 1126 4059 1130 4063
rect 1158 4058 1162 4062
rect 1222 4059 1226 4063
rect 1310 4058 1314 4062
rect 1398 4058 1402 4062
rect 1422 4058 1426 4062
rect 1462 4058 1466 4062
rect 1494 4058 1498 4062
rect 1542 4058 1546 4062
rect 1582 4058 1586 4062
rect 1614 4059 1618 4063
rect 1678 4058 1682 4062
rect 1710 4059 1714 4063
rect 1758 4058 1762 4062
rect 1838 4058 1842 4062
rect 1878 4058 1882 4062
rect 1910 4058 1914 4062
rect 1918 4058 1922 4062
rect 1966 4058 1970 4062
rect 2014 4058 2018 4062
rect 2062 4058 2066 4062
rect 2110 4058 2114 4062
rect 2190 4058 2194 4062
rect 2262 4058 2266 4062
rect 2286 4058 2290 4062
rect 2334 4058 2338 4062
rect 2358 4058 2362 4062
rect 2406 4058 2410 4062
rect 2446 4058 2450 4062
rect 2494 4058 2498 4062
rect 2534 4058 2538 4062
rect 2582 4058 2586 4062
rect 2622 4058 2626 4062
rect 2670 4058 2674 4062
rect 2710 4058 2714 4062
rect 2798 4058 2802 4062
rect 2830 4058 2834 4062
rect 2846 4058 2850 4062
rect 2894 4058 2898 4062
rect 2910 4058 2914 4062
rect 2926 4058 2930 4062
rect 2998 4058 3002 4062
rect 3038 4058 3042 4062
rect 3134 4058 3138 4062
rect 3190 4058 3194 4062
rect 3198 4058 3202 4062
rect 3222 4058 3226 4062
rect 3262 4058 3266 4062
rect 3302 4058 3306 4062
rect 3342 4058 3346 4062
rect 3382 4058 3386 4062
rect 3446 4058 3450 4062
rect 3510 4058 3514 4062
rect 3558 4058 3562 4062
rect 3590 4058 3594 4062
rect 3622 4058 3626 4062
rect 3662 4058 3666 4062
rect 3702 4058 3706 4062
rect 3726 4058 3730 4062
rect 3750 4058 3754 4062
rect 3782 4058 3786 4062
rect 3806 4058 3810 4062
rect 3814 4058 3818 4062
rect 3830 4058 3834 4062
rect 3854 4058 3858 4062
rect 3878 4058 3882 4062
rect 3918 4058 3922 4062
rect 3926 4058 3930 4062
rect 3950 4058 3954 4062
rect 3966 4058 3970 4062
rect 3982 4058 3986 4062
rect 4030 4058 4034 4062
rect 4070 4058 4074 4062
rect 4094 4058 4098 4062
rect 4126 4058 4130 4062
rect 4150 4058 4154 4062
rect 4166 4058 4170 4062
rect 4182 4058 4186 4062
rect 4222 4058 4226 4062
rect 4238 4058 4242 4062
rect 4262 4058 4266 4062
rect 4270 4058 4274 4062
rect 4302 4058 4306 4062
rect 4326 4058 4330 4062
rect 4390 4058 4394 4062
rect 4398 4058 4402 4062
rect 4422 4058 4426 4062
rect 4430 4058 4434 4062
rect 4470 4058 4474 4062
rect 4502 4058 4506 4062
rect 4534 4058 4538 4062
rect 4566 4058 4570 4062
rect 4582 4058 4586 4062
rect 366 4048 370 4052
rect 486 4048 490 4052
rect 598 4048 602 4052
rect 670 4048 674 4052
rect 710 4048 714 4052
rect 774 4048 778 4052
rect 798 4048 802 4052
rect 846 4048 850 4052
rect 894 4048 898 4052
rect 934 4048 938 4052
rect 1070 4048 1074 4052
rect 1318 4048 1322 4052
rect 1486 4048 1490 4052
rect 1502 4048 1506 4052
rect 1742 4048 1746 4052
rect 2078 4048 2082 4052
rect 2118 4048 2122 4052
rect 2126 4048 2130 4052
rect 2182 4048 2186 4052
rect 2214 4048 2218 4052
rect 2254 4048 2258 4052
rect 2334 4048 2338 4052
rect 2350 4048 2354 4052
rect 2422 4048 2426 4052
rect 2502 4048 2506 4052
rect 2630 4048 2634 4052
rect 2702 4048 2706 4052
rect 2750 4048 2754 4052
rect 2774 4048 2778 4052
rect 2806 4048 2810 4052
rect 2838 4048 2842 4052
rect 2902 4048 2906 4052
rect 3198 4048 3202 4052
rect 3214 4048 3218 4052
rect 3574 4048 3578 4052
rect 3606 4048 3610 4052
rect 3734 4048 3738 4052
rect 3766 4048 3770 4052
rect 3798 4048 3802 4052
rect 3830 4048 3834 4052
rect 3838 4048 3842 4052
rect 3894 4048 3898 4052
rect 3934 4048 3938 4052
rect 3958 4048 3962 4052
rect 3966 4048 3970 4052
rect 4022 4048 4026 4052
rect 4110 4048 4114 4052
rect 4254 4048 4258 4052
rect 4270 4048 4274 4052
rect 4414 4048 4418 4052
rect 4446 4048 4450 4052
rect 4454 4048 4458 4052
rect 4486 4048 4490 4052
rect 4598 4048 4602 4052
rect 374 4038 378 4042
rect 430 4038 434 4042
rect 462 4038 466 4042
rect 606 4038 610 4042
rect 678 4038 682 4042
rect 830 4038 834 4042
rect 854 4038 858 4042
rect 1174 4038 1178 4042
rect 1302 4038 1306 4042
rect 1822 4038 1826 4042
rect 1934 4038 1938 4042
rect 1958 4038 1962 4042
rect 2006 4038 2010 4042
rect 2102 4038 2106 4042
rect 2142 4038 2146 4042
rect 2198 4038 2202 4042
rect 2230 4038 2234 4042
rect 2270 4038 2274 4042
rect 2326 4038 2330 4042
rect 2366 4038 2370 4042
rect 2414 4038 2418 4042
rect 2438 4038 2442 4042
rect 2486 4038 2490 4042
rect 2518 4038 2522 4042
rect 2590 4038 2594 4042
rect 2614 4038 2618 4042
rect 2718 4038 2722 4042
rect 2734 4038 2738 4042
rect 2790 4038 2794 4042
rect 2822 4038 2826 4042
rect 2910 4038 2914 4042
rect 2926 4038 2930 4042
rect 2958 4038 2962 4042
rect 3046 4038 3050 4042
rect 3094 4038 3098 4042
rect 3230 4038 3234 4042
rect 3718 4038 3722 4042
rect 3910 4038 3914 4042
rect 3942 4038 3946 4042
rect 4286 4038 4290 4042
rect 4318 4038 4322 4042
rect 4350 4038 4354 4042
rect 4470 4038 4474 4042
rect 4542 4038 4546 4042
rect 1310 4028 1314 4032
rect 94 4018 98 4022
rect 214 4018 218 4022
rect 294 4018 298 4022
rect 390 4018 394 4022
rect 470 4018 474 4022
rect 622 4018 626 4022
rect 702 4018 706 4022
rect 734 4018 738 4022
rect 1038 4018 1042 4022
rect 1334 4018 1338 4022
rect 1966 4018 1970 4022
rect 2014 4018 2018 4022
rect 2110 4018 2114 4022
rect 2174 4018 2178 4022
rect 2190 4018 2194 4022
rect 2278 4018 2282 4022
rect 2374 4018 2378 4022
rect 2494 4018 2498 4022
rect 2622 4018 2626 4022
rect 2646 4018 2650 4022
rect 2726 4018 2730 4022
rect 2798 4018 2802 4022
rect 2830 4018 2834 4022
rect 2862 4018 2866 4022
rect 2894 4018 2898 4022
rect 2934 4018 2938 4022
rect 3334 4018 3338 4022
rect 3622 4018 3626 4022
rect 3726 4018 3730 4022
rect 3854 4018 3858 4022
rect 3918 4018 3922 4022
rect 4334 4018 4338 4022
rect 498 4003 502 4007
rect 505 4003 509 4007
rect 1522 4003 1526 4007
rect 1529 4003 1533 4007
rect 2546 4003 2550 4007
rect 2553 4003 2557 4007
rect 3570 4003 3574 4007
rect 3577 4003 3581 4007
rect 70 3988 74 3992
rect 238 3988 242 3992
rect 286 3988 290 3992
rect 398 3988 402 3992
rect 502 3988 506 3992
rect 566 3988 570 3992
rect 694 3988 698 3992
rect 886 3988 890 3992
rect 1006 3988 1010 3992
rect 1214 3988 1218 3992
rect 1430 3988 1434 3992
rect 1494 3988 1498 3992
rect 1646 3988 1650 3992
rect 1758 3988 1762 3992
rect 1782 3988 1786 3992
rect 1814 3988 1818 3992
rect 1870 3988 1874 3992
rect 2334 3988 2338 3992
rect 2470 3988 2474 3992
rect 2750 3988 2754 3992
rect 2990 3988 2994 3992
rect 3030 3988 3034 3992
rect 3174 3988 3178 3992
rect 3270 3988 3274 3992
rect 3342 3988 3346 3992
rect 3382 3988 3386 3992
rect 3438 3988 3442 3992
rect 3494 3988 3498 3992
rect 3766 3988 3770 3992
rect 4150 3988 4154 3992
rect 4326 3988 4330 3992
rect 4518 3988 4522 3992
rect 2622 3978 2626 3982
rect 3414 3978 3418 3982
rect 350 3968 354 3972
rect 734 3968 738 3972
rect 1230 3968 1234 3972
rect 1974 3968 1978 3972
rect 2342 3968 2346 3972
rect 2614 3968 2618 3972
rect 2710 3968 2714 3972
rect 2830 3968 2834 3972
rect 3334 3968 3338 3972
rect 3390 3968 3394 3972
rect 3446 3968 3450 3972
rect 4542 3968 4546 3972
rect 4582 3968 4586 3972
rect 326 3958 330 3962
rect 430 3958 434 3962
rect 814 3958 818 3962
rect 830 3958 834 3962
rect 854 3958 858 3962
rect 1406 3958 1410 3962
rect 1526 3958 1530 3962
rect 1766 3958 1770 3962
rect 1798 3958 1802 3962
rect 1926 3958 1930 3962
rect 1990 3958 1994 3962
rect 2094 3958 2098 3962
rect 2126 3958 2130 3962
rect 2150 3958 2154 3962
rect 2206 3958 2210 3962
rect 2246 3958 2250 3962
rect 2318 3958 2322 3962
rect 2598 3958 2602 3962
rect 2630 3958 2634 3962
rect 2670 3958 2674 3962
rect 2694 3958 2698 3962
rect 2742 3958 2746 3962
rect 2798 3958 2802 3962
rect 2862 3958 2866 3962
rect 2894 3958 2898 3962
rect 3142 3958 3146 3962
rect 3254 3958 3258 3962
rect 3350 3958 3354 3962
rect 3382 3958 3386 3962
rect 3422 3958 3426 3962
rect 3430 3958 3434 3962
rect 3550 3958 3554 3962
rect 3566 3958 3570 3962
rect 3582 3958 3586 3962
rect 3646 3958 3650 3962
rect 3710 3958 3714 3962
rect 3982 3958 3986 3962
rect 4022 3958 4026 3962
rect 4086 3958 4090 3962
rect 4334 3958 4338 3962
rect 4430 3958 4434 3962
rect 4478 3958 4482 3962
rect 46 3948 50 3952
rect 126 3948 130 3952
rect 222 3948 226 3952
rect 254 3948 258 3952
rect 270 3948 274 3952
rect 302 3948 306 3952
rect 334 3948 338 3952
rect 358 3948 362 3952
rect 446 3948 450 3952
rect 462 3948 466 3952
rect 478 3948 482 3952
rect 510 3948 514 3952
rect 630 3947 634 3951
rect 742 3948 746 3952
rect 926 3947 930 3951
rect 958 3948 962 3952
rect 1038 3948 1042 3952
rect 1046 3948 1050 3952
rect 1150 3948 1154 3952
rect 1182 3947 1186 3951
rect 1270 3948 1274 3952
rect 1342 3948 1346 3952
rect 1374 3947 1378 3951
rect 1582 3948 1586 3952
rect 1606 3947 1610 3951
rect 1662 3948 1666 3952
rect 1694 3947 1698 3951
rect 1782 3948 1786 3952
rect 1814 3948 1818 3952
rect 1886 3948 1890 3952
rect 1894 3948 1898 3952
rect 1918 3948 1922 3952
rect 1982 3948 1986 3952
rect 1998 3948 2002 3952
rect 2046 3948 2050 3952
rect 2182 3948 2186 3952
rect 2214 3948 2218 3952
rect 2358 3948 2362 3952
rect 2390 3948 2394 3952
rect 2422 3948 2426 3952
rect 2454 3948 2458 3952
rect 2518 3948 2522 3952
rect 2558 3948 2562 3952
rect 2606 3948 2610 3952
rect 2702 3948 2706 3952
rect 2734 3948 2738 3952
rect 206 3938 210 3942
rect 230 3938 234 3942
rect 262 3938 266 3942
rect 278 3938 282 3942
rect 302 3938 306 3942
rect 310 3938 314 3942
rect 326 3938 330 3942
rect 374 3938 378 3942
rect 382 3938 386 3942
rect 406 3938 410 3942
rect 414 3938 418 3942
rect 470 3938 474 3942
rect 486 3938 490 3942
rect 550 3938 554 3942
rect 598 3938 602 3942
rect 614 3938 618 3942
rect 758 3938 762 3942
rect 814 3938 818 3942
rect 838 3938 842 3942
rect 862 3938 866 3942
rect 894 3938 898 3942
rect 1110 3938 1114 3942
rect 1294 3938 1298 3942
rect 1486 3938 1490 3942
rect 1678 3938 1682 3942
rect 1790 3938 1794 3942
rect 1822 3938 1826 3942
rect 1838 3938 1842 3942
rect 1862 3938 1866 3942
rect 2926 3947 2930 3951
rect 2958 3948 2962 3952
rect 3022 3948 3026 3952
rect 3094 3948 3098 3952
rect 3262 3948 3266 3952
rect 3294 3948 3298 3952
rect 3342 3948 3346 3952
rect 3374 3948 3378 3952
rect 3438 3948 3442 3952
rect 3470 3948 3474 3952
rect 3478 3948 3482 3952
rect 3510 3948 3514 3952
rect 3526 3948 3530 3952
rect 3542 3948 3546 3952
rect 3590 3948 3594 3952
rect 3606 3948 3610 3952
rect 3630 3948 3634 3952
rect 3726 3948 3730 3952
rect 3782 3948 3786 3952
rect 3798 3948 3802 3952
rect 3814 3948 3818 3952
rect 3830 3948 3834 3952
rect 3854 3948 3858 3952
rect 3870 3948 3874 3952
rect 3886 3948 3890 3952
rect 3918 3948 3922 3952
rect 3926 3948 3930 3952
rect 3966 3948 3970 3952
rect 4006 3948 4010 3952
rect 4062 3948 4066 3952
rect 4102 3948 4106 3952
rect 4134 3948 4138 3952
rect 4166 3948 4170 3952
rect 4198 3948 4202 3952
rect 4206 3948 4210 3952
rect 4238 3948 4242 3952
rect 4246 3948 4250 3952
rect 4278 3948 4282 3952
rect 4318 3948 4322 3952
rect 4358 3948 4362 3952
rect 4374 3948 4378 3952
rect 4414 3948 4418 3952
rect 4446 3948 4450 3952
rect 4462 3948 4466 3952
rect 4486 3948 4490 3952
rect 4526 3948 4530 3952
rect 4542 3948 4546 3952
rect 4566 3958 4570 3962
rect 2070 3938 2074 3942
rect 2078 3938 2082 3942
rect 2134 3938 2138 3942
rect 2158 3938 2162 3942
rect 2190 3938 2194 3942
rect 2550 3938 2554 3942
rect 2662 3938 2666 3942
rect 2686 3938 2690 3942
rect 2774 3938 2778 3942
rect 2782 3938 2786 3942
rect 2806 3938 2810 3942
rect 2830 3938 2834 3942
rect 2838 3938 2842 3942
rect 3126 3938 3130 3942
rect 3158 3938 3162 3942
rect 3230 3938 3234 3942
rect 3238 3938 3242 3942
rect 3302 3938 3306 3942
rect 3318 3938 3322 3942
rect 3358 3938 3362 3942
rect 3406 3938 3410 3942
rect 3518 3938 3522 3942
rect 3550 3938 3554 3942
rect 3614 3938 3618 3942
rect 3622 3938 3626 3942
rect 3654 3938 3658 3942
rect 3662 3938 3666 3942
rect 3694 3938 3698 3942
rect 3734 3938 3738 3942
rect 3774 3938 3778 3942
rect 3806 3938 3810 3942
rect 3862 3938 3866 3942
rect 3878 3938 3882 3942
rect 3902 3938 3906 3942
rect 3934 3938 3938 3942
rect 3950 3938 3954 3942
rect 3958 3938 3962 3942
rect 3974 3938 3978 3942
rect 3990 3938 3994 3942
rect 4126 3938 4130 3942
rect 4174 3938 4178 3942
rect 4190 3938 4194 3942
rect 4214 3938 4218 3942
rect 4238 3938 4242 3942
rect 4254 3938 4258 3942
rect 4294 3938 4298 3942
rect 4310 3938 4314 3942
rect 4350 3938 4354 3942
rect 4366 3938 4370 3942
rect 4382 3938 4386 3942
rect 4438 3938 4442 3942
rect 4470 3938 4474 3942
rect 4502 3938 4506 3942
rect 4518 3938 4522 3942
rect 4534 3938 4538 3942
rect 4582 3938 4586 3942
rect 6 3928 10 3932
rect 38 3928 42 3932
rect 70 3928 74 3932
rect 102 3928 106 3932
rect 214 3928 218 3932
rect 342 3928 346 3932
rect 542 3928 546 3932
rect 702 3928 706 3932
rect 798 3928 802 3932
rect 1406 3928 1410 3932
rect 1502 3928 1506 3932
rect 1510 3928 1514 3932
rect 1606 3928 1610 3932
rect 1830 3928 1834 3932
rect 1870 3928 1874 3932
rect 1958 3928 1962 3932
rect 2094 3928 2098 3932
rect 2326 3928 2330 3932
rect 2342 3928 2346 3932
rect 2726 3928 2730 3932
rect 2806 3928 2810 3932
rect 2862 3928 2866 3932
rect 3310 3928 3314 3932
rect 3462 3928 3466 3932
rect 3670 3928 3674 3932
rect 3822 3928 3826 3932
rect 3830 3928 3834 3932
rect 3838 3928 3842 3932
rect 3902 3928 3906 3932
rect 3950 3928 3954 3932
rect 4038 3928 4042 3932
rect 4334 3928 4338 3932
rect 4398 3928 4402 3932
rect 4486 3928 4490 3932
rect 4598 3928 4602 3932
rect 142 3918 146 3922
rect 206 3918 210 3922
rect 446 3918 450 3922
rect 710 3918 714 3922
rect 830 3918 834 3922
rect 846 3918 850 3922
rect 870 3918 874 3922
rect 1022 3918 1026 3922
rect 1118 3918 1122 3922
rect 1310 3918 1314 3922
rect 1430 3918 1434 3922
rect 1542 3918 1546 3922
rect 1934 3918 1938 3922
rect 1982 3918 1986 3922
rect 2014 3918 2018 3922
rect 2126 3918 2130 3922
rect 2150 3918 2154 3922
rect 2206 3918 2210 3922
rect 2230 3918 2234 3922
rect 2254 3918 2258 3922
rect 2318 3918 2322 3922
rect 2374 3918 2378 3922
rect 2406 3918 2410 3922
rect 2438 3918 2442 3922
rect 2494 3918 2498 3922
rect 2582 3918 2586 3922
rect 2638 3918 2642 3922
rect 2678 3918 2682 3922
rect 2718 3918 2722 3922
rect 2798 3918 2802 3922
rect 2854 3918 2858 3922
rect 2894 3918 2898 3922
rect 3006 3918 3010 3922
rect 3142 3918 3146 3922
rect 3494 3918 3498 3922
rect 3910 3918 3914 3922
rect 3998 3918 4002 3922
rect 4190 3918 4194 3922
rect 4222 3918 4226 3922
rect 4270 3918 4274 3922
rect 4294 3918 4298 3922
rect 4446 3918 4450 3922
rect 1002 3903 1006 3907
rect 1009 3903 1013 3907
rect 2026 3903 2030 3907
rect 2033 3903 2037 3907
rect 3050 3903 3054 3907
rect 3057 3903 3061 3907
rect 4082 3903 4086 3907
rect 4089 3903 4093 3907
rect 110 3888 114 3892
rect 230 3888 234 3892
rect 326 3888 330 3892
rect 374 3888 378 3892
rect 382 3888 386 3892
rect 430 3888 434 3892
rect 574 3888 578 3892
rect 614 3888 618 3892
rect 742 3888 746 3892
rect 934 3888 938 3892
rect 1150 3888 1154 3892
rect 1502 3888 1506 3892
rect 1526 3888 1530 3892
rect 1622 3888 1626 3892
rect 1734 3888 1738 3892
rect 1790 3888 1794 3892
rect 3166 3888 3170 3892
rect 3174 3888 3178 3892
rect 3454 3888 3458 3892
rect 3462 3888 3466 3892
rect 3750 3888 3754 3892
rect 3758 3888 3762 3892
rect 3798 3888 3802 3892
rect 3814 3888 3818 3892
rect 3926 3888 3930 3892
rect 4054 3888 4058 3892
rect 4390 3888 4394 3892
rect 4438 3888 4442 3892
rect 4510 3888 4514 3892
rect 6 3878 10 3882
rect 694 3878 698 3882
rect 718 3878 722 3882
rect 774 3878 778 3882
rect 790 3878 794 3882
rect 798 3878 802 3882
rect 854 3878 858 3882
rect 910 3878 914 3882
rect 982 3878 986 3882
rect 1270 3878 1274 3882
rect 1318 3878 1322 3882
rect 1438 3878 1442 3882
rect 1958 3878 1962 3882
rect 1974 3878 1978 3882
rect 2390 3878 2394 3882
rect 2438 3878 2442 3882
rect 2494 3878 2498 3882
rect 2726 3878 2730 3882
rect 2750 3878 2754 3882
rect 2982 3878 2986 3882
rect 3142 3878 3146 3882
rect 3326 3878 3330 3882
rect 30 3868 34 3872
rect 158 3868 162 3872
rect 214 3868 218 3872
rect 270 3868 274 3872
rect 318 3868 322 3872
rect 342 3866 346 3870
rect 350 3868 354 3872
rect 358 3868 362 3872
rect 398 3866 402 3870
rect 414 3868 418 3872
rect 462 3868 466 3872
rect 518 3868 522 3872
rect 582 3868 586 3872
rect 630 3868 634 3872
rect 638 3868 642 3872
rect 686 3868 690 3872
rect 710 3868 714 3872
rect 918 3868 922 3872
rect 934 3868 938 3872
rect 1038 3868 1042 3872
rect 1070 3868 1074 3872
rect 1158 3868 1162 3872
rect 1190 3868 1194 3872
rect 1214 3868 1218 3872
rect 1254 3868 1258 3872
rect 1270 3868 1274 3872
rect 1326 3868 1330 3872
rect 1606 3868 1610 3872
rect 1718 3868 1722 3872
rect 1726 3868 1730 3872
rect 1758 3868 1762 3872
rect 1902 3868 1906 3872
rect 1926 3868 1930 3872
rect 2022 3868 2026 3872
rect 2110 3868 2114 3872
rect 2174 3868 2178 3872
rect 2438 3868 2442 3872
rect 2462 3868 2466 3872
rect 2646 3868 2650 3872
rect 3422 3878 3426 3882
rect 3702 3878 3706 3882
rect 3790 3878 3794 3882
rect 3878 3878 3882 3882
rect 3942 3878 3946 3882
rect 4046 3878 4050 3882
rect 4446 3878 4450 3882
rect 2894 3868 2898 3872
rect 2910 3868 2914 3872
rect 3206 3868 3210 3872
rect 3310 3868 3314 3872
rect 3398 3868 3402 3872
rect 3430 3868 3434 3872
rect 46 3859 50 3863
rect 78 3858 82 3862
rect 142 3859 146 3863
rect 302 3858 306 3862
rect 510 3859 514 3863
rect 710 3858 714 3862
rect 758 3858 762 3862
rect 838 3858 842 3862
rect 870 3858 874 3862
rect 950 3858 954 3862
rect 1102 3858 1106 3862
rect 1166 3858 1170 3862
rect 1190 3858 1194 3862
rect 1206 3858 1210 3862
rect 1222 3858 1226 3862
rect 1278 3858 1282 3862
rect 1294 3858 1298 3862
rect 1310 3858 1314 3862
rect 1374 3858 1378 3862
rect 1382 3858 1386 3862
rect 1406 3858 1410 3862
rect 1438 3859 1442 3863
rect 1462 3858 1466 3862
rect 1558 3858 1562 3862
rect 1590 3859 1594 3863
rect 1662 3858 1666 3862
rect 1686 3859 1690 3863
rect 1774 3858 1778 3862
rect 1830 3858 1834 3862
rect 1862 3859 1866 3863
rect 1910 3858 1914 3862
rect 1950 3858 1954 3862
rect 1998 3858 2002 3862
rect 374 3848 378 3852
rect 670 3848 674 3852
rect 862 3848 866 3852
rect 902 3848 906 3852
rect 934 3848 938 3852
rect 1182 3848 1186 3852
rect 1230 3848 1234 3852
rect 1790 3848 1794 3852
rect 1894 3848 1898 3852
rect 206 3838 210 3842
rect 814 3838 818 3842
rect 878 3838 882 3842
rect 1342 3838 1346 3842
rect 1734 3838 1738 3842
rect 2006 3838 2010 3842
rect 2046 3838 2050 3842
rect 2086 3858 2090 3862
rect 2118 3858 2122 3862
rect 2150 3858 2154 3862
rect 2182 3858 2186 3862
rect 2214 3858 2218 3862
rect 2246 3858 2250 3862
rect 2270 3858 2274 3862
rect 2294 3858 2298 3862
rect 2342 3858 2346 3862
rect 2358 3858 2362 3862
rect 2414 3858 2418 3862
rect 2470 3858 2474 3862
rect 2518 3858 2522 3862
rect 2574 3858 2578 3862
rect 2606 3858 2610 3862
rect 2062 3848 2066 3852
rect 2094 3848 2098 3852
rect 2126 3848 2130 3852
rect 2158 3848 2162 3852
rect 2190 3848 2194 3852
rect 2222 3848 2226 3852
rect 2254 3848 2258 3852
rect 2350 3848 2354 3852
rect 2374 3848 2378 3852
rect 2502 3848 2506 3852
rect 2566 3848 2570 3852
rect 2598 3848 2602 3852
rect 2630 3848 2634 3852
rect 2078 3838 2082 3842
rect 2110 3838 2114 3842
rect 2142 3838 2146 3842
rect 2174 3838 2178 3842
rect 2206 3838 2210 3842
rect 2238 3838 2242 3842
rect 2262 3838 2266 3842
rect 2334 3838 2338 3842
rect 2422 3838 2426 3842
rect 2462 3838 2466 3842
rect 2550 3838 2554 3842
rect 2614 3838 2618 3842
rect 2662 3838 2666 3842
rect 2702 3858 2706 3862
rect 2750 3858 2754 3862
rect 2782 3858 2786 3862
rect 2814 3858 2818 3862
rect 2838 3858 2842 3862
rect 2878 3858 2882 3862
rect 3438 3866 3442 3870
rect 3542 3868 3546 3872
rect 3574 3868 3578 3872
rect 3598 3868 3602 3872
rect 3670 3868 3674 3872
rect 3678 3868 3682 3872
rect 2918 3858 2922 3862
rect 2942 3858 2946 3862
rect 3006 3858 3010 3862
rect 3022 3858 3026 3862
rect 3038 3858 3042 3862
rect 3086 3858 3090 3862
rect 3102 3858 3106 3862
rect 3118 3858 3122 3862
rect 3230 3858 3234 3862
rect 3294 3859 3298 3863
rect 3734 3866 3738 3870
rect 3782 3868 3786 3872
rect 3838 3868 3842 3872
rect 3846 3868 3850 3872
rect 3918 3868 3922 3872
rect 3934 3868 3938 3872
rect 3982 3868 3986 3872
rect 4014 3868 4018 3872
rect 4038 3868 4042 3872
rect 4062 3868 4066 3872
rect 4102 3868 4106 3872
rect 4142 3868 4146 3872
rect 4158 3868 4162 3872
rect 4214 3868 4218 3872
rect 4230 3868 4234 3872
rect 4270 3868 4274 3872
rect 4302 3868 4306 3872
rect 4334 3868 4338 3872
rect 4430 3868 4434 3872
rect 4462 3868 4466 3872
rect 4478 3868 4482 3872
rect 4502 3868 4506 3872
rect 4534 3868 4538 3872
rect 4558 3868 4562 3872
rect 3406 3858 3410 3862
rect 3518 3858 3522 3862
rect 3582 3858 3586 3862
rect 3678 3858 3682 3862
rect 3702 3858 3706 3862
rect 3718 3858 3722 3862
rect 3774 3858 3778 3862
rect 3806 3858 3810 3862
rect 3830 3858 3834 3862
rect 3846 3858 3850 3862
rect 3894 3858 3898 3862
rect 3910 3858 3914 3862
rect 3934 3858 3938 3862
rect 3974 3858 3978 3862
rect 3990 3858 3994 3862
rect 4030 3858 4034 3862
rect 4078 3858 4082 3862
rect 4166 3858 4170 3862
rect 4198 3858 4202 3862
rect 4206 3858 4210 3862
rect 4222 3858 4226 3862
rect 4238 3858 4242 3862
rect 4270 3858 4274 3862
rect 4294 3858 4298 3862
rect 4334 3858 4338 3862
rect 4374 3858 4378 3862
rect 4406 3858 4410 3862
rect 4454 3858 4458 3862
rect 4486 3858 4490 3862
rect 4494 3858 4498 3862
rect 4526 3858 4530 3862
rect 4590 3858 4594 3862
rect 2678 3848 2682 3852
rect 2750 3848 2754 3852
rect 2790 3848 2794 3852
rect 2822 3848 2826 3852
rect 2830 3848 2834 3852
rect 2886 3848 2890 3852
rect 2894 3848 2898 3852
rect 3030 3848 3034 3852
rect 3078 3848 3082 3852
rect 3110 3848 3114 3852
rect 3398 3848 3402 3852
rect 3598 3848 3602 3852
rect 3758 3848 3762 3852
rect 3814 3848 3818 3852
rect 3870 3848 3874 3852
rect 3894 3848 3898 3852
rect 4006 3848 4010 3852
rect 4062 3848 4066 3852
rect 4078 3848 4082 3852
rect 4126 3848 4130 3852
rect 4246 3848 4250 3852
rect 4278 3848 4282 3852
rect 4310 3848 4314 3852
rect 4366 3848 4370 3852
rect 2702 3838 2706 3842
rect 2742 3838 2746 3842
rect 2774 3838 2778 3842
rect 2806 3838 2810 3842
rect 2846 3838 2850 3842
rect 2870 3838 2874 3842
rect 3014 3838 3018 3842
rect 3046 3838 3050 3842
rect 3070 3838 3074 3842
rect 3126 3838 3130 3842
rect 2534 3828 2538 3832
rect 2638 3828 2642 3832
rect 3974 3828 3978 3832
rect 14 3818 18 3822
rect 782 3818 786 3822
rect 966 3818 970 3822
rect 1358 3818 1362 3822
rect 1390 3818 1394 3822
rect 1934 3818 1938 3822
rect 1966 3818 1970 3822
rect 2054 3818 2058 3822
rect 2150 3818 2154 3822
rect 2214 3818 2218 3822
rect 2246 3818 2250 3822
rect 2286 3818 2290 3822
rect 2310 3818 2314 3822
rect 2342 3818 2346 3822
rect 2430 3818 2434 3822
rect 2590 3818 2594 3822
rect 2622 3818 2626 3822
rect 2670 3818 2674 3822
rect 2782 3818 2786 3822
rect 2798 3818 2802 3822
rect 2854 3818 2858 3822
rect 2878 3818 2882 3822
rect 2934 3818 2938 3822
rect 2974 3818 2978 3822
rect 3038 3818 3042 3822
rect 3118 3818 3122 3822
rect 3390 3818 3394 3822
rect 3614 3818 3618 3822
rect 4142 3818 4146 3822
rect 4462 3818 4466 3822
rect 4542 3818 4546 3822
rect 498 3803 502 3807
rect 505 3803 509 3807
rect 1522 3803 1526 3807
rect 1529 3803 1533 3807
rect 2546 3803 2550 3807
rect 2553 3803 2557 3807
rect 3570 3803 3574 3807
rect 3577 3803 3581 3807
rect 238 3788 242 3792
rect 334 3788 338 3792
rect 430 3788 434 3792
rect 614 3788 618 3792
rect 902 3788 906 3792
rect 1126 3788 1130 3792
rect 1174 3788 1178 3792
rect 1198 3788 1202 3792
rect 1662 3788 1666 3792
rect 1878 3788 1882 3792
rect 1958 3788 1962 3792
rect 2118 3788 2122 3792
rect 2150 3788 2154 3792
rect 2190 3788 2194 3792
rect 2334 3788 2338 3792
rect 2414 3788 2418 3792
rect 2750 3788 2754 3792
rect 2774 3788 2778 3792
rect 2854 3788 2858 3792
rect 3766 3788 3770 3792
rect 3862 3788 3866 3792
rect 3926 3788 3930 3792
rect 4190 3788 4194 3792
rect 4214 3788 4218 3792
rect 4438 3788 4442 3792
rect 1694 3778 1698 3782
rect 2126 3778 2130 3782
rect 2374 3778 2378 3782
rect 1510 3768 1514 3772
rect 2262 3768 2266 3772
rect 2326 3768 2330 3772
rect 2702 3768 2706 3772
rect 2766 3768 2770 3772
rect 2862 3768 2866 3772
rect 2966 3768 2970 3772
rect 3030 3768 3034 3772
rect 3718 3768 3722 3772
rect 4510 3768 4514 3772
rect 38 3757 42 3761
rect 654 3758 658 3762
rect 774 3758 778 3762
rect 1326 3758 1330 3762
rect 1446 3758 1450 3762
rect 1678 3758 1682 3762
rect 94 3748 98 3752
rect 126 3748 130 3752
rect 142 3748 146 3752
rect 174 3747 178 3751
rect 270 3747 274 3751
rect 366 3747 370 3751
rect 558 3748 562 3752
rect 750 3748 754 3752
rect 766 3748 770 3752
rect 790 3748 794 3752
rect 838 3747 842 3751
rect 966 3748 970 3752
rect 1062 3747 1066 3751
rect 1134 3748 1138 3752
rect 1166 3748 1170 3752
rect 1190 3748 1194 3752
rect 1262 3748 1266 3752
rect 1294 3747 1298 3751
rect 1398 3748 1402 3752
rect 1406 3748 1410 3752
rect 1438 3748 1442 3752
rect 1478 3748 1482 3752
rect 1542 3748 1546 3752
rect 1574 3747 1578 3751
rect 1678 3748 1682 3752
rect 1742 3748 1746 3752
rect 1774 3747 1778 3751
rect 1814 3748 1818 3752
rect 1838 3758 1842 3762
rect 1854 3748 1858 3752
rect 1878 3748 1882 3752
rect 1902 3758 1906 3762
rect 1974 3758 1978 3762
rect 2174 3758 2178 3762
rect 2310 3758 2314 3762
rect 2342 3758 2346 3762
rect 2494 3758 2498 3762
rect 2518 3758 2522 3762
rect 2526 3758 2530 3762
rect 2606 3758 2610 3762
rect 2686 3758 2690 3762
rect 2806 3758 2810 3762
rect 2894 3758 2898 3762
rect 2950 3758 2954 3762
rect 2990 3758 2994 3762
rect 3014 3758 3018 3762
rect 3038 3758 3042 3762
rect 3094 3758 3098 3762
rect 3118 3758 3122 3762
rect 3142 3758 3146 3762
rect 3254 3758 3258 3762
rect 3270 3758 3274 3762
rect 3406 3758 3410 3762
rect 3414 3758 3418 3762
rect 3446 3758 3450 3762
rect 1918 3748 1922 3752
rect 2014 3748 2018 3752
rect 2054 3747 2058 3751
rect 2078 3748 2082 3752
rect 2222 3748 2226 3752
rect 2230 3748 2234 3752
rect 2278 3748 2282 3752
rect 2318 3748 2322 3752
rect 2390 3748 2394 3752
rect 2398 3748 2402 3752
rect 2454 3748 2458 3752
rect 2542 3748 2546 3752
rect 2710 3748 2714 3752
rect 2774 3748 2778 3752
rect 2854 3748 2858 3752
rect 3110 3748 3114 3752
rect 3126 3748 3130 3752
rect 3190 3748 3194 3752
rect 3222 3748 3226 3752
rect 3270 3748 3274 3752
rect 3326 3747 3330 3751
rect 3358 3748 3362 3752
rect 3398 3748 3402 3752
rect 3446 3748 3450 3752
rect 3462 3748 3466 3752
rect 3518 3747 3522 3751
rect 3542 3748 3546 3752
rect 3854 3758 3858 3762
rect 4110 3758 4114 3762
rect 4142 3758 4146 3762
rect 4294 3758 4298 3762
rect 4310 3758 4314 3762
rect 4358 3758 4362 3762
rect 4478 3758 4482 3762
rect 4526 3758 4530 3762
rect 4582 3758 4586 3762
rect 3734 3748 3738 3752
rect 3798 3748 3802 3752
rect 3806 3748 3810 3752
rect 3838 3748 3842 3752
rect 3846 3748 3850 3752
rect 3878 3748 3882 3752
rect 3926 3748 3930 3752
rect 3934 3748 3938 3752
rect 3966 3748 3970 3752
rect 3974 3748 3978 3752
rect 4006 3748 4010 3752
rect 4014 3748 4018 3752
rect 4054 3748 4058 3752
rect 4086 3748 4090 3752
rect 4126 3748 4130 3752
rect 4158 3748 4162 3752
rect 4174 3748 4178 3752
rect 4230 3748 4234 3752
rect 4262 3748 4266 3752
rect 4278 3748 4282 3752
rect 4326 3748 4330 3752
rect 4334 3748 4338 3752
rect 4366 3748 4370 3752
rect 4398 3748 4402 3752
rect 4406 3748 4410 3752
rect 4462 3748 4466 3752
rect 4486 3748 4490 3752
rect 4518 3748 4522 3752
rect 4566 3748 4570 3752
rect 22 3738 26 3742
rect 62 3738 66 3742
rect 118 3738 122 3742
rect 286 3738 290 3742
rect 502 3738 506 3742
rect 622 3738 626 3742
rect 670 3738 674 3742
rect 678 3738 682 3742
rect 726 3738 730 3742
rect 758 3738 762 3742
rect 774 3738 778 3742
rect 822 3738 826 3742
rect 934 3738 938 3742
rect 1046 3738 1050 3742
rect 1070 3738 1074 3742
rect 1142 3738 1146 3742
rect 1158 3738 1162 3742
rect 1198 3738 1202 3742
rect 1214 3738 1218 3742
rect 1358 3738 1362 3742
rect 1374 3738 1378 3742
rect 1414 3738 1418 3742
rect 1422 3738 1426 3742
rect 1430 3738 1434 3742
rect 1470 3738 1474 3742
rect 1606 3738 1610 3742
rect 1806 3738 1810 3742
rect 1862 3738 1866 3742
rect 1870 3738 1874 3742
rect 1934 3738 1938 3742
rect 1950 3738 1954 3742
rect 1990 3738 1994 3742
rect 2158 3738 2162 3742
rect 2198 3738 2202 3742
rect 2262 3738 2266 3742
rect 2358 3738 2362 3742
rect 2422 3738 2426 3742
rect 2510 3738 2514 3742
rect 2534 3738 2538 3742
rect 2822 3738 2826 3742
rect 2878 3738 2882 3742
rect 2886 3738 2890 3742
rect 2910 3738 2914 3742
rect 2934 3738 2938 3742
rect 2942 3738 2946 3742
rect 2966 3738 2970 3742
rect 2974 3738 2978 3742
rect 2998 3738 3002 3742
rect 3022 3738 3026 3742
rect 3102 3738 3106 3742
rect 3150 3738 3154 3742
rect 3166 3738 3170 3742
rect 3246 3738 3250 3742
rect 3310 3738 3314 3742
rect 3414 3738 3418 3742
rect 3438 3738 3442 3742
rect 3534 3738 3538 3742
rect 3606 3738 3610 3742
rect 3710 3738 3714 3742
rect 3734 3738 3738 3742
rect 3830 3738 3834 3742
rect 3942 3738 3946 3742
rect 3958 3738 3962 3742
rect 3982 3738 3986 3742
rect 3998 3738 4002 3742
rect 4022 3738 4026 3742
rect 4038 3738 4042 3742
rect 4078 3738 4082 3742
rect 4134 3738 4138 3742
rect 4166 3738 4170 3742
rect 4206 3738 4210 3742
rect 4238 3738 4242 3742
rect 4270 3738 4274 3742
rect 4334 3738 4338 3742
rect 4374 3738 4378 3742
rect 4382 3738 4386 3742
rect 4398 3738 4402 3742
rect 4422 3738 4426 3742
rect 4454 3738 4458 3742
rect 4486 3738 4490 3742
rect 4510 3738 4514 3742
rect 4550 3738 4554 3742
rect 6 3728 10 3732
rect 86 3728 90 3732
rect 126 3728 130 3732
rect 174 3728 178 3732
rect 366 3728 370 3732
rect 550 3728 554 3732
rect 734 3728 738 3732
rect 870 3728 874 3732
rect 918 3728 922 3732
rect 1182 3728 1186 3732
rect 1358 3728 1362 3732
rect 1478 3728 1482 3732
rect 1494 3728 1498 3732
rect 1678 3728 1682 3732
rect 1934 3728 1938 3732
rect 2134 3728 2138 3732
rect 2142 3728 2146 3732
rect 2182 3728 2186 3732
rect 2262 3728 2266 3732
rect 2734 3728 2738 3732
rect 2742 3728 2746 3732
rect 2798 3728 2802 3732
rect 2830 3728 2834 3732
rect 2918 3728 2922 3732
rect 3046 3728 3050 3732
rect 3134 3728 3138 3732
rect 3214 3728 3218 3732
rect 3294 3728 3298 3732
rect 3486 3728 3490 3732
rect 3782 3728 3786 3732
rect 3806 3728 3810 3732
rect 3822 3728 3826 3732
rect 3870 3728 3874 3732
rect 3894 3728 3898 3732
rect 3910 3728 3914 3732
rect 4446 3728 4450 3732
rect 126 3718 130 3722
rect 446 3718 450 3722
rect 710 3718 714 3722
rect 806 3718 810 3722
rect 910 3718 914 3722
rect 1014 3718 1018 3722
rect 1150 3718 1154 3722
rect 1830 3718 1834 3722
rect 2174 3718 2178 3722
rect 2294 3718 2298 3722
rect 2342 3718 2346 3722
rect 2446 3718 2450 3722
rect 2478 3718 2482 3722
rect 2502 3718 2506 3722
rect 2606 3718 2610 3722
rect 2622 3718 2626 3722
rect 2678 3718 2682 3722
rect 2702 3718 2706 3722
rect 2806 3718 2810 3722
rect 2902 3718 2906 3722
rect 2926 3718 2930 3722
rect 2990 3718 2994 3722
rect 3014 3718 3018 3722
rect 3094 3718 3098 3722
rect 3174 3718 3178 3722
rect 3390 3718 3394 3722
rect 3430 3718 3434 3722
rect 3590 3718 3594 3722
rect 3662 3718 3666 3722
rect 3814 3718 3818 3722
rect 3958 3718 3962 3722
rect 3998 3718 4002 3722
rect 4038 3718 4042 3722
rect 4070 3718 4074 3722
rect 3214 3708 3218 3712
rect 3294 3708 3298 3712
rect 1002 3703 1006 3707
rect 1009 3703 1013 3707
rect 2026 3703 2030 3707
rect 2033 3703 2037 3707
rect 3050 3703 3054 3707
rect 3057 3703 3061 3707
rect 4082 3703 4086 3707
rect 4089 3703 4093 3707
rect 3358 3698 3362 3702
rect 3486 3698 3490 3702
rect 3774 3698 3778 3702
rect 254 3688 258 3692
rect 422 3688 426 3692
rect 534 3688 538 3692
rect 838 3688 842 3692
rect 966 3688 970 3692
rect 990 3688 994 3692
rect 1110 3688 1114 3692
rect 1166 3688 1170 3692
rect 1310 3688 1314 3692
rect 1454 3688 1458 3692
rect 1654 3688 1658 3692
rect 1758 3688 1762 3692
rect 1854 3688 1858 3692
rect 1886 3688 1890 3692
rect 2006 3688 2010 3692
rect 2030 3688 2034 3692
rect 2358 3688 2362 3692
rect 2966 3688 2970 3692
rect 3062 3688 3066 3692
rect 3494 3688 3498 3692
rect 3782 3688 3786 3692
rect 4398 3688 4402 3692
rect 4430 3688 4434 3692
rect 6 3678 10 3682
rect 38 3678 42 3682
rect 46 3678 50 3682
rect 70 3678 74 3682
rect 142 3678 146 3682
rect 454 3678 458 3682
rect 590 3678 594 3682
rect 662 3678 666 3682
rect 734 3678 738 3682
rect 1046 3678 1050 3682
rect 1158 3678 1162 3682
rect 1302 3678 1306 3682
rect 2158 3678 2162 3682
rect 2238 3678 2242 3682
rect 2318 3678 2322 3682
rect 2326 3678 2330 3682
rect 2334 3678 2338 3682
rect 2342 3678 2346 3682
rect 2398 3678 2402 3682
rect 2446 3678 2450 3682
rect 2710 3678 2714 3682
rect 2758 3678 2762 3682
rect 2774 3678 2778 3682
rect 2894 3678 2898 3682
rect 2902 3678 2906 3682
rect 2974 3678 2978 3682
rect 3022 3678 3026 3682
rect 3358 3678 3362 3682
rect 3486 3678 3490 3682
rect 3774 3678 3778 3682
rect 102 3668 106 3672
rect 142 3668 146 3672
rect 158 3668 162 3672
rect 174 3668 178 3672
rect 262 3668 266 3672
rect 326 3668 330 3672
rect 342 3668 346 3672
rect 366 3668 370 3672
rect 630 3668 634 3672
rect 870 3668 874 3672
rect 918 3668 922 3672
rect 1142 3668 1146 3672
rect 1214 3668 1218 3672
rect 1246 3668 1250 3672
rect 1286 3668 1290 3672
rect 1358 3668 1362 3672
rect 1430 3668 1434 3672
rect 1446 3668 1450 3672
rect 1742 3668 1746 3672
rect 1806 3668 1810 3672
rect 1878 3668 1882 3672
rect 1934 3668 1938 3672
rect 1982 3668 1986 3672
rect 2078 3668 2082 3672
rect 2350 3668 2354 3672
rect 2534 3668 2538 3672
rect 2590 3668 2594 3672
rect 2638 3668 2642 3672
rect 2726 3668 2730 3672
rect 2902 3668 2906 3672
rect 2950 3668 2954 3672
rect 3038 3668 3042 3672
rect 3174 3668 3178 3672
rect 3310 3668 3314 3672
rect 3382 3668 3386 3672
rect 3414 3668 3418 3672
rect 3454 3668 3458 3672
rect 3534 3668 3538 3672
rect 3614 3668 3618 3672
rect 3726 3668 3730 3672
rect 3990 3668 3994 3672
rect 4022 3668 4026 3672
rect 4118 3668 4122 3672
rect 4150 3668 4154 3672
rect 4182 3668 4186 3672
rect 4214 3668 4218 3672
rect 4262 3668 4266 3672
rect 4286 3668 4290 3672
rect 4318 3668 4322 3672
rect 4486 3668 4490 3672
rect 4502 3668 4506 3672
rect 4542 3668 4546 3672
rect 4574 3668 4578 3672
rect 46 3658 50 3662
rect 134 3658 138 3662
rect 190 3659 194 3663
rect 222 3658 226 3662
rect 374 3658 378 3662
rect 454 3659 458 3663
rect 542 3658 546 3662
rect 582 3658 586 3662
rect 614 3658 618 3662
rect 662 3659 666 3663
rect 774 3659 778 3663
rect 806 3658 810 3662
rect 854 3658 858 3662
rect 862 3658 866 3662
rect 910 3658 914 3662
rect 974 3658 978 3662
rect 1054 3658 1058 3662
rect 1230 3659 1234 3663
rect 1374 3659 1378 3663
rect 1518 3659 1522 3663
rect 1590 3659 1594 3663
rect 1622 3658 1626 3662
rect 1726 3659 1730 3663
rect 1822 3659 1826 3663
rect 1878 3658 1882 3662
rect 1950 3659 1954 3663
rect 1990 3658 1994 3662
rect 2094 3659 2098 3663
rect 2134 3658 2138 3662
rect 2190 3658 2194 3662
rect 2214 3658 2218 3662
rect 2270 3658 2274 3662
rect 2302 3658 2306 3662
rect 2382 3658 2386 3662
rect 2414 3658 2418 3662
rect 2462 3658 2466 3662
rect 2494 3658 2498 3662
rect 2566 3658 2570 3662
rect 2582 3658 2586 3662
rect 2654 3658 2658 3662
rect 2694 3658 2698 3662
rect 2750 3658 2754 3662
rect 2798 3658 2802 3662
rect 2830 3658 2834 3662
rect 2870 3658 2874 3662
rect 2934 3658 2938 3662
rect 2998 3658 3002 3662
rect 3038 3658 3042 3662
rect 3086 3658 3090 3662
rect 3118 3658 3122 3662
rect 3134 3658 3138 3662
rect 3158 3658 3162 3662
rect 3214 3658 3218 3662
rect 3246 3658 3250 3662
rect 3262 3658 3266 3662
rect 3294 3658 3298 3662
rect 3334 3658 3338 3662
rect 3438 3658 3442 3662
rect 3462 3658 3466 3662
rect 3550 3658 3554 3662
rect 3630 3659 3634 3663
rect 3702 3658 3706 3662
rect 3750 3658 3754 3662
rect 3814 3658 3818 3662
rect 3830 3658 3834 3662
rect 3902 3659 3906 3663
rect 4030 3658 4034 3662
rect 4070 3658 4074 3662
rect 4110 3658 4114 3662
rect 4142 3658 4146 3662
rect 4174 3658 4178 3662
rect 4206 3658 4210 3662
rect 4254 3658 4258 3662
rect 4286 3658 4290 3662
rect 4310 3658 4314 3662
rect 4326 3658 4330 3662
rect 4374 3658 4378 3662
rect 4382 3658 4386 3662
rect 4414 3658 4418 3662
rect 4446 3658 4450 3662
rect 4478 3658 4482 3662
rect 4518 3658 4522 3662
rect 4534 3658 4538 3662
rect 4542 3658 4546 3662
rect 118 3649 122 3653
rect 630 3648 634 3652
rect 846 3648 850 3652
rect 1118 3648 1122 3652
rect 1262 3648 1266 3652
rect 1406 3648 1410 3652
rect 2126 3648 2130 3652
rect 2198 3648 2202 3652
rect 2206 3648 2210 3652
rect 2278 3648 2282 3652
rect 2310 3648 2314 3652
rect 2366 3648 2370 3652
rect 2374 3648 2378 3652
rect 2454 3648 2458 3652
rect 2486 3648 2490 3652
rect 2518 3648 2522 3652
rect 2558 3648 2562 3652
rect 2638 3648 2642 3652
rect 2646 3648 2650 3652
rect 2702 3648 2706 3652
rect 2790 3648 2794 3652
rect 2814 3648 2818 3652
rect 2822 3648 2826 3652
rect 2942 3648 2946 3652
rect 2966 3648 2970 3652
rect 3054 3648 3058 3652
rect 3078 3648 3082 3652
rect 3110 3648 3114 3652
rect 3166 3648 3170 3652
rect 3182 3648 3186 3652
rect 3190 3648 3194 3652
rect 3222 3648 3226 3652
rect 3254 3648 3258 3652
rect 3366 3648 3370 3652
rect 3446 3648 3450 3652
rect 3734 3648 3738 3652
rect 4014 3648 4018 3652
rect 4030 3648 4034 3652
rect 4046 3648 4050 3652
rect 4094 3648 4098 3652
rect 4126 3648 4130 3652
rect 4158 3648 4162 3652
rect 4190 3648 4194 3652
rect 4518 3648 4522 3652
rect 726 3638 730 3642
rect 822 3638 826 3642
rect 1854 3638 1858 3642
rect 2006 3638 2010 3642
rect 2142 3638 2146 3642
rect 2158 3638 2162 3642
rect 2182 3638 2186 3642
rect 2190 3638 2194 3642
rect 2222 3638 2226 3642
rect 2262 3638 2266 3642
rect 2294 3638 2298 3642
rect 2390 3638 2394 3642
rect 2414 3638 2418 3642
rect 2470 3638 2474 3642
rect 2502 3638 2506 3642
rect 2534 3638 2538 3642
rect 2574 3638 2578 3642
rect 2662 3638 2666 3642
rect 2686 3638 2690 3642
rect 2734 3638 2738 3642
rect 2798 3638 2802 3642
rect 2806 3638 2810 3642
rect 2838 3638 2842 3642
rect 2862 3638 2866 3642
rect 2926 3638 2930 3642
rect 3006 3638 3010 3642
rect 3070 3638 3074 3642
rect 3126 3638 3130 3642
rect 3150 3638 3154 3642
rect 3206 3638 3210 3642
rect 3238 3638 3242 3642
rect 3406 3638 3410 3642
rect 3950 3638 3954 3642
rect 4502 3638 4506 3642
rect 3214 3628 3218 3632
rect 3278 3628 3282 3632
rect 742 3618 746 3622
rect 990 3618 994 3622
rect 1662 3618 1666 3622
rect 2134 3618 2138 3622
rect 2190 3618 2194 3622
rect 2302 3618 2306 3622
rect 2422 3618 2426 3622
rect 2478 3618 2482 3622
rect 2494 3618 2498 3622
rect 2654 3618 2658 3622
rect 2678 3618 2682 3622
rect 2766 3618 2770 3622
rect 2830 3618 2834 3622
rect 2870 3618 2874 3622
rect 2934 3618 2938 3622
rect 3014 3618 3018 3622
rect 3102 3618 3106 3622
rect 3142 3618 3146 3622
rect 3246 3618 3250 3622
rect 3334 3618 3338 3622
rect 3694 3618 3698 3622
rect 3750 3618 3754 3622
rect 4326 3618 4330 3622
rect 4358 3618 4362 3622
rect 4462 3618 4466 3622
rect 498 3603 502 3607
rect 505 3603 509 3607
rect 1522 3603 1526 3607
rect 1529 3603 1533 3607
rect 2546 3603 2550 3607
rect 2553 3603 2557 3607
rect 3570 3603 3574 3607
rect 3577 3603 3581 3607
rect 382 3588 386 3592
rect 1238 3588 1242 3592
rect 1406 3588 1410 3592
rect 1622 3588 1626 3592
rect 1886 3588 1890 3592
rect 1982 3588 1986 3592
rect 2022 3588 2026 3592
rect 2110 3588 2114 3592
rect 2198 3588 2202 3592
rect 2318 3588 2322 3592
rect 2462 3588 2466 3592
rect 2518 3588 2522 3592
rect 2846 3588 2850 3592
rect 2942 3588 2946 3592
rect 2990 3588 2994 3592
rect 3078 3588 3082 3592
rect 3406 3588 3410 3592
rect 3718 3588 3722 3592
rect 1918 3578 1922 3582
rect 2534 3578 2538 3582
rect 3606 3578 3610 3582
rect 190 3568 194 3572
rect 286 3568 290 3572
rect 886 3568 890 3572
rect 1142 3568 1146 3572
rect 1750 3568 1754 3572
rect 1942 3568 1946 3572
rect 2454 3568 2458 3572
rect 2502 3568 2506 3572
rect 2854 3568 2858 3572
rect 2878 3568 2882 3572
rect 2950 3568 2954 3572
rect 2998 3568 3002 3572
rect 3742 3568 3746 3572
rect 3870 3568 3874 3572
rect 534 3558 538 3562
rect 734 3558 738 3562
rect 790 3558 794 3562
rect 1382 3558 1386 3562
rect 1862 3558 1866 3562
rect 1902 3558 1906 3562
rect 22 3548 26 3552
rect 94 3548 98 3552
rect 126 3547 130 3551
rect 158 3548 162 3552
rect 230 3548 234 3552
rect 318 3547 322 3551
rect 342 3548 346 3552
rect 406 3548 410 3552
rect 438 3548 442 3552
rect 670 3548 674 3552
rect 774 3548 778 3552
rect 846 3548 850 3552
rect 1078 3547 1082 3551
rect 1174 3547 1178 3551
rect 1246 3548 1250 3552
rect 1262 3548 1266 3552
rect 1350 3547 1354 3551
rect 1398 3548 1402 3552
rect 1438 3548 1442 3552
rect 1446 3548 1450 3552
rect 1518 3547 1522 3551
rect 1630 3548 1634 3552
rect 1686 3548 1690 3552
rect 1718 3547 1722 3551
rect 1782 3548 1786 3552
rect 1814 3547 1818 3551
rect 1918 3548 1922 3552
rect 1998 3558 2002 3562
rect 2006 3558 2010 3562
rect 2126 3558 2130 3562
rect 2142 3558 2146 3562
rect 2294 3558 2298 3562
rect 2430 3558 2434 3562
rect 2438 3558 2442 3562
rect 2470 3558 2474 3562
rect 2494 3558 2498 3562
rect 2598 3558 2602 3562
rect 2638 3558 2642 3562
rect 2646 3558 2650 3562
rect 2670 3558 2674 3562
rect 2694 3558 2698 3562
rect 2774 3558 2778 3562
rect 2814 3558 2818 3562
rect 3014 3558 3018 3562
rect 3086 3558 3090 3562
rect 3110 3558 3114 3562
rect 3150 3558 3154 3562
rect 3190 3558 3194 3562
rect 3230 3558 3234 3562
rect 3286 3558 3290 3562
rect 3310 3558 3314 3562
rect 3334 3558 3338 3562
rect 3390 3558 3394 3562
rect 3430 3558 3434 3562
rect 3438 3558 3442 3562
rect 3462 3558 3466 3562
rect 3510 3558 3514 3562
rect 3726 3558 3730 3562
rect 4238 3558 4242 3562
rect 4510 3558 4514 3562
rect 4534 3558 4538 3562
rect 1958 3548 1962 3552
rect 1982 3548 1986 3552
rect 2022 3548 2026 3552
rect 2054 3548 2058 3552
rect 2070 3548 2074 3552
rect 2110 3548 2114 3552
rect 2126 3548 2130 3552
rect 2158 3548 2162 3552
rect 2166 3548 2170 3552
rect 2190 3548 2194 3552
rect 62 3538 66 3542
rect 78 3538 82 3542
rect 222 3538 226 3542
rect 406 3538 410 3542
rect 486 3538 490 3542
rect 494 3538 498 3542
rect 558 3538 562 3542
rect 566 3538 570 3542
rect 630 3538 634 3542
rect 646 3538 650 3542
rect 758 3538 762 3542
rect 766 3538 770 3542
rect 782 3538 786 3542
rect 806 3538 810 3542
rect 894 3538 898 3542
rect 966 3538 970 3542
rect 1038 3538 1042 3542
rect 1062 3538 1066 3542
rect 1158 3538 1162 3542
rect 1198 3538 1202 3542
rect 1246 3538 1250 3542
rect 1270 3538 1274 3542
rect 1334 3538 1338 3542
rect 1406 3538 1410 3542
rect 1422 3538 1426 3542
rect 1534 3538 1538 3542
rect 1558 3538 1562 3542
rect 1862 3538 1866 3542
rect 1878 3538 1882 3542
rect 1910 3538 1914 3542
rect 1966 3538 1970 3542
rect 1974 3538 1978 3542
rect 2030 3538 2034 3542
rect 2086 3538 2090 3542
rect 2134 3538 2138 3542
rect 2262 3547 2266 3551
rect 2382 3547 2386 3551
rect 2446 3548 2450 3552
rect 2790 3548 2794 3552
rect 2846 3548 2850 3552
rect 2894 3548 2898 3552
rect 2942 3548 2946 3552
rect 2990 3548 2994 3552
rect 3150 3548 3154 3552
rect 3342 3548 3346 3552
rect 3374 3548 3378 3552
rect 3398 3548 3402 3552
rect 3494 3548 3498 3552
rect 2278 3538 2282 3542
rect 2310 3538 2314 3542
rect 2414 3538 2418 3542
rect 2486 3538 2490 3542
rect 2510 3538 2514 3542
rect 2550 3538 2554 3542
rect 2686 3538 2690 3542
rect 2790 3538 2794 3542
rect 3046 3538 3050 3542
rect 3110 3538 3114 3542
rect 3126 3538 3130 3542
rect 3134 3538 3138 3542
rect 3542 3547 3546 3551
rect 3574 3548 3578 3552
rect 3654 3547 3658 3551
rect 3686 3548 3690 3552
rect 3742 3548 3746 3552
rect 3798 3547 3802 3551
rect 3918 3547 3922 3551
rect 3950 3548 3954 3552
rect 4014 3547 4018 3551
rect 4126 3547 4130 3551
rect 4270 3547 4274 3551
rect 4366 3548 4370 3552
rect 4422 3547 4426 3551
rect 4566 3548 4570 3552
rect 4574 3548 4578 3552
rect 3174 3538 3178 3542
rect 3246 3538 3250 3542
rect 3286 3538 3290 3542
rect 3318 3538 3322 3542
rect 3390 3538 3394 3542
rect 3414 3538 3418 3542
rect 3422 3538 3426 3542
rect 3438 3538 3442 3542
rect 3806 3538 3810 3542
rect 3886 3538 3890 3542
rect 3998 3538 4002 3542
rect 4038 3538 4042 3542
rect 4110 3538 4114 3542
rect 4214 3538 4218 3542
rect 4254 3538 4258 3542
rect 4342 3538 4346 3542
rect 4350 3538 4354 3542
rect 4406 3538 4410 3542
rect 4494 3538 4498 3542
rect 4518 3538 4522 3542
rect 4566 3538 4570 3542
rect 6 3528 10 3532
rect 22 3528 26 3532
rect 86 3528 90 3532
rect 390 3528 394 3532
rect 406 3528 410 3532
rect 446 3528 450 3532
rect 494 3528 498 3532
rect 662 3528 666 3532
rect 1078 3528 1082 3532
rect 1382 3528 1386 3532
rect 1438 3528 1442 3532
rect 1646 3528 1650 3532
rect 1846 3528 1850 3532
rect 2046 3528 2050 3532
rect 2382 3528 2386 3532
rect 2422 3528 2426 3532
rect 2526 3528 2530 3532
rect 2558 3528 2562 3532
rect 2606 3528 2610 3532
rect 2654 3528 2658 3532
rect 2822 3528 2826 3532
rect 2878 3528 2882 3532
rect 2918 3528 2922 3532
rect 2966 3528 2970 3532
rect 3062 3528 3066 3532
rect 3094 3528 3098 3532
rect 3222 3528 3226 3532
rect 3254 3528 3258 3532
rect 3470 3528 3474 3532
rect 3510 3528 3514 3532
rect 3766 3528 3770 3532
rect 4334 3528 4338 3532
rect 46 3518 50 3522
rect 422 3518 426 3522
rect 534 3518 538 3522
rect 542 3518 546 3522
rect 726 3518 730 3522
rect 734 3518 738 3522
rect 1454 3518 1458 3522
rect 1638 3518 1642 3522
rect 1654 3518 1658 3522
rect 2302 3518 2306 3522
rect 2470 3518 2474 3522
rect 2590 3518 2594 3522
rect 2638 3518 2642 3522
rect 2694 3518 2698 3522
rect 2758 3518 2762 3522
rect 2774 3518 2778 3522
rect 2814 3518 2818 3522
rect 2910 3518 2914 3522
rect 3014 3518 3018 3522
rect 3110 3518 3114 3522
rect 3150 3518 3154 3522
rect 3198 3518 3202 3522
rect 3230 3518 3234 3522
rect 3286 3518 3290 3522
rect 3310 3518 3314 3522
rect 3334 3518 3338 3522
rect 3358 3518 3362 3522
rect 3462 3518 3466 3522
rect 3862 3518 3866 3522
rect 3870 3518 3874 3522
rect 3982 3518 3986 3522
rect 4094 3518 4098 3522
rect 4382 3518 4386 3522
rect 4486 3518 4490 3522
rect 4510 3518 4514 3522
rect 4590 3518 4594 3522
rect 3470 3508 3474 3512
rect 3766 3508 3770 3512
rect 1002 3503 1006 3507
rect 1009 3503 1013 3507
rect 2026 3503 2030 3507
rect 2033 3503 2037 3507
rect 3050 3503 3054 3507
rect 3057 3503 3061 3507
rect 4082 3503 4086 3507
rect 4089 3503 4093 3507
rect 3550 3498 3554 3502
rect 3750 3498 3754 3502
rect 3910 3498 3914 3502
rect 126 3488 130 3492
rect 190 3488 194 3492
rect 318 3488 322 3492
rect 382 3488 386 3492
rect 1022 3488 1026 3492
rect 1134 3488 1138 3492
rect 1510 3488 1514 3492
rect 1798 3488 1802 3492
rect 1910 3488 1914 3492
rect 1958 3488 1962 3492
rect 1974 3488 1978 3492
rect 2078 3488 2082 3492
rect 2174 3488 2178 3492
rect 2326 3488 2330 3492
rect 2414 3488 2418 3492
rect 2486 3488 2490 3492
rect 2582 3488 2586 3492
rect 3246 3488 3250 3492
rect 3382 3488 3386 3492
rect 3414 3488 3418 3492
rect 3430 3488 3434 3492
rect 3718 3488 3722 3492
rect 3806 3488 3810 3492
rect 4006 3488 4010 3492
rect 4182 3488 4186 3492
rect 4318 3488 4322 3492
rect 6 3478 10 3482
rect 70 3478 74 3482
rect 134 3478 138 3482
rect 230 3478 234 3482
rect 318 3478 322 3482
rect 382 3478 386 3482
rect 414 3478 418 3482
rect 470 3478 474 3482
rect 750 3478 754 3482
rect 830 3478 834 3482
rect 1414 3478 1418 3482
rect 1574 3478 1578 3482
rect 1894 3478 1898 3482
rect 2086 3478 2090 3482
rect 2134 3478 2138 3482
rect 2182 3478 2186 3482
rect 2198 3478 2202 3482
rect 2422 3478 2426 3482
rect 2526 3478 2530 3482
rect 2622 3478 2626 3482
rect 2862 3478 2866 3482
rect 2878 3478 2882 3482
rect 3038 3478 3042 3482
rect 3078 3478 3082 3482
rect 3510 3478 3514 3482
rect 3550 3478 3554 3482
rect 3750 3478 3754 3482
rect 3910 3478 3914 3482
rect 4038 3478 4042 3482
rect 22 3468 26 3472
rect 62 3468 66 3472
rect 126 3468 130 3472
rect 150 3468 154 3472
rect 286 3468 290 3472
rect 318 3468 322 3472
rect 422 3468 426 3472
rect 446 3468 450 3472
rect 526 3468 530 3472
rect 574 3468 578 3472
rect 662 3468 666 3472
rect 846 3468 850 3472
rect 942 3468 946 3472
rect 1078 3468 1082 3472
rect 1198 3468 1202 3472
rect 1246 3468 1250 3472
rect 1270 3468 1274 3472
rect 1334 3468 1338 3472
rect 1398 3468 1402 3472
rect 1430 3468 1434 3472
rect 1446 3468 1450 3472
rect 1494 3468 1498 3472
rect 1686 3468 1690 3472
rect 1782 3468 1786 3472
rect 1894 3468 1898 3472
rect 1934 3468 1938 3472
rect 1998 3468 2002 3472
rect 2038 3468 2042 3472
rect 2054 3468 2058 3472
rect 2150 3468 2154 3472
rect 2278 3468 2282 3472
rect 2294 3468 2298 3472
rect 2342 3468 2346 3472
rect 2398 3468 2402 3472
rect 2422 3468 2426 3472
rect 2438 3468 2442 3472
rect 2462 3468 2466 3472
rect 2718 3468 2722 3472
rect 3014 3468 3018 3472
rect 3054 3468 3058 3472
rect 3206 3468 3210 3472
rect 3262 3468 3266 3472
rect 3374 3468 3378 3472
rect 3398 3468 3402 3472
rect 3438 3468 3442 3472
rect 3446 3468 3450 3472
rect 3462 3468 3466 3472
rect 3518 3468 3522 3472
rect 3622 3468 3626 3472
rect 3662 3468 3666 3472
rect 3742 3468 3746 3472
rect 3862 3468 3866 3472
rect 3950 3468 3954 3472
rect 4110 3468 4114 3472
rect 4206 3468 4210 3472
rect 4286 3468 4290 3472
rect 4294 3468 4298 3472
rect 4326 3468 4330 3472
rect 4366 3468 4370 3472
rect 4382 3468 4386 3472
rect 4486 3468 4490 3472
rect 4502 3468 4506 3472
rect 4558 3468 4562 3472
rect 78 3458 82 3462
rect 118 3458 122 3462
rect 174 3458 178 3462
rect 214 3458 218 3462
rect 246 3458 250 3462
rect 310 3458 314 3462
rect 374 3458 378 3462
rect 510 3458 514 3462
rect 518 3458 522 3462
rect 558 3459 562 3463
rect 654 3459 658 3463
rect 750 3459 754 3463
rect 870 3458 874 3462
rect 894 3458 898 3462
rect 958 3459 962 3463
rect 1070 3459 1074 3463
rect 1206 3459 1210 3463
rect 1238 3458 1242 3462
rect 1254 3458 1258 3462
rect 1310 3458 1314 3462
rect 1342 3459 1346 3463
rect 1422 3458 1426 3462
rect 1438 3458 1442 3462
rect 1454 3458 1458 3462
rect 1478 3458 1482 3462
rect 1574 3459 1578 3463
rect 1670 3459 1674 3463
rect 1766 3459 1770 3463
rect 1830 3458 1834 3462
rect 1862 3459 1866 3463
rect 1926 3458 1930 3462
rect 1942 3458 1946 3462
rect 1990 3458 1994 3462
rect 1998 3458 2002 3462
rect 2030 3458 2034 3462
rect 2102 3458 2106 3462
rect 2150 3458 2154 3462
rect 2158 3458 2162 3462
rect 2222 3458 2226 3462
rect 2254 3458 2258 3462
rect 2310 3458 2314 3462
rect 2350 3458 2354 3462
rect 2374 3458 2378 3462
rect 2470 3458 2474 3462
rect 2502 3458 2506 3462
rect 2566 3458 2570 3462
rect 2606 3458 2610 3462
rect 2622 3458 2626 3462
rect 2654 3458 2658 3462
rect 2686 3458 2690 3462
rect 2710 3458 2714 3462
rect 2742 3458 2746 3462
rect 2782 3458 2786 3462
rect 2806 3458 2810 3462
rect 2822 3458 2826 3462
rect 2838 3458 2842 3462
rect 2902 3458 2906 3462
rect 2934 3458 2938 3462
rect 2966 3458 2970 3462
rect 2998 3458 3002 3462
rect 3038 3458 3042 3462
rect 3102 3458 3106 3462
rect 3134 3458 3138 3462
rect 3166 3458 3170 3462
rect 3222 3458 3226 3462
rect 3286 3458 3290 3462
rect 3326 3458 3330 3462
rect 3350 3458 3354 3462
rect 3486 3458 3490 3462
rect 3574 3458 3578 3462
rect 3598 3458 3602 3462
rect 3654 3459 3658 3463
rect 3686 3458 3690 3462
rect 3726 3458 3730 3462
rect 3774 3458 3778 3462
rect 3790 3458 3794 3462
rect 3886 3458 3890 3462
rect 3942 3459 3946 3463
rect 4038 3459 4042 3463
rect 4222 3459 4226 3463
rect 4302 3458 4306 3462
rect 4350 3458 4354 3462
rect 4390 3458 4394 3462
rect 4430 3458 4434 3462
rect 4454 3458 4458 3462
rect 4518 3458 4522 3462
rect 4566 3458 4570 3462
rect 438 3448 442 3452
rect 462 3448 466 3452
rect 486 3448 490 3452
rect 502 3448 506 3452
rect 1374 3448 1378 3452
rect 1462 3448 1466 3452
rect 2078 3448 2082 3452
rect 2094 3448 2098 3452
rect 2182 3448 2186 3452
rect 2190 3448 2194 3452
rect 2214 3448 2218 3452
rect 2238 3448 2242 3452
rect 2246 3448 2250 3452
rect 2286 3448 2290 3452
rect 2326 3448 2330 3452
rect 2358 3448 2362 3452
rect 2366 3448 2370 3452
rect 2414 3448 2418 3452
rect 2446 3448 2450 3452
rect 2486 3448 2490 3452
rect 2494 3448 2498 3452
rect 2526 3448 2530 3452
rect 2614 3448 2618 3452
rect 2662 3448 2666 3452
rect 2694 3448 2698 3452
rect 2702 3448 2706 3452
rect 2734 3448 2738 3452
rect 2790 3448 2794 3452
rect 2798 3448 2802 3452
rect 2830 3448 2834 3452
rect 2878 3448 2882 3452
rect 2894 3448 2898 3452
rect 2926 3448 2930 3452
rect 2958 3448 2962 3452
rect 2990 3448 2994 3452
rect 3046 3448 3050 3452
rect 3086 3448 3090 3452
rect 3094 3448 3098 3452
rect 3126 3448 3130 3452
rect 3158 3448 3162 3452
rect 3190 3448 3194 3452
rect 3214 3448 3218 3452
rect 3278 3448 3282 3452
rect 3334 3448 3338 3452
rect 3390 3448 3394 3452
rect 3414 3448 3418 3452
rect 3462 3448 3466 3452
rect 3598 3448 3602 3452
rect 3606 3448 3610 3452
rect 3742 3448 3746 3452
rect 3790 3448 3794 3452
rect 3870 3448 3874 3452
rect 3886 3448 3890 3452
rect 4318 3448 4322 3452
rect 4350 3448 4354 3452
rect 4366 3448 4370 3452
rect 4438 3448 4442 3452
rect 4502 3448 4506 3452
rect 4510 3448 4514 3452
rect 4542 3448 4546 3452
rect 446 3438 450 3442
rect 718 3438 722 3442
rect 830 3438 834 3442
rect 926 3438 930 3442
rect 1294 3438 1298 3442
rect 1910 3438 1914 3442
rect 1974 3438 1978 3442
rect 2230 3438 2234 3442
rect 2262 3438 2266 3442
rect 2342 3438 2346 3442
rect 2382 3438 2386 3442
rect 2510 3438 2514 3442
rect 2574 3438 2578 3442
rect 2598 3438 2602 3442
rect 2646 3438 2650 3442
rect 2686 3438 2690 3442
rect 2718 3438 2722 3442
rect 2750 3438 2754 3442
rect 2774 3438 2778 3442
rect 2814 3438 2818 3442
rect 2846 3438 2850 3442
rect 2910 3438 2914 3442
rect 2942 3438 2946 3442
rect 2966 3438 2970 3442
rect 2974 3438 2978 3442
rect 2998 3438 3002 3442
rect 3030 3438 3034 3442
rect 3110 3438 3114 3442
rect 3142 3438 3146 3442
rect 3174 3438 3178 3442
rect 3206 3438 3210 3442
rect 3230 3438 3234 3442
rect 3294 3438 3298 3442
rect 3318 3438 3322 3442
rect 3358 3438 3362 3442
rect 3518 3438 3522 3442
rect 3534 3438 3538 3442
rect 4526 3438 4530 3442
rect 4550 3438 4554 3442
rect 814 3428 818 3432
rect 30 3418 34 3422
rect 430 3418 434 3422
rect 622 3418 626 3422
rect 1142 3418 1146 3422
rect 1606 3418 1610 3422
rect 1702 3418 1706 3422
rect 2118 3418 2122 3422
rect 2206 3418 2210 3422
rect 2254 3418 2258 3422
rect 2374 3418 2378 3422
rect 2606 3418 2610 3422
rect 2654 3418 2658 3422
rect 2686 3418 2690 3422
rect 2758 3418 2762 3422
rect 2782 3418 2786 3422
rect 2838 3418 2842 3422
rect 2886 3418 2890 3422
rect 2902 3418 2906 3422
rect 2934 3418 2938 3422
rect 3102 3418 3106 3422
rect 3134 3418 3138 3422
rect 3166 3418 3170 3422
rect 3222 3418 3226 3422
rect 3286 3418 3290 3422
rect 3326 3418 3330 3422
rect 3350 3418 3354 3422
rect 3614 3418 3618 3422
rect 3806 3418 3810 3422
rect 4102 3418 4106 3422
rect 498 3403 502 3407
rect 505 3403 509 3407
rect 1522 3403 1526 3407
rect 1529 3403 1533 3407
rect 2546 3403 2550 3407
rect 2553 3403 2557 3407
rect 3570 3403 3574 3407
rect 3577 3403 3581 3407
rect 310 3388 314 3392
rect 1094 3388 1098 3392
rect 1494 3388 1498 3392
rect 1942 3388 1946 3392
rect 2166 3388 2170 3392
rect 2190 3388 2194 3392
rect 2238 3388 2242 3392
rect 2358 3388 2362 3392
rect 2486 3388 2490 3392
rect 2622 3388 2626 3392
rect 2662 3388 2666 3392
rect 2702 3388 2706 3392
rect 2742 3388 2746 3392
rect 2854 3388 2858 3392
rect 3046 3388 3050 3392
rect 4190 3388 4194 3392
rect 2118 3378 2122 3382
rect 3734 3378 3738 3382
rect 790 3368 794 3372
rect 1190 3368 1194 3372
rect 1910 3368 1914 3372
rect 1958 3368 1962 3372
rect 2518 3368 2522 3372
rect 2614 3368 2618 3372
rect 2750 3368 2754 3372
rect 2782 3368 2786 3372
rect 2846 3368 2850 3372
rect 2918 3368 2922 3372
rect 2998 3368 3002 3372
rect 3358 3368 3362 3372
rect 3478 3368 3482 3372
rect 3486 3368 3490 3372
rect 3502 3368 3506 3372
rect 38 3357 42 3361
rect 438 3358 442 3362
rect 558 3358 562 3362
rect 606 3358 610 3362
rect 654 3358 658 3362
rect 1222 3358 1226 3362
rect 1334 3358 1338 3362
rect 1638 3358 1642 3362
rect 1670 3358 1674 3362
rect 1806 3358 1810 3362
rect 1926 3358 1930 3362
rect 2054 3358 2058 3362
rect 2142 3358 2146 3362
rect 2150 3358 2154 3362
rect 2206 3358 2210 3362
rect 2254 3358 2258 3362
rect 2262 3358 2266 3362
rect 2366 3358 2370 3362
rect 2510 3358 2514 3362
rect 2550 3358 2554 3362
rect 2590 3358 2594 3362
rect 2598 3358 2602 3362
rect 2630 3358 2634 3362
rect 2646 3358 2650 3362
rect 2678 3358 2682 3362
rect 2774 3358 2778 3362
rect 2790 3358 2794 3362
rect 2830 3358 2834 3362
rect 2886 3358 2890 3362
rect 2926 3358 2930 3362
rect 2934 3358 2938 3362
rect 2966 3358 2970 3362
rect 2974 3358 2978 3362
rect 3006 3358 3010 3362
rect 3110 3358 3114 3362
rect 3118 3358 3122 3362
rect 3158 3358 3162 3362
rect 3166 3358 3170 3362
rect 3190 3358 3194 3362
rect 3214 3358 3218 3362
rect 3238 3358 3242 3362
rect 3286 3358 3290 3362
rect 3302 3358 3306 3362
rect 3310 3358 3314 3362
rect 3350 3358 3354 3362
rect 3398 3358 3402 3362
rect 3406 3358 3410 3362
rect 3742 3368 3746 3372
rect 3838 3368 3842 3372
rect 3526 3358 3530 3362
rect 3550 3358 3554 3362
rect 3638 3358 3642 3362
rect 3678 3358 3682 3362
rect 3886 3358 3890 3362
rect 4334 3358 4338 3362
rect 4502 3358 4506 3362
rect 4550 3358 4554 3362
rect 4590 3358 4594 3362
rect 62 3348 66 3352
rect 110 3347 114 3351
rect 206 3347 210 3351
rect 294 3348 298 3352
rect 366 3348 370 3352
rect 422 3348 426 3352
rect 470 3347 474 3351
rect 566 3348 570 3352
rect 726 3347 730 3351
rect 822 3347 826 3351
rect 846 3348 850 3352
rect 926 3348 930 3352
rect 942 3348 946 3352
rect 1030 3347 1034 3351
rect 1134 3348 1138 3352
rect 1198 3348 1202 3352
rect 1230 3348 1234 3352
rect 1262 3347 1266 3351
rect 1294 3348 1298 3352
rect 1414 3348 1418 3352
rect 1446 3347 1450 3351
rect 1478 3348 1482 3352
rect 1526 3348 1530 3352
rect 1542 3348 1546 3352
rect 1558 3348 1562 3352
rect 1566 3348 1570 3352
rect 1582 3348 1586 3352
rect 1606 3348 1610 3352
rect 1630 3348 1634 3352
rect 1662 3348 1666 3352
rect 1694 3348 1698 3352
rect 1734 3348 1738 3352
rect 1766 3347 1770 3351
rect 1846 3348 1850 3352
rect 1878 3347 1882 3351
rect 1950 3348 1954 3352
rect 1990 3348 1994 3352
rect 2022 3347 2026 3351
rect 2078 3348 2082 3352
rect 2086 3348 2090 3352
rect 2102 3348 2106 3352
rect 2118 3348 2122 3352
rect 2166 3348 2170 3352
rect 2190 3348 2194 3352
rect 2310 3348 2314 3352
rect 2342 3348 2346 3352
rect 2510 3348 2514 3352
rect 2606 3348 2610 3352
rect 2742 3348 2746 3352
rect 2854 3348 2858 3352
rect 2990 3348 2994 3352
rect 3062 3348 3066 3352
rect 3270 3348 3274 3352
rect 3326 3348 3330 3352
rect 3454 3348 3458 3352
rect 3462 3348 3466 3352
rect 3622 3348 3626 3352
rect 3646 3348 3650 3352
rect 3670 3348 3674 3352
rect 3694 3348 3698 3352
rect 22 3338 26 3342
rect 62 3338 66 3342
rect 190 3338 194 3342
rect 334 3338 338 3342
rect 374 3338 378 3342
rect 414 3338 418 3342
rect 486 3338 490 3342
rect 582 3338 586 3342
rect 630 3338 634 3342
rect 678 3338 682 3342
rect 710 3338 714 3342
rect 854 3338 858 3342
rect 1014 3338 1018 3342
rect 1062 3338 1066 3342
rect 1110 3338 1114 3342
rect 1206 3338 1210 3342
rect 1222 3338 1226 3342
rect 1358 3338 1362 3342
rect 1502 3338 1506 3342
rect 1550 3338 1554 3342
rect 1574 3338 1578 3342
rect 1590 3338 1594 3342
rect 1662 3338 1666 3342
rect 1694 3338 1698 3342
rect 1782 3338 1786 3342
rect 1894 3338 1898 3342
rect 1950 3338 1954 3342
rect 2094 3338 2098 3342
rect 2126 3338 2130 3342
rect 2174 3338 2178 3342
rect 2182 3338 2186 3342
rect 2230 3338 2234 3342
rect 2278 3338 2282 3342
rect 2286 3338 2290 3342
rect 2318 3338 2322 3342
rect 2382 3338 2386 3342
rect 2390 3338 2394 3342
rect 2454 3338 2458 3342
rect 2478 3338 2482 3342
rect 2526 3338 2530 3342
rect 2534 3338 2538 3342
rect 2574 3338 2578 3342
rect 2654 3338 2658 3342
rect 2678 3338 2682 3342
rect 2694 3338 2698 3342
rect 2766 3338 2770 3342
rect 2806 3338 2810 3342
rect 2814 3338 2818 3342
rect 2902 3338 2906 3342
rect 2910 3338 2914 3342
rect 2950 3338 2954 3342
rect 2958 3338 2962 3342
rect 2974 3338 2978 3342
rect 3030 3338 3034 3342
rect 3086 3338 3090 3342
rect 3094 3338 3098 3342
rect 3134 3338 3138 3342
rect 3142 3338 3146 3342
rect 3182 3338 3186 3342
rect 3230 3338 3234 3342
rect 3254 3338 3258 3342
rect 3262 3338 3266 3342
rect 3286 3338 3290 3342
rect 3326 3338 3330 3342
rect 3374 3338 3378 3342
rect 3382 3338 3386 3342
rect 3422 3338 3426 3342
rect 3430 3338 3434 3342
rect 3478 3338 3482 3342
rect 3502 3338 3506 3342
rect 3526 3338 3530 3342
rect 3550 3338 3554 3342
rect 3574 3338 3578 3342
rect 3774 3347 3778 3351
rect 3806 3348 3810 3352
rect 3862 3348 3866 3352
rect 3918 3347 3922 3351
rect 4022 3348 4026 3352
rect 4126 3347 4130 3351
rect 4222 3347 4226 3351
rect 4294 3348 4298 3352
rect 4310 3348 4314 3352
rect 4326 3348 4330 3352
rect 4350 3348 4354 3352
rect 4390 3347 4394 3351
rect 4454 3348 4458 3352
rect 4478 3348 4482 3352
rect 4526 3348 4530 3352
rect 3686 3338 3690 3342
rect 3726 3338 3730 3342
rect 3830 3338 3834 3342
rect 3886 3338 3890 3342
rect 3902 3338 3906 3342
rect 3934 3338 3938 3342
rect 4030 3338 4034 3342
rect 4070 3338 4074 3342
rect 4230 3338 4234 3342
rect 4302 3338 4306 3342
rect 4318 3338 4322 3342
rect 4358 3338 4362 3342
rect 4406 3338 4410 3342
rect 4414 3338 4418 3342
rect 4486 3338 4490 3342
rect 4534 3338 4538 3342
rect 4558 3338 4562 3342
rect 6 3328 10 3332
rect 70 3328 74 3332
rect 110 3328 114 3332
rect 254 3328 258 3332
rect 302 3328 306 3332
rect 318 3328 322 3332
rect 382 3328 386 3332
rect 398 3328 402 3332
rect 598 3328 602 3332
rect 646 3328 650 3332
rect 694 3328 698 3332
rect 1918 3328 1922 3332
rect 2134 3328 2138 3332
rect 2214 3328 2218 3332
rect 2350 3328 2354 3332
rect 2462 3328 2466 3332
rect 2686 3328 2690 3332
rect 2710 3328 2714 3332
rect 2878 3328 2882 3332
rect 3030 3328 3034 3332
rect 3126 3328 3130 3332
rect 3198 3328 3202 3332
rect 3246 3328 3250 3332
rect 3318 3328 3322 3332
rect 3598 3328 3602 3332
rect 3718 3328 3722 3332
rect 3846 3328 3850 3332
rect 4126 3328 4130 3332
rect 4270 3328 4274 3332
rect 174 3318 178 3322
rect 270 3318 274 3322
rect 374 3318 378 3322
rect 438 3318 442 3322
rect 534 3318 538 3322
rect 606 3318 610 3322
rect 654 3318 658 3322
rect 886 3318 890 3322
rect 982 3318 986 3322
rect 1326 3318 1330 3322
rect 1494 3318 1498 3322
rect 1702 3318 1706 3322
rect 2262 3318 2266 3322
rect 2366 3318 2370 3322
rect 2550 3318 2554 3322
rect 2590 3318 2594 3322
rect 2630 3318 2634 3322
rect 2790 3318 2794 3322
rect 2830 3318 2834 3322
rect 2886 3318 2890 3322
rect 2934 3318 2938 3322
rect 3006 3318 3010 3322
rect 3110 3318 3114 3322
rect 3158 3318 3162 3322
rect 3166 3318 3170 3322
rect 3302 3318 3306 3322
rect 3350 3318 3354 3322
rect 3358 3318 3362 3322
rect 3398 3318 3402 3322
rect 3406 3318 3410 3322
rect 3494 3318 3498 3322
rect 3518 3318 3522 3322
rect 3542 3318 3546 3322
rect 3558 3318 3562 3322
rect 3638 3318 3642 3322
rect 3982 3318 3986 3322
rect 4494 3318 4498 3322
rect 4542 3318 4546 3322
rect 4566 3318 4570 3322
rect 3718 3308 3722 3312
rect 3846 3308 3850 3312
rect 1002 3303 1006 3307
rect 1009 3303 1013 3307
rect 2026 3303 2030 3307
rect 2033 3303 2037 3307
rect 3050 3303 3054 3307
rect 3057 3303 3061 3307
rect 4082 3303 4086 3307
rect 4089 3303 4093 3307
rect 3438 3298 3442 3302
rect 3598 3298 3602 3302
rect 3742 3298 3746 3302
rect 294 3288 298 3292
rect 430 3288 434 3292
rect 1030 3288 1034 3292
rect 1126 3288 1130 3292
rect 1222 3288 1226 3292
rect 1518 3288 1522 3292
rect 1822 3288 1826 3292
rect 2030 3288 2034 3292
rect 2126 3288 2130 3292
rect 2246 3288 2250 3292
rect 2278 3288 2282 3292
rect 2286 3288 2290 3292
rect 2390 3288 2394 3292
rect 2462 3288 2466 3292
rect 2502 3288 2506 3292
rect 2526 3288 2530 3292
rect 2534 3288 2538 3292
rect 2630 3288 2634 3292
rect 2654 3288 2658 3292
rect 2678 3288 2682 3292
rect 2702 3288 2706 3292
rect 2766 3288 2770 3292
rect 2814 3288 2818 3292
rect 2846 3288 2850 3292
rect 2854 3288 2858 3292
rect 2894 3288 2898 3292
rect 2910 3288 2914 3292
rect 2926 3288 2930 3292
rect 2950 3288 2954 3292
rect 3006 3288 3010 3292
rect 3030 3288 3034 3292
rect 3038 3288 3042 3292
rect 3126 3288 3130 3292
rect 3134 3288 3138 3292
rect 3230 3288 3234 3292
rect 3254 3288 3258 3292
rect 3286 3288 3290 3292
rect 3310 3288 3314 3292
rect 3334 3288 3338 3292
rect 4206 3288 4210 3292
rect 4494 3288 4498 3292
rect 4510 3288 4514 3292
rect 230 3278 234 3282
rect 246 3278 250 3282
rect 262 3278 266 3282
rect 334 3278 338 3282
rect 462 3278 466 3282
rect 470 3278 474 3282
rect 518 3278 522 3282
rect 726 3278 730 3282
rect 774 3278 778 3282
rect 854 3278 858 3282
rect 1062 3278 1066 3282
rect 1422 3278 1426 3282
rect 110 3268 114 3272
rect 230 3268 234 3272
rect 254 3268 258 3272
rect 286 3268 290 3272
rect 302 3268 306 3272
rect 334 3268 338 3272
rect 342 3268 346 3272
rect 382 3268 386 3272
rect 398 3268 402 3272
rect 1486 3278 1490 3282
rect 2062 3278 2066 3282
rect 2094 3278 2098 3282
rect 2190 3278 2194 3282
rect 2558 3278 2562 3282
rect 2974 3278 2978 3282
rect 3222 3278 3226 3282
rect 3390 3278 3394 3282
rect 3438 3278 3442 3282
rect 3598 3278 3602 3282
rect 3702 3278 3706 3282
rect 3742 3278 3746 3282
rect 3862 3278 3866 3282
rect 542 3268 546 3272
rect 806 3268 810 3272
rect 822 3268 826 3272
rect 1238 3268 1242 3272
rect 1334 3268 1338 3272
rect 1438 3268 1442 3272
rect 1478 3268 1482 3272
rect 1502 3268 1506 3272
rect 1806 3268 1810 3272
rect 1902 3268 1906 3272
rect 1918 3268 1922 3272
rect 1934 3268 1938 3272
rect 4014 3278 4018 3282
rect 4366 3278 4370 3282
rect 4534 3278 4538 3282
rect 2222 3268 2226 3272
rect 2254 3268 2258 3272
rect 2342 3268 2346 3272
rect 2398 3268 2402 3272
rect 2406 3268 2410 3272
rect 2430 3268 2434 3272
rect 2478 3268 2482 3272
rect 2502 3268 2506 3272
rect 2558 3268 2562 3272
rect 38 3258 42 3262
rect 62 3258 66 3262
rect 126 3259 130 3263
rect 214 3258 218 3262
rect 278 3258 282 3262
rect 310 3258 314 3262
rect 342 3258 346 3262
rect 358 3258 362 3262
rect 366 3258 370 3262
rect 414 3258 418 3262
rect 446 3258 450 3262
rect 558 3259 562 3263
rect 582 3258 586 3262
rect 654 3259 658 3263
rect 678 3258 682 3262
rect 750 3258 754 3262
rect 790 3258 794 3262
rect 814 3258 818 3262
rect 854 3259 858 3263
rect 958 3258 962 3262
rect 982 3258 986 3262
rect 1062 3259 1066 3263
rect 1158 3259 1162 3263
rect 1190 3258 1194 3262
rect 1262 3258 1266 3262
rect 1366 3258 1370 3262
rect 1446 3258 1450 3262
rect 1462 3258 1466 3262
rect 1550 3258 1554 3262
rect 1582 3259 1586 3263
rect 1646 3258 1650 3262
rect 1678 3259 1682 3263
rect 1790 3259 1794 3263
rect 1886 3259 1890 3263
rect 1926 3258 1930 3262
rect 1982 3258 1986 3262
rect 2014 3258 2018 3262
rect 2094 3259 2098 3263
rect 2190 3259 2194 3263
rect 2230 3258 2234 3262
rect 2262 3258 2266 3262
rect 2350 3259 2354 3263
rect 2622 3268 2626 3272
rect 2646 3268 2650 3272
rect 2670 3268 2674 3272
rect 2710 3268 2714 3272
rect 2750 3268 2754 3272
rect 2766 3268 2770 3272
rect 2806 3268 2810 3272
rect 2830 3268 2834 3272
rect 2870 3268 2874 3272
rect 2878 3268 2882 3272
rect 2918 3268 2922 3272
rect 2942 3268 2946 3272
rect 2966 3268 2970 3272
rect 2990 3268 2994 3272
rect 3014 3268 3018 3272
rect 3054 3268 3058 3272
rect 3078 3268 3082 3272
rect 3094 3268 3098 3272
rect 3150 3268 3154 3272
rect 3158 3268 3162 3272
rect 3174 3268 3178 3272
rect 3246 3268 3250 3272
rect 3278 3268 3282 3272
rect 3302 3268 3306 3272
rect 3342 3268 3346 3272
rect 3526 3268 3530 3272
rect 3662 3268 3666 3272
rect 3766 3268 3770 3272
rect 3806 3268 3810 3272
rect 3902 3268 3906 3272
rect 3982 3268 3986 3272
rect 4030 3268 4034 3272
rect 4102 3268 4106 3272
rect 4110 3268 4114 3272
rect 4126 3268 4130 3272
rect 4214 3268 4218 3272
rect 4246 3268 4250 3272
rect 4278 3268 4282 3272
rect 4414 3268 4418 3272
rect 2438 3258 2442 3262
rect 2462 3258 2466 3262
rect 2598 3258 2602 3262
rect 2614 3258 2618 3262
rect 2718 3258 2722 3262
rect 2742 3258 2746 3262
rect 2798 3258 2802 3262
rect 3086 3258 3090 3262
rect 3198 3258 3202 3262
rect 3366 3258 3370 3262
rect 3406 3258 3410 3262
rect 3422 3258 3426 3262
rect 3502 3258 3506 3262
rect 3566 3258 3570 3262
rect 3670 3259 3674 3263
rect 3718 3258 3722 3262
rect 3798 3259 3802 3263
rect 3894 3259 3898 3263
rect 4014 3258 4018 3262
rect 4142 3259 4146 3263
rect 4222 3258 4226 3262
rect 4254 3258 4258 3262
rect 4342 3258 4346 3262
rect 4366 3258 4370 3262
rect 4430 3259 4434 3263
rect 4526 3258 4530 3262
rect 4550 3258 4554 3262
rect 238 3248 242 3252
rect 286 3248 290 3252
rect 374 3248 378 3252
rect 422 3248 426 3252
rect 798 3248 802 3252
rect 1422 3248 1426 3252
rect 1462 3248 1466 3252
rect 1950 3248 1954 3252
rect 2278 3248 2282 3252
rect 2382 3248 2386 3252
rect 2454 3248 2458 3252
rect 2462 3248 2466 3252
rect 2502 3248 2506 3252
rect 2534 3248 2538 3252
rect 2614 3248 2618 3252
rect 2638 3248 2642 3252
rect 2662 3248 2666 3252
rect 2686 3248 2690 3252
rect 2694 3248 2698 3252
rect 2766 3248 2770 3252
rect 2822 3248 2826 3252
rect 2846 3248 2850 3252
rect 2854 3248 2858 3252
rect 2894 3248 2898 3252
rect 2926 3248 2930 3252
rect 2950 3248 2954 3252
rect 2990 3248 2994 3252
rect 3006 3248 3010 3252
rect 3030 3248 3034 3252
rect 3038 3248 3042 3252
rect 3110 3248 3114 3252
rect 3126 3248 3130 3252
rect 3134 3248 3138 3252
rect 3174 3248 3178 3252
rect 3230 3248 3234 3252
rect 3254 3248 3258 3252
rect 3294 3248 3298 3252
rect 3318 3248 3322 3252
rect 3350 3248 3354 3252
rect 3398 3248 3402 3252
rect 3542 3248 3546 3252
rect 3702 3248 3706 3252
rect 3750 3248 3754 3252
rect 4006 3248 4010 3252
rect 4238 3248 4242 3252
rect 4254 3248 4258 3252
rect 4270 3248 4274 3252
rect 4302 3248 4306 3252
rect 4574 3248 4578 3252
rect 622 3238 626 3242
rect 718 3238 722 3242
rect 758 3238 762 3242
rect 1718 3238 1722 3242
rect 2246 3238 2250 3242
rect 2406 3238 2410 3242
rect 3606 3238 3610 3242
rect 3942 3238 3946 3242
rect 4190 3238 4194 3242
rect 782 3228 786 3232
rect 94 3218 98 3222
rect 190 3218 194 3222
rect 406 3218 410 3222
rect 494 3218 498 3222
rect 526 3218 530 3222
rect 766 3218 770 3222
rect 918 3218 922 3222
rect 1318 3218 1322 3222
rect 1414 3218 1418 3222
rect 1614 3218 1618 3222
rect 1990 3218 1994 3222
rect 3446 3218 3450 3222
rect 3558 3218 3562 3222
rect 3758 3218 3762 3222
rect 498 3203 502 3207
rect 505 3203 509 3207
rect 1522 3203 1526 3207
rect 1529 3203 1533 3207
rect 2546 3203 2550 3207
rect 2553 3203 2557 3207
rect 3570 3203 3574 3207
rect 3577 3203 3581 3207
rect 38 3188 42 3192
rect 86 3188 90 3192
rect 206 3188 210 3192
rect 294 3188 298 3192
rect 302 3188 306 3192
rect 366 3188 370 3192
rect 382 3188 386 3192
rect 1014 3188 1018 3192
rect 1102 3188 1106 3192
rect 1118 3188 1122 3192
rect 1358 3188 1362 3192
rect 1950 3188 1954 3192
rect 2166 3188 2170 3192
rect 2214 3188 2218 3192
rect 2310 3188 2314 3192
rect 2366 3188 2370 3192
rect 2710 3188 2714 3192
rect 2822 3188 2826 3192
rect 2902 3188 2906 3192
rect 3006 3188 3010 3192
rect 3214 3188 3218 3192
rect 3518 3188 3522 3192
rect 3766 3188 3770 3192
rect 238 3178 242 3182
rect 1550 3178 1554 3182
rect 4070 3178 4074 3182
rect 4406 3178 4410 3182
rect 30 3168 34 3172
rect 78 3168 82 3172
rect 198 3168 202 3172
rect 230 3168 234 3172
rect 286 3168 290 3172
rect 342 3168 346 3172
rect 358 3168 362 3172
rect 1630 3168 1634 3172
rect 1846 3168 1850 3172
rect 2078 3168 2082 3172
rect 46 3158 50 3162
rect 94 3158 98 3162
rect 3278 3168 3282 3172
rect 3646 3168 3650 3172
rect 3950 3168 3954 3172
rect 4438 3168 4442 3172
rect 214 3158 218 3162
rect 246 3158 250 3162
rect 270 3158 274 3162
rect 374 3158 378 3162
rect 446 3158 450 3162
rect 1334 3158 1338 3162
rect 1414 3158 1418 3162
rect 1662 3158 1666 3162
rect 1694 3158 1698 3162
rect 2078 3158 2082 3162
rect 6 3148 10 3152
rect 38 3148 42 3152
rect 54 3148 58 3152
rect 86 3148 90 3152
rect 150 3148 154 3152
rect 238 3148 242 3152
rect 278 3148 282 3152
rect 302 3148 306 3152
rect 342 3148 346 3152
rect 366 3148 370 3152
rect 382 3148 386 3152
rect 406 3148 410 3152
rect 422 3148 426 3152
rect 510 3148 514 3152
rect 526 3148 530 3152
rect 566 3148 570 3152
rect 598 3147 602 3151
rect 694 3147 698 3151
rect 790 3147 794 3151
rect 894 3148 898 3152
rect 1150 3148 1154 3152
rect 1166 3148 1170 3152
rect 1246 3148 1250 3152
rect 1310 3148 1314 3152
rect 118 3138 122 3142
rect 158 3138 162 3142
rect 198 3138 202 3142
rect 262 3138 266 3142
rect 430 3138 434 3142
rect 486 3138 490 3142
rect 494 3138 498 3142
rect 518 3138 522 3142
rect 534 3138 538 3142
rect 550 3138 554 3142
rect 582 3138 586 3142
rect 678 3138 682 3142
rect 902 3138 906 3142
rect 958 3138 962 3142
rect 1030 3138 1034 3142
rect 1318 3138 1322 3142
rect 1334 3138 1338 3142
rect 1374 3148 1378 3152
rect 1406 3148 1410 3152
rect 1438 3148 1442 3152
rect 1478 3148 1482 3152
rect 1526 3148 1530 3152
rect 1574 3148 1578 3152
rect 1582 3148 1586 3152
rect 1598 3148 1602 3152
rect 1614 3148 1618 3152
rect 1622 3148 1626 3152
rect 1662 3148 1666 3152
rect 1686 3148 1690 3152
rect 1718 3148 1722 3152
rect 1734 3148 1738 3152
rect 1774 3148 1778 3152
rect 1806 3147 1810 3151
rect 1918 3147 1922 3151
rect 2014 3147 2018 3151
rect 2094 3148 2098 3152
rect 2110 3148 2114 3152
rect 2126 3158 2130 3162
rect 2182 3158 2186 3162
rect 2230 3158 2234 3162
rect 2238 3158 2242 3162
rect 2254 3158 2258 3162
rect 2270 3158 2274 3162
rect 2342 3158 2346 3162
rect 2142 3148 2146 3152
rect 2166 3148 2170 3152
rect 2254 3148 2258 3152
rect 2278 3148 2282 3152
rect 2286 3148 2290 3152
rect 2318 3148 2322 3152
rect 2406 3158 2410 3162
rect 2414 3158 2418 3162
rect 2438 3158 2442 3162
rect 2462 3158 2466 3162
rect 2486 3158 2490 3162
rect 2510 3158 2514 3162
rect 2534 3158 2538 3162
rect 2606 3158 2610 3162
rect 2622 3158 2626 3162
rect 2630 3158 2634 3162
rect 2654 3158 2658 3162
rect 2662 3158 2666 3162
rect 2678 3158 2682 3162
rect 2734 3158 2738 3162
rect 2774 3158 2778 3162
rect 2782 3158 2786 3162
rect 2838 3158 2842 3162
rect 2862 3158 2866 3162
rect 2918 3158 2922 3162
rect 2934 3158 2938 3162
rect 2966 3158 2970 3162
rect 3022 3158 3026 3162
rect 3070 3158 3074 3162
rect 3102 3158 3106 3162
rect 3110 3158 3114 3162
rect 3150 3158 3154 3162
rect 3158 3158 3162 3162
rect 3182 3158 3186 3162
rect 3238 3158 3242 3162
rect 3254 3158 3258 3162
rect 3326 3158 3330 3162
rect 2366 3148 2370 3152
rect 2390 3148 2394 3152
rect 2398 3148 2402 3152
rect 2598 3148 2602 3152
rect 2726 3148 2730 3152
rect 2806 3148 2810 3152
rect 2886 3148 2890 3152
rect 2990 3148 2994 3152
rect 3230 3148 3234 3152
rect 3358 3158 3362 3162
rect 3670 3158 3674 3162
rect 3686 3158 3690 3162
rect 3758 3158 3762 3162
rect 4262 3158 4266 3162
rect 4294 3158 4298 3162
rect 4414 3158 4418 3162
rect 4422 3158 4426 3162
rect 4478 3158 4482 3162
rect 4558 3158 4562 3162
rect 4590 3158 4594 3162
rect 3374 3148 3378 3152
rect 1438 3138 1442 3142
rect 1534 3138 1538 3142
rect 1550 3138 1554 3142
rect 1566 3138 1570 3142
rect 1582 3138 1586 3142
rect 1606 3138 1610 3142
rect 1614 3138 1618 3142
rect 1646 3138 1650 3142
rect 1686 3138 1690 3142
rect 1718 3138 1722 3142
rect 2094 3138 2098 3142
rect 2150 3138 2154 3142
rect 2158 3138 2162 3142
rect 2206 3138 2210 3142
rect 2262 3138 2266 3142
rect 2294 3138 2298 3142
rect 2318 3138 2322 3142
rect 2374 3138 2378 3142
rect 2430 3138 2434 3142
rect 2454 3138 2458 3142
rect 2478 3138 2482 3142
rect 2502 3138 2506 3142
rect 2526 3138 2530 3142
rect 2550 3138 2554 3142
rect 2574 3138 2578 3142
rect 2622 3138 2626 3142
rect 2646 3138 2650 3142
rect 2670 3138 2674 3142
rect 2678 3138 2682 3142
rect 2694 3138 2698 3142
rect 2750 3138 2754 3142
rect 2758 3138 2762 3142
rect 2798 3138 2802 3142
rect 2862 3138 2866 3142
rect 2878 3138 2882 3142
rect 2934 3138 2938 3142
rect 2982 3138 2986 3142
rect 3038 3138 3042 3142
rect 3046 3138 3050 3142
rect 3086 3138 3090 3142
rect 3126 3138 3130 3142
rect 3430 3147 3434 3151
rect 3502 3148 3506 3152
rect 3574 3147 3578 3151
rect 3686 3148 3690 3152
rect 3742 3148 3746 3152
rect 3758 3148 3762 3152
rect 3822 3148 3826 3152
rect 3886 3147 3890 3151
rect 3918 3148 3922 3152
rect 3982 3147 3986 3151
rect 4014 3148 4018 3152
rect 4070 3148 4074 3152
rect 4198 3147 4202 3151
rect 4230 3148 4234 3152
rect 4278 3148 4282 3152
rect 4294 3148 4298 3152
rect 3174 3138 3178 3142
rect 3198 3138 3202 3142
rect 3254 3138 3258 3142
rect 3286 3138 3290 3142
rect 3302 3138 3306 3142
rect 3310 3138 3314 3142
rect 3350 3138 3354 3142
rect 3366 3138 3370 3142
rect 3414 3138 3418 3142
rect 3582 3138 3586 3142
rect 3662 3138 3666 3142
rect 3966 3138 3970 3142
rect 4046 3138 4050 3142
rect 4078 3138 4082 3142
rect 4102 3138 4106 3142
rect 4270 3138 4274 3142
rect 4326 3147 4330 3151
rect 4358 3148 4362 3152
rect 4430 3148 4434 3152
rect 4462 3148 4466 3152
rect 4486 3148 4490 3152
rect 4510 3148 4514 3152
rect 4534 3148 4538 3152
rect 4454 3138 4458 3142
rect 4566 3138 4570 3142
rect 6 3128 10 3132
rect 54 3128 58 3132
rect 102 3128 106 3132
rect 174 3128 178 3132
rect 182 3128 186 3132
rect 254 3128 258 3132
rect 318 3128 322 3132
rect 326 3128 330 3132
rect 398 3128 402 3132
rect 422 3128 426 3132
rect 454 3128 458 3132
rect 542 3128 546 3132
rect 790 3128 794 3132
rect 1238 3128 1242 3132
rect 1510 3128 1514 3132
rect 1918 3128 1922 3132
rect 2014 3128 2018 3132
rect 2062 3128 2066 3132
rect 2078 3128 2082 3132
rect 2190 3128 2194 3132
rect 2302 3128 2306 3132
rect 2614 3128 2618 3132
rect 2846 3128 2850 3132
rect 2870 3128 2874 3132
rect 2926 3128 2930 3132
rect 2950 3128 2954 3132
rect 3030 3128 3034 3132
rect 3142 3128 3146 3132
rect 3166 3128 3170 3132
rect 3190 3128 3194 3132
rect 3398 3128 3402 3132
rect 3710 3128 3714 3132
rect 3718 3128 3722 3132
rect 158 3118 162 3122
rect 662 3118 666 3122
rect 758 3118 762 3122
rect 854 3118 858 3122
rect 950 3118 954 3122
rect 1302 3118 1306 3122
rect 1390 3118 1394 3122
rect 1494 3118 1498 3122
rect 2414 3118 2418 3122
rect 2438 3118 2442 3122
rect 2462 3118 2466 3122
rect 2486 3118 2490 3122
rect 2510 3118 2514 3122
rect 2534 3118 2538 3122
rect 2582 3118 2586 3122
rect 2710 3118 2714 3122
rect 2734 3118 2738 3122
rect 2774 3118 2778 3122
rect 2782 3118 2786 3122
rect 3070 3118 3074 3122
rect 3102 3118 3106 3122
rect 3214 3118 3218 3122
rect 3238 3118 3242 3122
rect 3270 3118 3274 3122
rect 3294 3118 3298 3122
rect 3334 3118 3338 3122
rect 3494 3118 3498 3122
rect 3518 3118 3522 3122
rect 3638 3118 3642 3122
rect 3654 3118 3658 3122
rect 4158 3118 4162 3122
rect 4390 3118 4394 3122
rect 4558 3118 4562 3122
rect 4574 3118 4578 3122
rect 3398 3108 3402 3112
rect 3710 3108 3714 3112
rect 3718 3108 3722 3112
rect 1002 3103 1006 3107
rect 1009 3103 1013 3107
rect 2026 3103 2030 3107
rect 2033 3103 2037 3107
rect 3050 3103 3054 3107
rect 3057 3103 3061 3107
rect 4082 3103 4086 3107
rect 4089 3103 4093 3107
rect 3286 3098 3290 3102
rect 3454 3098 3458 3102
rect 3566 3098 3570 3102
rect 142 3088 146 3092
rect 238 3088 242 3092
rect 270 3088 274 3092
rect 350 3088 354 3092
rect 366 3088 370 3092
rect 438 3088 442 3092
rect 510 3088 514 3092
rect 526 3088 530 3092
rect 630 3088 634 3092
rect 894 3088 898 3092
rect 1102 3088 1106 3092
rect 1198 3088 1202 3092
rect 1294 3088 1298 3092
rect 1598 3088 1602 3092
rect 1694 3088 1698 3092
rect 1790 3088 1794 3092
rect 1886 3088 1890 3092
rect 1982 3088 1986 3092
rect 2126 3088 2130 3092
rect 2158 3088 2162 3092
rect 2222 3088 2226 3092
rect 2278 3088 2282 3092
rect 2342 3088 2346 3092
rect 2406 3088 2410 3092
rect 2494 3088 2498 3092
rect 2598 3088 2602 3092
rect 2630 3088 2634 3092
rect 2670 3088 2674 3092
rect 2718 3088 2722 3092
rect 2758 3088 2762 3092
rect 2774 3088 2778 3092
rect 2838 3088 2842 3092
rect 2862 3088 2866 3092
rect 2894 3088 2898 3092
rect 2934 3088 2938 3092
rect 2974 3088 2978 3092
rect 3014 3088 3018 3092
rect 3030 3088 3034 3092
rect 3094 3088 3098 3092
rect 3174 3088 3178 3092
rect 3198 3088 3202 3092
rect 3222 3088 3226 3092
rect 3246 3088 3250 3092
rect 3814 3088 3818 3092
rect 4110 3088 4114 3092
rect 4406 3088 4410 3092
rect 4446 3088 4450 3092
rect 38 3078 42 3082
rect 6 3068 10 3072
rect 326 3078 330 3082
rect 390 3078 394 3082
rect 430 3078 434 3082
rect 470 3078 474 3082
rect 662 3078 666 3082
rect 686 3078 690 3082
rect 774 3078 778 3082
rect 62 3068 66 3072
rect 190 3068 194 3072
rect 246 3068 250 3072
rect 262 3068 266 3072
rect 334 3068 338 3072
rect 1518 3078 1522 3082
rect 1726 3078 1730 3082
rect 2414 3078 2418 3082
rect 2510 3078 2514 3082
rect 2814 3078 2818 3082
rect 2846 3078 2850 3082
rect 2854 3078 2858 3082
rect 3286 3078 3290 3082
rect 3454 3078 3458 3082
rect 3566 3078 3570 3082
rect 4206 3078 4210 3082
rect 4278 3078 4282 3082
rect 4486 3078 4490 3082
rect 582 3068 586 3072
rect 630 3068 634 3072
rect 646 3068 650 3072
rect 702 3068 706 3072
rect 726 3068 730 3072
rect 758 3068 762 3072
rect 774 3068 778 3072
rect 798 3068 802 3072
rect 910 3068 914 3072
rect 1022 3068 1026 3072
rect 1150 3068 1154 3072
rect 1238 3068 1242 3072
rect 1310 3068 1314 3072
rect 1326 3068 1330 3072
rect 1350 3068 1354 3072
rect 1382 3068 1386 3072
rect 1398 3068 1402 3072
rect 1438 3068 1442 3072
rect 1454 3068 1458 3072
rect 1486 3068 1490 3072
rect 1502 3068 1506 3072
rect 1550 3068 1554 3072
rect 1590 3068 1594 3072
rect 1678 3068 1682 3072
rect 1774 3068 1778 3072
rect 1870 3068 1874 3072
rect 1918 3068 1922 3072
rect 1966 3068 1970 3072
rect 2014 3068 2018 3072
rect 2030 3068 2034 3072
rect 2094 3068 2098 3072
rect 2150 3068 2154 3072
rect 2182 3068 2186 3072
rect 2214 3068 2218 3072
rect 2254 3068 2258 3072
rect 2286 3068 2290 3072
rect 2318 3068 2322 3072
rect 2382 3068 2386 3072
rect 2430 3068 2434 3072
rect 2454 3068 2458 3072
rect 2486 3068 2490 3072
rect 2510 3068 2514 3072
rect 2526 3068 2530 3072
rect 2566 3068 2570 3072
rect 2614 3068 2618 3072
rect 2654 3068 2658 3072
rect 2678 3068 2682 3072
rect 2750 3068 2754 3072
rect 2766 3068 2770 3072
rect 2822 3068 2826 3072
rect 2878 3068 2882 3072
rect 2902 3068 2906 3072
rect 2910 3068 2914 3072
rect 2974 3068 2978 3072
rect 2990 3068 2994 3072
rect 2998 3068 3002 3072
rect 3022 3068 3026 3072
rect 3038 3068 3042 3072
rect 3062 3068 3066 3072
rect 3086 3068 3090 3072
rect 3110 3068 3114 3072
rect 3158 3068 3162 3072
rect 3182 3068 3186 3072
rect 3206 3068 3210 3072
rect 3230 3068 3234 3072
rect 3270 3068 3274 3072
rect 3454 3068 3458 3072
rect 3494 3068 3498 3072
rect 3518 3068 3522 3072
rect 3582 3068 3586 3072
rect 3630 3068 3634 3072
rect 3710 3068 3714 3072
rect 3726 3068 3730 3072
rect 3942 3068 3946 3072
rect 3998 3068 4002 3072
rect 4014 3068 4018 3072
rect 4118 3068 4122 3072
rect 4174 3068 4178 3072
rect 4294 3068 4298 3072
rect 4350 3068 4354 3072
rect 4390 3068 4394 3072
rect 4438 3068 4442 3072
rect 4462 3068 4466 3072
rect 4534 3068 4538 3072
rect 4566 3068 4570 3072
rect 6 3058 10 3062
rect 38 3058 42 3062
rect 78 3059 82 3063
rect 110 3058 114 3062
rect 174 3059 178 3063
rect 262 3058 266 3062
rect 294 3058 298 3062
rect 326 3058 330 3062
rect 430 3058 434 3062
rect 598 3058 602 3062
rect 622 3058 626 3062
rect 654 3058 658 3062
rect 702 3058 706 3062
rect 750 3058 754 3062
rect 846 3058 850 3062
rect 862 3058 866 3062
rect 934 3058 938 3062
rect 1046 3058 1050 3062
rect 1142 3058 1146 3062
rect 1230 3059 1234 3063
rect 1302 3058 1306 3062
rect 1366 3058 1370 3062
rect 1374 3058 1378 3062
rect 1406 3058 1410 3062
rect 1526 3058 1530 3062
rect 1542 3058 1546 3062
rect 1558 3058 1562 3062
rect 1590 3058 1594 3062
rect 1662 3059 1666 3063
rect 1758 3059 1762 3063
rect 1854 3059 1858 3063
rect 1950 3059 1954 3063
rect 2046 3059 2050 3063
rect 2102 3058 2106 3062
rect 2142 3058 2146 3062
rect 2174 3058 2178 3062
rect 2206 3058 2210 3062
rect 2238 3058 2242 3062
rect 2262 3058 2266 3062
rect 2294 3058 2298 3062
rect 2310 3058 2314 3062
rect 2366 3058 2370 3062
rect 2414 3058 2418 3062
rect 2462 3058 2466 3062
rect 2574 3058 2578 3062
rect 2598 3058 2602 3062
rect 2654 3058 2658 3062
rect 2702 3058 2706 3062
rect 2790 3058 2794 3062
rect 2918 3058 2922 3062
rect 2942 3058 2946 3062
rect 3294 3058 3298 3062
rect 3326 3058 3330 3062
rect 3382 3059 3386 3063
rect 3414 3058 3418 3062
rect 3494 3058 3498 3062
rect 3526 3058 3530 3062
rect 3542 3058 3546 3062
rect 3614 3059 3618 3063
rect 3686 3058 3690 3062
rect 3750 3058 3754 3062
rect 3862 3058 3866 3062
rect 3934 3059 3938 3063
rect 4030 3059 4034 3063
rect 4062 3058 4066 3062
rect 4126 3058 4130 3062
rect 4174 3058 4178 3062
rect 4206 3059 4210 3063
rect 4278 3058 4282 3062
rect 4302 3058 4306 3062
rect 4350 3058 4354 3062
rect 4358 3058 4362 3062
rect 4510 3058 4514 3062
rect 4542 3058 4546 3062
rect 46 3048 50 3052
rect 286 3048 290 3052
rect 350 3048 354 3052
rect 390 3048 394 3052
rect 494 3048 498 3052
rect 590 3048 594 3052
rect 718 3048 722 3052
rect 774 3048 778 3052
rect 782 3048 786 3052
rect 1326 3048 1330 3052
rect 1414 3048 1418 3052
rect 1462 3048 1466 3052
rect 1566 3048 1570 3052
rect 2206 3048 2210 3052
rect 2222 3048 2226 3052
rect 2278 3048 2282 3052
rect 2294 3048 2298 3052
rect 2438 3048 2442 3052
rect 2478 3048 2482 3052
rect 2510 3048 2514 3052
rect 2590 3048 2594 3052
rect 2598 3048 2602 3052
rect 2670 3048 2674 3052
rect 2726 3048 2730 3052
rect 2750 3048 2754 3052
rect 2774 3048 2778 3052
rect 2838 3048 2842 3052
rect 2862 3048 2866 3052
rect 2886 3048 2890 3052
rect 2934 3048 2938 3052
rect 2974 3048 2978 3052
rect 3014 3048 3018 3052
rect 3038 3048 3042 3052
rect 3046 3048 3050 3052
rect 3110 3048 3114 3052
rect 3126 3048 3130 3052
rect 3150 3048 3154 3052
rect 3174 3048 3178 3052
rect 3198 3048 3202 3052
rect 3222 3048 3226 3052
rect 3246 3048 3250 3052
rect 3254 3048 3258 3052
rect 3318 3048 3322 3052
rect 3470 3048 3474 3052
rect 3502 3048 3506 3052
rect 4150 3048 4154 3052
rect 4278 3048 4282 3052
rect 4318 3048 4322 3052
rect 4382 3048 4386 3052
rect 4406 3048 4410 3052
rect 4454 3048 4458 3052
rect 4470 3048 4474 3052
rect 4478 3048 4482 3052
rect 4526 3048 4530 3052
rect 4558 3048 4562 3052
rect 4582 3048 4586 3052
rect 30 3038 34 3042
rect 302 3038 306 3042
rect 606 3038 610 3042
rect 670 3038 674 3042
rect 990 3038 994 3042
rect 1382 3038 1386 3042
rect 2118 3038 2122 3042
rect 2158 3038 2162 3042
rect 2190 3038 2194 3042
rect 2310 3038 2314 3042
rect 2350 3038 2354 3042
rect 2406 3038 2410 3042
rect 2534 3038 2538 3042
rect 3270 3038 3274 3042
rect 3446 3038 3450 3042
rect 3790 3038 3794 3042
rect 4326 3038 4330 3042
rect 310 3018 314 3022
rect 526 3018 530 3022
rect 598 3018 602 3022
rect 742 3018 746 3022
rect 3142 3018 3146 3022
rect 3302 3018 3306 3022
rect 3342 3018 3346 3022
rect 3486 3018 3490 3022
rect 3678 3018 3682 3022
rect 3702 3018 3706 3022
rect 3806 3018 3810 3022
rect 4574 3018 4578 3022
rect 498 3003 502 3007
rect 505 3003 509 3007
rect 1522 3003 1526 3007
rect 1529 3003 1533 3007
rect 2546 3003 2550 3007
rect 2553 3003 2557 3007
rect 3570 3003 3574 3007
rect 3577 3003 3581 3007
rect 110 2988 114 2992
rect 190 2988 194 2992
rect 270 2988 274 2992
rect 374 2988 378 2992
rect 1182 2988 1186 2992
rect 1278 2988 1282 2992
rect 1286 2988 1290 2992
rect 1582 2988 1586 2992
rect 1854 2988 1858 2992
rect 2142 2988 2146 2992
rect 2158 2988 2162 2992
rect 2166 2988 2170 2992
rect 2294 2988 2298 2992
rect 2318 2988 2322 2992
rect 2566 2988 2570 2992
rect 2734 2988 2738 2992
rect 2910 2988 2914 2992
rect 3230 2988 3234 2992
rect 3454 2988 3458 2992
rect 3630 2988 3634 2992
rect 3878 2988 3882 2992
rect 4094 2988 4098 2992
rect 4278 2988 4282 2992
rect 4310 2988 4314 2992
rect 4358 2988 4362 2992
rect 4526 2988 4530 2992
rect 2310 2978 2314 2982
rect 590 2968 594 2972
rect 598 2968 602 2972
rect 990 2968 994 2972
rect 1014 2968 1018 2972
rect 1470 2968 1474 2972
rect 1870 2968 1874 2972
rect 1966 2968 1970 2972
rect 2470 2968 2474 2972
rect 2622 2968 2626 2972
rect 2638 2968 2642 2972
rect 2646 2968 2650 2972
rect 2694 2968 2698 2972
rect 2838 2968 2842 2972
rect 2886 2968 2890 2972
rect 2950 2968 2954 2972
rect 3054 2968 3058 2972
rect 3094 2968 3098 2972
rect 3118 2968 3122 2972
rect 3134 2968 3138 2972
rect 3182 2968 3186 2972
rect 3206 2968 3210 2972
rect 3262 2968 3266 2972
rect 3270 2968 3274 2972
rect 3286 2968 3290 2972
rect 3846 2968 3850 2972
rect 4558 2968 4562 2972
rect 494 2958 498 2962
rect 46 2947 50 2951
rect 150 2948 154 2952
rect 254 2948 258 2952
rect 310 2947 314 2951
rect 342 2948 346 2952
rect 406 2947 410 2951
rect 438 2948 442 2952
rect 534 2958 538 2962
rect 550 2958 554 2962
rect 1078 2958 1082 2962
rect 1422 2958 1426 2962
rect 2262 2958 2266 2962
rect 2414 2958 2418 2962
rect 534 2948 538 2952
rect 582 2948 586 2952
rect 630 2948 634 2952
rect 638 2948 642 2952
rect 670 2948 674 2952
rect 678 2948 682 2952
rect 710 2948 714 2952
rect 718 2948 722 2952
rect 782 2948 786 2952
rect 790 2948 794 2952
rect 822 2948 826 2952
rect 14 2938 18 2942
rect 62 2938 66 2942
rect 158 2938 162 2942
rect 246 2938 250 2942
rect 478 2938 482 2942
rect 542 2938 546 2942
rect 566 2938 570 2942
rect 622 2938 626 2942
rect 646 2938 650 2942
rect 662 2938 666 2942
rect 686 2938 690 2942
rect 702 2938 706 2942
rect 734 2938 738 2942
rect 926 2947 930 2951
rect 1070 2948 1074 2952
rect 1126 2948 1130 2952
rect 1222 2948 1226 2952
rect 1350 2947 1354 2951
rect 1382 2948 1386 2952
rect 1398 2948 1402 2952
rect 1414 2948 1418 2952
rect 1534 2947 1538 2951
rect 1662 2947 1666 2951
rect 1758 2947 1762 2951
rect 1814 2948 1818 2952
rect 1846 2948 1850 2952
rect 1910 2948 1914 2952
rect 2014 2947 2018 2951
rect 2230 2947 2234 2951
rect 2382 2947 2386 2951
rect 2454 2948 2458 2952
rect 2502 2958 2506 2962
rect 2510 2958 2514 2962
rect 2542 2958 2546 2962
rect 2662 2958 2666 2962
rect 2718 2958 2722 2962
rect 2766 2958 2770 2962
rect 2806 2958 2810 2962
rect 2486 2948 2490 2952
rect 2510 2948 2514 2952
rect 2566 2948 2570 2952
rect 2734 2948 2738 2952
rect 2790 2948 2794 2952
rect 2910 2948 2914 2952
rect 2934 2958 2938 2962
rect 2974 2958 2978 2962
rect 3022 2958 3026 2962
rect 3030 2958 3034 2962
rect 3214 2958 3218 2962
rect 3358 2958 3362 2962
rect 3646 2958 3650 2962
rect 3710 2958 3714 2962
rect 4350 2958 4354 2962
rect 4510 2958 4514 2962
rect 4550 2958 4554 2962
rect 4558 2958 4562 2962
rect 2982 2948 2986 2952
rect 3230 2948 3234 2952
rect 3342 2948 3346 2952
rect 750 2938 754 2942
rect 774 2938 778 2942
rect 798 2938 802 2942
rect 814 2938 818 2942
rect 830 2938 834 2942
rect 894 2938 898 2942
rect 910 2938 914 2942
rect 998 2938 1002 2942
rect 1038 2938 1042 2942
rect 1070 2938 1074 2942
rect 1134 2938 1138 2942
rect 1222 2938 1226 2942
rect 1342 2938 1346 2942
rect 1382 2938 1386 2942
rect 1406 2938 1410 2942
rect 1446 2938 1450 2942
rect 1550 2938 1554 2942
rect 1678 2938 1682 2942
rect 1742 2938 1746 2942
rect 1918 2938 1922 2942
rect 2030 2938 2034 2942
rect 2054 2938 2058 2942
rect 2126 2938 2130 2942
rect 2278 2938 2282 2942
rect 2366 2938 2370 2942
rect 2430 2938 2434 2942
rect 2454 2938 2458 2942
rect 2478 2938 2482 2942
rect 2510 2938 2514 2942
rect 2534 2938 2538 2942
rect 2598 2938 2602 2942
rect 2622 2938 2626 2942
rect 2662 2938 2666 2942
rect 2686 2938 2690 2942
rect 2710 2938 2714 2942
rect 2758 2938 2762 2942
rect 2806 2938 2810 2942
rect 2830 2938 2834 2942
rect 2862 2938 2866 2942
rect 2958 2938 2962 2942
rect 2974 2938 2978 2942
rect 3390 2947 3394 2951
rect 3422 2948 3426 2952
rect 3486 2947 3490 2951
rect 3518 2948 3522 2952
rect 3662 2948 3666 2952
rect 3726 2948 3730 2952
rect 3782 2947 3786 2951
rect 3854 2948 3858 2952
rect 3918 2948 3922 2952
rect 3998 2947 4002 2951
rect 4198 2947 4202 2951
rect 4270 2948 4274 2952
rect 4286 2948 4290 2952
rect 4318 2948 4322 2952
rect 4334 2948 4338 2952
rect 2998 2938 3002 2942
rect 3006 2938 3010 2942
rect 3030 2938 3034 2942
rect 3070 2938 3074 2942
rect 3086 2938 3090 2942
rect 3118 2938 3122 2942
rect 3134 2938 3138 2942
rect 3158 2938 3162 2942
rect 3166 2938 3170 2942
rect 3190 2938 3194 2942
rect 3238 2938 3242 2942
rect 3246 2938 3250 2942
rect 3286 2938 3290 2942
rect 3310 2938 3314 2942
rect 3358 2938 3362 2942
rect 3574 2938 3578 2942
rect 3718 2938 3722 2942
rect 3790 2938 3794 2942
rect 3870 2938 3874 2942
rect 4014 2938 4018 2942
rect 4102 2938 4106 2942
rect 4166 2938 4170 2942
rect 4182 2938 4186 2942
rect 4398 2947 4402 2951
rect 4486 2948 4490 2952
rect 4566 2948 4570 2952
rect 4294 2938 4298 2942
rect 4318 2938 4322 2942
rect 4326 2938 4330 2942
rect 4382 2938 4386 2942
rect 4534 2938 4538 2942
rect 4550 2938 4554 2942
rect 6 2928 10 2932
rect 166 2928 170 2932
rect 606 2928 610 2932
rect 1086 2928 1090 2932
rect 1462 2928 1466 2932
rect 2134 2928 2138 2932
rect 2150 2928 2154 2932
rect 2230 2928 2234 2932
rect 2286 2928 2290 2932
rect 2302 2928 2306 2932
rect 2438 2928 2442 2932
rect 2446 2928 2450 2932
rect 2590 2928 2594 2932
rect 2758 2928 2762 2932
rect 2822 2928 2826 2932
rect 2886 2928 2890 2932
rect 3014 2928 3018 2932
rect 3318 2928 3322 2932
rect 3686 2928 3690 2932
rect 3694 2928 3698 2932
rect 3750 2928 3754 2932
rect 4366 2928 4370 2932
rect 4462 2928 4466 2932
rect 4470 2928 4474 2932
rect 4518 2928 4522 2932
rect 158 2918 162 2922
rect 190 2918 194 2922
rect 270 2918 274 2922
rect 470 2918 474 2922
rect 614 2918 618 2922
rect 654 2918 658 2922
rect 694 2918 698 2922
rect 766 2918 770 2922
rect 806 2918 810 2922
rect 1694 2918 1698 2922
rect 1798 2918 1802 2922
rect 1830 2918 1834 2922
rect 1950 2918 1954 2922
rect 2262 2918 2266 2922
rect 2414 2918 2418 2922
rect 2614 2918 2618 2922
rect 2638 2918 2642 2922
rect 2654 2918 2658 2922
rect 2670 2918 2674 2922
rect 2694 2918 2698 2922
rect 2846 2918 2850 2922
rect 2870 2918 2874 2922
rect 2966 2918 2970 2922
rect 3078 2918 3082 2922
rect 3102 2918 3106 2922
rect 3118 2918 3122 2922
rect 3150 2918 3154 2922
rect 3182 2918 3186 2922
rect 3206 2918 3210 2922
rect 3262 2918 3266 2922
rect 3278 2918 3282 2922
rect 3302 2918 3306 2922
rect 3550 2918 3554 2922
rect 3646 2918 3650 2922
rect 3702 2918 3706 2922
rect 3854 2918 3858 2922
rect 3318 2908 3322 2912
rect 3686 2908 3690 2912
rect 3694 2908 3698 2912
rect 3750 2908 3754 2912
rect 1002 2903 1006 2907
rect 1009 2903 1013 2907
rect 2026 2903 2030 2907
rect 2033 2903 2037 2907
rect 3050 2903 3054 2907
rect 3057 2903 3061 2907
rect 4082 2903 4086 2907
rect 4089 2903 4093 2907
rect 2886 2898 2890 2902
rect 3070 2898 3074 2902
rect 3150 2898 3154 2902
rect 3478 2898 3482 2902
rect 3550 2898 3554 2902
rect 3710 2898 3714 2902
rect 3886 2898 3890 2902
rect 3894 2898 3898 2902
rect 46 2888 50 2892
rect 254 2888 258 2892
rect 462 2888 466 2892
rect 510 2888 514 2892
rect 574 2888 578 2892
rect 598 2888 602 2892
rect 662 2888 666 2892
rect 982 2888 986 2892
rect 1086 2888 1090 2892
rect 1094 2888 1098 2892
rect 1278 2888 1282 2892
rect 1374 2888 1378 2892
rect 1382 2888 1386 2892
rect 1494 2888 1498 2892
rect 1846 2888 1850 2892
rect 1942 2888 1946 2892
rect 2054 2888 2058 2892
rect 2150 2888 2154 2892
rect 2246 2888 2250 2892
rect 2342 2888 2346 2892
rect 2438 2888 2442 2892
rect 2542 2888 2546 2892
rect 2670 2888 2674 2892
rect 2718 2888 2722 2892
rect 2750 2888 2754 2892
rect 2774 2888 2778 2892
rect 2790 2888 2794 2892
rect 2902 2888 2906 2892
rect 3126 2888 3130 2892
rect 3238 2888 3242 2892
rect 3278 2888 3282 2892
rect 3326 2888 3330 2892
rect 3342 2888 3346 2892
rect 4030 2888 4034 2892
rect 4238 2888 4242 2892
rect 4334 2888 4338 2892
rect 4358 2888 4362 2892
rect 4406 2888 4410 2892
rect 6 2878 10 2882
rect 22 2878 26 2882
rect 78 2878 82 2882
rect 86 2878 90 2882
rect 158 2878 162 2882
rect 190 2878 194 2882
rect 318 2878 322 2882
rect 334 2878 338 2882
rect 62 2868 66 2872
rect 102 2868 106 2872
rect 134 2868 138 2872
rect 438 2868 442 2872
rect 542 2878 546 2882
rect 614 2878 618 2882
rect 670 2878 674 2882
rect 742 2878 746 2882
rect 862 2878 866 2882
rect 950 2878 954 2882
rect 1022 2878 1026 2882
rect 1630 2878 1634 2882
rect 1838 2878 1842 2882
rect 2886 2878 2890 2882
rect 2982 2878 2986 2882
rect 3070 2878 3074 2882
rect 3150 2878 3154 2882
rect 3334 2878 3338 2882
rect 3478 2878 3482 2882
rect 3550 2878 3554 2882
rect 3710 2878 3714 2882
rect 3886 2878 3890 2882
rect 3894 2878 3898 2882
rect 4142 2878 4146 2882
rect 4454 2878 4458 2882
rect 478 2868 482 2872
rect 494 2868 498 2872
rect 550 2868 554 2872
rect 582 2868 586 2872
rect 662 2868 666 2872
rect 710 2868 714 2872
rect 886 2868 890 2872
rect 918 2868 922 2872
rect 958 2868 962 2872
rect 1134 2868 1138 2872
rect 1222 2868 1226 2872
rect 1294 2868 1298 2872
rect 1462 2868 1466 2872
rect 1550 2868 1554 2872
rect 1590 2868 1594 2872
rect 1646 2868 1650 2872
rect 1662 2868 1666 2872
rect 1678 2868 1682 2872
rect 1742 2868 1746 2872
rect 1774 2868 1778 2872
rect 1806 2868 1810 2872
rect 1822 2868 1826 2872
rect 1838 2868 1842 2872
rect 1926 2868 1930 2872
rect 2022 2868 2026 2872
rect 2230 2868 2234 2872
rect 2326 2868 2330 2872
rect 2422 2868 2426 2872
rect 2518 2868 2522 2872
rect 2566 2868 2570 2872
rect 2606 2868 2610 2872
rect 2630 2868 2634 2872
rect 2678 2868 2682 2872
rect 2710 2868 2714 2872
rect 2750 2868 2754 2872
rect 2774 2868 2778 2872
rect 2838 2868 2842 2872
rect 2886 2868 2890 2872
rect 2910 2868 2914 2872
rect 2958 2868 2962 2872
rect 3014 2868 3018 2872
rect 3222 2868 3226 2872
rect 3246 2868 3250 2872
rect 3254 2868 3258 2872
rect 3318 2868 3322 2872
rect 3422 2868 3426 2872
rect 3502 2868 3506 2872
rect 3598 2868 3602 2872
rect 3710 2868 3714 2872
rect 3758 2868 3762 2872
rect 54 2858 58 2862
rect 134 2858 138 2862
rect 190 2859 194 2863
rect 294 2858 298 2862
rect 366 2859 370 2863
rect 390 2858 394 2862
rect 518 2858 522 2862
rect 558 2858 562 2862
rect 630 2858 634 2862
rect 654 2858 658 2862
rect 694 2858 698 2862
rect 702 2858 706 2862
rect 742 2859 746 2863
rect 814 2858 818 2862
rect 878 2858 882 2862
rect 894 2858 898 2862
rect 910 2858 914 2862
rect 1030 2858 1034 2862
rect 1158 2859 1162 2863
rect 1214 2859 1218 2863
rect 1310 2859 1314 2863
rect 1446 2859 1450 2863
rect 1558 2859 1562 2863
rect 1598 2858 1602 2862
rect 1614 2858 1618 2862
rect 1638 2858 1642 2862
rect 1670 2858 1674 2862
rect 1766 2858 1770 2862
rect 1910 2859 1914 2863
rect 2006 2859 2010 2863
rect 2086 2858 2090 2862
rect 2118 2859 2122 2863
rect 2182 2858 2186 2862
rect 2214 2859 2218 2863
rect 2310 2859 2314 2863
rect 2374 2858 2378 2862
rect 2406 2859 2410 2863
rect 2478 2858 2482 2862
rect 2502 2859 2506 2863
rect 2574 2858 2578 2862
rect 2598 2858 2602 2862
rect 2654 2858 2658 2862
rect 2702 2858 2706 2862
rect 2726 2858 2730 2862
rect 2806 2858 2810 2862
rect 2814 2858 2818 2862
rect 2854 2858 2858 2862
rect 2862 2858 2866 2862
rect 2942 2858 2946 2862
rect 2966 2858 2970 2862
rect 3046 2858 3050 2862
rect 3094 2858 3098 2862
rect 3118 2858 3122 2862
rect 3142 2858 3146 2862
rect 3174 2858 3178 2862
rect 3190 2858 3194 2862
rect 3294 2858 3298 2862
rect 3398 2858 3402 2862
rect 3454 2858 3458 2862
rect 3518 2858 3522 2862
rect 3526 2858 3530 2862
rect 3606 2858 3610 2862
rect 3694 2858 3698 2862
rect 3726 2858 3730 2862
rect 3734 2858 3738 2862
rect 3774 2859 3778 2863
rect 3950 2868 3954 2872
rect 4158 2868 4162 2872
rect 4254 2868 4258 2872
rect 4342 2868 4346 2872
rect 4398 2868 4402 2872
rect 4422 2868 4426 2872
rect 4582 2868 4586 2872
rect 4598 2868 4602 2872
rect 3846 2858 3850 2862
rect 3862 2858 3866 2862
rect 3918 2858 3922 2862
rect 3966 2859 3970 2863
rect 4078 2859 4082 2863
rect 4110 2858 4114 2862
rect 4174 2859 4178 2863
rect 4270 2859 4274 2863
rect 4382 2858 4386 2862
rect 4390 2858 4394 2862
rect 4422 2858 4426 2862
rect 4454 2859 4458 2863
rect 4478 2858 4482 2862
rect 4558 2858 4562 2862
rect 118 2849 122 2853
rect 278 2849 282 2853
rect 494 2848 498 2852
rect 574 2848 578 2852
rect 686 2848 690 2852
rect 838 2848 842 2852
rect 942 2848 946 2852
rect 974 2848 978 2852
rect 1614 2848 1618 2852
rect 1646 2848 1650 2852
rect 1750 2848 1754 2852
rect 1782 2848 1786 2852
rect 2534 2848 2538 2852
rect 2606 2848 2610 2852
rect 2622 2848 2626 2852
rect 2670 2848 2674 2852
rect 2726 2848 2730 2852
rect 2758 2848 2762 2852
rect 2774 2848 2778 2852
rect 2846 2848 2850 2852
rect 2910 2848 2914 2852
rect 2950 2848 2954 2852
rect 2998 2848 3002 2852
rect 3190 2848 3194 2852
rect 3230 2848 3234 2852
rect 3270 2848 3274 2852
rect 3438 2848 3442 2852
rect 3478 2848 3482 2852
rect 3510 2848 3514 2852
rect 3670 2848 3674 2852
rect 3742 2848 3746 2852
rect 3846 2848 3850 2852
rect 3934 2848 3938 2852
rect 4358 2848 4362 2852
rect 4542 2848 4546 2852
rect 4582 2848 4586 2852
rect 430 2838 434 2842
rect 446 2838 450 2842
rect 2262 2838 2266 2842
rect 3502 2838 3506 2842
rect 4014 2838 4018 2842
rect 4566 2838 4570 2842
rect 542 2828 546 2832
rect 806 2828 810 2832
rect 3662 2828 3666 2832
rect 590 2818 594 2822
rect 630 2818 634 2822
rect 814 2818 818 2822
rect 1686 2818 1690 2822
rect 3006 2818 3010 2822
rect 3030 2818 3034 2822
rect 3094 2818 3098 2822
rect 3174 2818 3178 2822
rect 3454 2818 3458 2822
rect 3686 2818 3690 2822
rect 3838 2818 3842 2822
rect 3918 2818 3922 2822
rect 4030 2818 4034 2822
rect 498 2803 502 2807
rect 505 2803 509 2807
rect 1522 2803 1526 2807
rect 1529 2803 1533 2807
rect 2546 2803 2550 2807
rect 2553 2803 2557 2807
rect 3570 2803 3574 2807
rect 3577 2803 3581 2807
rect 990 2788 994 2792
rect 1182 2788 1186 2792
rect 1734 2788 1738 2792
rect 1902 2788 1906 2792
rect 2190 2788 2194 2792
rect 2926 2788 2930 2792
rect 3078 2788 3082 2792
rect 4094 2788 4098 2792
rect 4222 2788 4226 2792
rect 4414 2788 4418 2792
rect 4598 2788 4602 2792
rect 1910 2778 1914 2782
rect 2094 2778 2098 2782
rect 2542 2778 2546 2782
rect 3742 2778 3746 2782
rect 254 2768 258 2772
rect 1278 2768 1282 2772
rect 1470 2768 1474 2772
rect 1926 2768 1930 2772
rect 2358 2768 2362 2772
rect 2382 2768 2386 2772
rect 2406 2768 2410 2772
rect 2438 2768 2442 2772
rect 2734 2768 2738 2772
rect 2774 2768 2778 2772
rect 2822 2768 2826 2772
rect 2838 2768 2842 2772
rect 2918 2768 2922 2772
rect 3726 2768 3730 2772
rect 4078 2768 4082 2772
rect 350 2758 354 2762
rect 470 2758 474 2762
rect 614 2758 618 2762
rect 630 2758 634 2762
rect 694 2758 698 2762
rect 822 2758 826 2762
rect 854 2758 858 2762
rect 1886 2758 1890 2762
rect 22 2748 26 2752
rect 38 2748 42 2752
rect 102 2748 106 2752
rect 134 2748 138 2752
rect 6 2738 10 2742
rect 190 2747 194 2751
rect 302 2748 306 2752
rect 398 2748 402 2752
rect 550 2748 554 2752
rect 590 2748 594 2752
rect 622 2748 626 2752
rect 638 2748 642 2752
rect 646 2748 650 2752
rect 686 2748 690 2752
rect 710 2748 714 2752
rect 758 2748 762 2752
rect 830 2748 834 2752
rect 838 2748 842 2752
rect 870 2748 874 2752
rect 910 2747 914 2751
rect 1022 2747 1026 2751
rect 1118 2747 1122 2751
rect 1238 2748 1242 2752
rect 1310 2747 1314 2751
rect 1414 2748 1418 2752
rect 1518 2747 1522 2751
rect 1550 2748 1554 2752
rect 1590 2748 1594 2752
rect 1678 2748 1682 2752
rect 1726 2748 1730 2752
rect 1758 2748 1762 2752
rect 1766 2748 1770 2752
rect 1782 2748 1786 2752
rect 1798 2748 1802 2752
rect 1806 2748 1810 2752
rect 1822 2748 1826 2752
rect 1846 2748 1850 2752
rect 1974 2747 1978 2751
rect 2022 2748 2026 2752
rect 2134 2748 2138 2752
rect 2334 2758 2338 2762
rect 2478 2758 2482 2762
rect 2614 2758 2618 2762
rect 2662 2758 2666 2762
rect 2710 2758 2714 2762
rect 2846 2758 2850 2762
rect 2934 2758 2938 2762
rect 2942 2758 2946 2762
rect 3006 2758 3010 2762
rect 3062 2758 3066 2762
rect 3102 2758 3106 2762
rect 3198 2758 3202 2762
rect 3246 2758 3250 2762
rect 3350 2758 3354 2762
rect 3398 2758 3402 2762
rect 3646 2758 3650 2762
rect 3750 2758 3754 2762
rect 3798 2758 3802 2762
rect 3982 2758 3986 2762
rect 4302 2758 4306 2762
rect 2158 2747 2162 2751
rect 2254 2747 2258 2751
rect 2318 2748 2322 2752
rect 2326 2748 2330 2752
rect 2462 2748 2466 2752
rect 2598 2748 2602 2752
rect 2646 2748 2650 2752
rect 2694 2748 2698 2752
rect 2766 2748 2770 2752
rect 2862 2748 2866 2752
rect 2942 2748 2946 2752
rect 2958 2748 2962 2752
rect 3046 2748 3050 2752
rect 3078 2748 3082 2752
rect 3126 2748 3130 2752
rect 3182 2748 3186 2752
rect 3222 2748 3226 2752
rect 3246 2748 3250 2752
rect 3278 2747 3282 2751
rect 3310 2748 3314 2752
rect 3366 2748 3370 2752
rect 3414 2748 3418 2752
rect 3470 2747 3474 2751
rect 3502 2748 3506 2752
rect 3582 2747 3586 2751
rect 3678 2747 3682 2751
rect 3870 2747 3874 2751
rect 4030 2747 4034 2751
rect 4158 2747 4162 2751
rect 4238 2748 4242 2752
rect 4262 2748 4266 2752
rect 4302 2748 4306 2752
rect 4374 2748 4378 2752
rect 4462 2748 4466 2752
rect 78 2738 82 2742
rect 142 2738 146 2742
rect 206 2738 210 2742
rect 302 2738 306 2742
rect 390 2738 394 2742
rect 398 2738 402 2742
rect 502 2738 506 2742
rect 598 2738 602 2742
rect 614 2738 618 2742
rect 654 2738 658 2742
rect 718 2738 722 2742
rect 734 2738 738 2742
rect 846 2738 850 2742
rect 862 2738 866 2742
rect 878 2738 882 2742
rect 926 2738 930 2742
rect 1030 2738 1034 2742
rect 1102 2738 1106 2742
rect 1222 2738 1226 2742
rect 1590 2738 1594 2742
rect 1614 2738 1618 2742
rect 1686 2738 1690 2742
rect 1726 2738 1730 2742
rect 1750 2738 1754 2742
rect 1758 2738 1762 2742
rect 1790 2738 1794 2742
rect 1806 2738 1810 2742
rect 1830 2738 1834 2742
rect 1862 2738 1866 2742
rect 1990 2738 1994 2742
rect 2086 2738 2090 2742
rect 2222 2738 2226 2742
rect 2270 2738 2274 2742
rect 2286 2738 2290 2742
rect 2302 2738 2306 2742
rect 2310 2738 2314 2742
rect 2342 2738 2346 2742
rect 2366 2738 2370 2742
rect 2390 2738 2394 2742
rect 2414 2738 2418 2742
rect 2486 2738 2490 2742
rect 2702 2738 2706 2742
rect 2718 2738 2722 2742
rect 2742 2738 2746 2742
rect 2798 2738 2802 2742
rect 2822 2738 2826 2742
rect 2894 2738 2898 2742
rect 2918 2738 2922 2742
rect 2990 2738 2994 2742
rect 3014 2738 3018 2742
rect 3406 2738 3410 2742
rect 3566 2738 3570 2742
rect 3662 2738 3666 2742
rect 3774 2738 3778 2742
rect 3822 2738 3826 2742
rect 3854 2738 3858 2742
rect 3982 2738 3986 2742
rect 3998 2738 4002 2742
rect 4014 2738 4018 2742
rect 4118 2738 4122 2742
rect 4142 2738 4146 2742
rect 4230 2738 4234 2742
rect 4286 2738 4290 2742
rect 4534 2747 4538 2751
rect 4310 2738 4314 2742
rect 4350 2738 4354 2742
rect 4398 2738 4402 2742
rect 4478 2738 4482 2742
rect 22 2728 26 2732
rect 86 2728 90 2732
rect 158 2728 162 2732
rect 558 2728 562 2732
rect 1310 2728 1314 2732
rect 1406 2728 1410 2732
rect 1846 2728 1850 2732
rect 1894 2728 1898 2732
rect 2438 2728 2442 2732
rect 2574 2728 2578 2732
rect 2622 2728 2626 2732
rect 2670 2728 2674 2732
rect 2886 2728 2890 2732
rect 2982 2728 2986 2732
rect 3102 2728 3106 2732
rect 3150 2728 3154 2732
rect 3158 2728 3162 2732
rect 3206 2728 3210 2732
rect 3278 2728 3282 2732
rect 3390 2728 3394 2732
rect 3438 2728 3442 2732
rect 3790 2728 3794 2732
rect 3838 2728 3842 2732
rect 3942 2728 3946 2732
rect 4278 2728 4282 2732
rect 4310 2728 4314 2732
rect 4406 2728 4410 2732
rect 78 2718 82 2722
rect 142 2718 146 2722
rect 486 2718 490 2722
rect 670 2718 674 2722
rect 694 2718 698 2722
rect 814 2718 818 2722
rect 974 2718 978 2722
rect 1086 2718 1090 2722
rect 1374 2718 1378 2722
rect 1582 2718 1586 2722
rect 1606 2718 1610 2722
rect 2350 2718 2354 2722
rect 2374 2718 2378 2722
rect 2398 2718 2402 2722
rect 2430 2718 2434 2722
rect 2478 2718 2482 2722
rect 2542 2718 2546 2722
rect 2614 2718 2618 2722
rect 2662 2718 2666 2722
rect 2726 2718 2730 2722
rect 2774 2718 2778 2722
rect 2806 2718 2810 2722
rect 2830 2718 2834 2722
rect 2846 2718 2850 2722
rect 2902 2718 2906 2722
rect 3022 2718 3026 2722
rect 3110 2718 3114 2722
rect 3198 2718 3202 2722
rect 3342 2718 3346 2722
rect 3350 2718 3354 2722
rect 3550 2718 3554 2722
rect 3934 2718 3938 2722
rect 3966 2718 3970 2722
rect 3990 2718 3994 2722
rect 4126 2718 4130 2722
rect 4254 2718 4258 2722
rect 4270 2718 4274 2722
rect 4358 2718 4362 2722
rect 2438 2708 2442 2712
rect 2574 2708 2578 2712
rect 2622 2708 2626 2712
rect 2670 2708 2674 2712
rect 2886 2708 2890 2712
rect 3150 2708 3154 2712
rect 3158 2708 3162 2712
rect 3206 2708 3210 2712
rect 3390 2708 3394 2712
rect 3438 2708 3442 2712
rect 1002 2703 1006 2707
rect 1009 2703 1013 2707
rect 2026 2703 2030 2707
rect 2033 2703 2037 2707
rect 3050 2703 3054 2707
rect 3057 2703 3061 2707
rect 4082 2703 4086 2707
rect 4089 2703 4093 2707
rect 2214 2698 2218 2702
rect 2262 2698 2266 2702
rect 2310 2698 2314 2702
rect 2926 2698 2930 2702
rect 78 2688 82 2692
rect 870 2688 874 2692
rect 1078 2688 1082 2692
rect 1174 2688 1178 2692
rect 1270 2688 1274 2692
rect 1462 2688 1466 2692
rect 1558 2688 1562 2692
rect 1670 2688 1674 2692
rect 1702 2688 1706 2692
rect 1798 2688 1802 2692
rect 1894 2688 1898 2692
rect 2022 2688 2026 2692
rect 2118 2688 2122 2692
rect 2366 2688 2370 2692
rect 2390 2688 2394 2692
rect 2486 2688 2490 2692
rect 2950 2688 2954 2692
rect 2990 2688 2994 2692
rect 3038 2688 3042 2692
rect 3102 2688 3106 2692
rect 3358 2688 3362 2692
rect 3430 2688 3434 2692
rect 3518 2688 3522 2692
rect 3782 2688 3786 2692
rect 4358 2688 4362 2692
rect 4390 2688 4394 2692
rect 4598 2688 4602 2692
rect 6 2678 10 2682
rect 14 2678 18 2682
rect 22 2678 26 2682
rect 86 2678 90 2682
rect 158 2678 162 2682
rect 502 2678 506 2682
rect 574 2678 578 2682
rect 582 2678 586 2682
rect 630 2678 634 2682
rect 646 2678 650 2682
rect 718 2678 722 2682
rect 2182 2678 2186 2682
rect 2214 2678 2218 2682
rect 2262 2678 2266 2682
rect 2310 2678 2314 2682
rect 2750 2678 2754 2682
rect 2926 2678 2930 2682
rect 3094 2678 3098 2682
rect 3230 2678 3234 2682
rect 3662 2678 3666 2682
rect 3710 2678 3714 2682
rect 3790 2678 3794 2682
rect 3798 2678 3802 2682
rect 3806 2678 3810 2682
rect 4030 2678 4034 2682
rect 4038 2678 4042 2682
rect 4214 2678 4218 2682
rect 4246 2678 4250 2682
rect 4262 2678 4266 2682
rect 4334 2678 4338 2682
rect 4350 2678 4354 2682
rect 4478 2678 4482 2682
rect 38 2668 42 2672
rect 78 2668 82 2672
rect 126 2668 130 2672
rect 142 2668 146 2672
rect 206 2668 210 2672
rect 302 2668 306 2672
rect 398 2668 402 2672
rect 598 2668 602 2672
rect 614 2668 618 2672
rect 654 2668 658 2672
rect 686 2668 690 2672
rect 702 2668 706 2672
rect 742 2668 746 2672
rect 774 2668 778 2672
rect 886 2668 890 2672
rect 1030 2668 1034 2672
rect 1222 2668 1226 2672
rect 1310 2668 1314 2672
rect 1382 2668 1386 2672
rect 1406 2668 1410 2672
rect 1478 2668 1482 2672
rect 1574 2668 1578 2672
rect 1614 2668 1618 2672
rect 1654 2668 1658 2672
rect 1670 2668 1674 2672
rect 1694 2668 1698 2672
rect 1990 2668 1994 2672
rect 2102 2668 2106 2672
rect 2582 2668 2586 2672
rect 2606 2668 2610 2672
rect 2718 2668 2722 2672
rect 2934 2668 2938 2672
rect 2950 2668 2954 2672
rect 3030 2668 3034 2672
rect 3182 2668 3186 2672
rect 70 2658 74 2662
rect 134 2658 138 2662
rect 190 2658 194 2662
rect 222 2659 226 2663
rect 254 2658 258 2662
rect 318 2659 322 2663
rect 350 2658 354 2662
rect 414 2659 418 2663
rect 486 2658 490 2662
rect 542 2658 546 2662
rect 566 2658 570 2662
rect 590 2658 594 2662
rect 606 2658 610 2662
rect 622 2658 626 2662
rect 646 2658 650 2662
rect 670 2658 674 2662
rect 694 2658 698 2662
rect 710 2658 714 2662
rect 734 2658 738 2662
rect 758 2658 762 2662
rect 766 2658 770 2662
rect 814 2658 818 2662
rect 838 2658 842 2662
rect 902 2659 906 2663
rect 934 2658 938 2662
rect 1014 2659 1018 2663
rect 1118 2658 1122 2662
rect 1142 2658 1146 2662
rect 1214 2658 1218 2662
rect 1326 2658 1330 2662
rect 1334 2658 1338 2662
rect 1398 2659 1402 2663
rect 1494 2659 1498 2663
rect 1590 2658 1594 2662
rect 1622 2658 1626 2662
rect 1638 2658 1642 2662
rect 1662 2658 1666 2662
rect 1694 2658 1698 2662
rect 1734 2658 1738 2662
rect 1766 2659 1770 2663
rect 1830 2658 1834 2662
rect 1862 2659 1866 2663
rect 1974 2659 1978 2663
rect 2086 2659 2090 2663
rect 2182 2659 2186 2663
rect 2238 2658 2242 2662
rect 2286 2658 2290 2662
rect 2334 2658 2338 2662
rect 2342 2658 2346 2662
rect 2382 2658 2386 2662
rect 2422 2658 2426 2662
rect 2454 2659 2458 2663
rect 2518 2658 2522 2662
rect 2550 2659 2554 2663
rect 2630 2658 2634 2662
rect 2726 2658 2730 2662
rect 2822 2658 2826 2662
rect 2854 2659 2858 2663
rect 3278 2668 3282 2672
rect 3342 2668 3346 2672
rect 3366 2668 3370 2672
rect 3382 2668 3386 2672
rect 3414 2668 3418 2672
rect 3438 2668 3442 2672
rect 3462 2668 3466 2672
rect 3534 2668 3538 2672
rect 3598 2668 3602 2672
rect 3646 2668 3650 2672
rect 3694 2668 3698 2672
rect 3742 2668 3746 2672
rect 3774 2668 3778 2672
rect 3854 2668 3858 2672
rect 3910 2668 3914 2672
rect 3942 2668 3946 2672
rect 4022 2668 4026 2672
rect 4054 2668 4058 2672
rect 4094 2668 4098 2672
rect 4126 2668 4130 2672
rect 4214 2668 4218 2672
rect 4230 2668 4234 2672
rect 4278 2668 4282 2672
rect 4310 2668 4314 2672
rect 4382 2668 4386 2672
rect 4406 2668 4410 2672
rect 4422 2668 4426 2672
rect 2902 2658 2906 2662
rect 2982 2658 2986 2662
rect 3006 2658 3010 2662
rect 3078 2658 3082 2662
rect 3158 2658 3162 2662
rect 3198 2658 3202 2662
rect 3214 2658 3218 2662
rect 3270 2659 3274 2663
rect 3382 2658 3386 2662
rect 3462 2658 3466 2662
rect 3734 2658 3738 2662
rect 3766 2658 3770 2662
rect 3838 2659 3842 2663
rect 3910 2658 3914 2662
rect 3966 2658 3970 2662
rect 3998 2658 4002 2662
rect 4054 2658 4058 2662
rect 4158 2658 4162 2662
rect 4198 2658 4202 2662
rect 4278 2658 4282 2662
rect 4286 2658 4290 2662
rect 4302 2658 4306 2662
rect 4318 2658 4322 2662
rect 4374 2658 4378 2662
rect 4454 2658 4458 2662
rect 4558 2658 4562 2662
rect 718 2648 722 2652
rect 750 2648 754 2652
rect 1606 2648 1610 2652
rect 1638 2648 1642 2652
rect 2254 2648 2258 2652
rect 2302 2648 2306 2652
rect 2350 2648 2354 2652
rect 2806 2648 2810 2652
rect 2886 2648 2890 2652
rect 2950 2648 2954 2652
rect 2990 2648 2994 2652
rect 3038 2648 3042 2652
rect 3198 2648 3202 2652
rect 3358 2648 3362 2652
rect 3382 2648 3386 2652
rect 3406 2648 3410 2652
rect 3430 2648 3434 2652
rect 3454 2648 3458 2652
rect 3622 2648 3626 2652
rect 3670 2648 3674 2652
rect 3718 2648 3722 2652
rect 3750 2648 3754 2652
rect 3934 2648 3938 2652
rect 3958 2648 3962 2652
rect 4070 2648 4074 2652
rect 4142 2648 4146 2652
rect 4206 2648 4210 2652
rect 4390 2648 4394 2652
rect 478 2638 482 2642
rect 966 2638 970 2642
rect 1366 2638 1370 2642
rect 1542 2638 1546 2642
rect 3318 2638 3322 2642
rect 3390 2638 3394 2642
rect 4174 2638 4178 2642
rect 4190 2638 4194 2642
rect 4318 2638 4322 2642
rect 2238 2628 2242 2632
rect 286 2618 290 2622
rect 382 2618 386 2622
rect 494 2618 498 2622
rect 662 2618 666 2622
rect 1078 2618 1082 2622
rect 2286 2618 2290 2622
rect 2686 2618 2690 2622
rect 2902 2618 2906 2622
rect 3334 2618 3338 2622
rect 3902 2618 3906 2622
rect 3918 2618 3922 2622
rect 3974 2618 3978 2622
rect 4062 2618 4066 2622
rect 4102 2618 4106 2622
rect 4134 2618 4138 2622
rect 4182 2618 4186 2622
rect 4286 2618 4290 2622
rect 4342 2618 4346 2622
rect 4598 2618 4602 2622
rect 498 2603 502 2607
rect 505 2603 509 2607
rect 1522 2603 1526 2607
rect 1529 2603 1533 2607
rect 2546 2603 2550 2607
rect 2553 2603 2557 2607
rect 3570 2603 3574 2607
rect 3577 2603 3581 2607
rect 750 2588 754 2592
rect 1022 2588 1026 2592
rect 1222 2588 1226 2592
rect 1342 2588 1346 2592
rect 1446 2588 1450 2592
rect 1454 2588 1458 2592
rect 1566 2588 1570 2592
rect 1678 2588 1682 2592
rect 1782 2588 1786 2592
rect 1790 2588 1794 2592
rect 2238 2588 2242 2592
rect 2302 2588 2306 2592
rect 2982 2588 2986 2592
rect 3006 2588 3010 2592
rect 3150 2588 3154 2592
rect 3278 2588 3282 2592
rect 3918 2588 3922 2592
rect 4118 2588 4122 2592
rect 1134 2568 1138 2572
rect 1910 2568 1914 2572
rect 1926 2568 1930 2572
rect 2006 2568 2010 2572
rect 2110 2568 2114 2572
rect 2174 2568 2178 2572
rect 2198 2568 2202 2572
rect 2294 2568 2298 2572
rect 2758 2568 2762 2572
rect 2870 2568 2874 2572
rect 2950 2568 2954 2572
rect 3582 2568 3586 2572
rect 3838 2568 3842 2572
rect 54 2557 58 2561
rect 654 2558 658 2562
rect 814 2558 818 2562
rect 830 2558 834 2562
rect 902 2558 906 2562
rect 1958 2558 1962 2562
rect 2214 2558 2218 2562
rect 22 2548 26 2552
rect 70 2548 74 2552
rect 134 2548 138 2552
rect 190 2547 194 2551
rect 286 2548 290 2552
rect 294 2548 298 2552
rect 422 2548 426 2552
rect 502 2548 506 2552
rect 558 2548 562 2552
rect 582 2547 586 2551
rect 638 2548 642 2552
rect 686 2547 690 2551
rect 758 2548 762 2552
rect 790 2548 794 2552
rect 822 2548 826 2552
rect 846 2548 850 2552
rect 862 2548 866 2552
rect 878 2548 882 2552
rect 894 2548 898 2552
rect 910 2548 914 2552
rect 926 2548 930 2552
rect 958 2547 962 2551
rect 990 2548 994 2552
rect 1070 2547 1074 2551
rect 1102 2548 1106 2552
rect 1142 2548 1146 2552
rect 1406 2548 1410 2552
rect 1518 2547 1522 2551
rect 1598 2548 1602 2552
rect 1630 2547 1634 2551
rect 1662 2548 1666 2552
rect 1726 2548 1730 2552
rect 1854 2547 1858 2551
rect 1942 2548 1946 2552
rect 2086 2548 2090 2552
rect 2142 2548 2146 2552
rect 2422 2558 2426 2562
rect 2238 2548 2242 2552
rect 2358 2548 2362 2552
rect 2470 2558 2474 2562
rect 2590 2558 2594 2562
rect 2678 2558 2682 2562
rect 2854 2558 2858 2562
rect 2926 2558 2930 2562
rect 2390 2547 2394 2551
rect 2446 2548 2450 2552
rect 2470 2548 2474 2552
rect 2542 2547 2546 2551
rect 2606 2548 2610 2552
rect 2662 2548 2666 2552
rect 2750 2548 2754 2552
rect 2790 2548 2794 2552
rect 2822 2547 2826 2551
rect 2878 2548 2882 2552
rect 2910 2548 2914 2552
rect 3022 2558 3026 2562
rect 3166 2558 3170 2562
rect 3286 2558 3290 2562
rect 3310 2558 3314 2562
rect 3334 2558 3338 2562
rect 3454 2558 3458 2562
rect 3462 2558 3466 2562
rect 3494 2558 3498 2562
rect 3542 2558 3546 2562
rect 3638 2558 3642 2562
rect 3654 2558 3658 2562
rect 3766 2558 3770 2562
rect 3926 2558 3930 2562
rect 3958 2558 3962 2562
rect 4062 2558 4066 2562
rect 4158 2558 4162 2562
rect 4246 2558 4250 2562
rect 3006 2548 3010 2552
rect 3078 2548 3082 2552
rect 3110 2547 3114 2551
rect 3150 2548 3154 2552
rect 3198 2547 3202 2551
rect 3310 2548 3314 2552
rect 3334 2548 3338 2552
rect 78 2538 82 2542
rect 142 2538 146 2542
rect 318 2538 322 2542
rect 382 2538 386 2542
rect 398 2538 402 2542
rect 598 2538 602 2542
rect 630 2538 634 2542
rect 694 2538 698 2542
rect 782 2538 786 2542
rect 798 2538 802 2542
rect 814 2538 818 2542
rect 854 2538 858 2542
rect 870 2538 874 2542
rect 886 2538 890 2542
rect 926 2538 930 2542
rect 1030 2538 1034 2542
rect 1206 2538 1210 2542
rect 1278 2538 1282 2542
rect 1398 2538 1402 2542
rect 1534 2538 1538 2542
rect 1726 2538 1730 2542
rect 1838 2538 1842 2542
rect 1870 2538 1874 2542
rect 1886 2538 1890 2542
rect 1910 2538 1914 2542
rect 1934 2538 1938 2542
rect 1974 2538 1978 2542
rect 1982 2538 1986 2542
rect 2014 2538 2018 2542
rect 2094 2538 2098 2542
rect 2118 2538 2122 2542
rect 2150 2538 2154 2542
rect 2174 2538 2178 2542
rect 2198 2538 2202 2542
rect 2270 2538 2274 2542
rect 2318 2538 2322 2542
rect 2422 2538 2426 2542
rect 2446 2538 2450 2542
rect 2558 2538 2562 2542
rect 2686 2538 2690 2542
rect 2878 2538 2882 2542
rect 2934 2538 2938 2542
rect 2966 2538 2970 2542
rect 2974 2538 2978 2542
rect 2998 2538 3002 2542
rect 3126 2538 3130 2542
rect 3142 2538 3146 2542
rect 3182 2538 3186 2542
rect 3270 2538 3274 2542
rect 3294 2538 3298 2542
rect 3318 2538 3322 2542
rect 3366 2547 3370 2551
rect 3462 2548 3466 2552
rect 3486 2548 3490 2552
rect 3566 2548 3570 2552
rect 3606 2548 3610 2552
rect 3630 2548 3634 2552
rect 3742 2548 3746 2552
rect 3798 2548 3802 2552
rect 3854 2548 3858 2552
rect 3878 2548 3882 2552
rect 3910 2548 3914 2552
rect 3942 2548 3946 2552
rect 3990 2548 3994 2552
rect 4078 2548 4082 2552
rect 4134 2548 4138 2552
rect 4142 2548 4146 2552
rect 4166 2548 4170 2552
rect 4206 2548 4210 2552
rect 4326 2558 4330 2562
rect 4510 2558 4514 2562
rect 4558 2558 4562 2562
rect 4270 2548 4274 2552
rect 4278 2548 4282 2552
rect 4406 2548 4410 2552
rect 4550 2548 4554 2552
rect 3350 2538 3354 2542
rect 3438 2538 3442 2542
rect 3486 2538 3490 2542
rect 3518 2538 3522 2542
rect 3566 2538 3570 2542
rect 3678 2538 3682 2542
rect 3734 2538 3738 2542
rect 3782 2538 3786 2542
rect 3822 2538 3826 2542
rect 3854 2538 3858 2542
rect 3886 2538 3890 2542
rect 3934 2538 3938 2542
rect 3966 2538 3970 2542
rect 3982 2538 3986 2542
rect 4038 2538 4042 2542
rect 4086 2538 4090 2542
rect 4198 2538 4202 2542
rect 4230 2538 4234 2542
rect 4310 2538 4314 2542
rect 4326 2538 4330 2542
rect 4334 2538 4338 2542
rect 4382 2538 4386 2542
rect 4414 2538 4418 2542
rect 4438 2538 4442 2542
rect 4470 2538 4474 2542
rect 4486 2538 4490 2542
rect 4494 2538 4498 2542
rect 4526 2538 4530 2542
rect 4574 2538 4578 2542
rect 6 2528 10 2532
rect 22 2528 26 2532
rect 38 2528 42 2532
rect 78 2528 82 2532
rect 158 2528 162 2532
rect 190 2528 194 2532
rect 486 2528 490 2532
rect 550 2528 554 2532
rect 614 2528 618 2532
rect 654 2528 658 2532
rect 1974 2528 1978 2532
rect 2262 2528 2266 2532
rect 2294 2528 2298 2532
rect 2310 2528 2314 2532
rect 2358 2528 2362 2532
rect 2390 2528 2394 2532
rect 2510 2528 2514 2532
rect 2630 2528 2634 2532
rect 2638 2528 2642 2532
rect 142 2518 146 2522
rect 254 2518 258 2522
rect 270 2518 274 2522
rect 478 2518 482 2522
rect 622 2518 626 2522
rect 830 2518 834 2522
rect 1894 2518 1898 2522
rect 1926 2518 1930 2522
rect 1958 2518 1962 2522
rect 1990 2518 1994 2522
rect 2102 2518 2106 2522
rect 2166 2518 2170 2522
rect 2190 2518 2194 2522
rect 2278 2518 2282 2522
rect 2582 2518 2586 2522
rect 2678 2518 2682 2522
rect 2958 2528 2962 2532
rect 3078 2528 3082 2532
rect 3534 2528 3538 2532
rect 3598 2528 3602 2532
rect 3646 2528 3650 2532
rect 3694 2528 3698 2532
rect 3702 2528 3706 2532
rect 3742 2528 3746 2532
rect 3894 2528 3898 2532
rect 3966 2528 3970 2532
rect 4046 2528 4050 2532
rect 4190 2528 4194 2532
rect 4254 2528 4258 2532
rect 4302 2528 4306 2532
rect 4350 2528 4354 2532
rect 4390 2528 4394 2532
rect 4406 2528 4410 2532
rect 4454 2528 4458 2532
rect 4462 2528 4466 2532
rect 2926 2518 2930 2522
rect 2942 2518 2946 2522
rect 3262 2518 3266 2522
rect 3430 2518 3434 2522
rect 3750 2518 3754 2522
rect 3814 2518 3818 2522
rect 3862 2518 3866 2522
rect 3974 2518 3978 2522
rect 4014 2518 4018 2522
rect 4182 2518 4186 2522
rect 4222 2518 4226 2522
rect 4342 2518 4346 2522
rect 4358 2518 4362 2522
rect 4366 2518 4370 2522
rect 4446 2518 4450 2522
rect 4526 2518 4530 2522
rect 2630 2508 2634 2512
rect 2638 2508 2642 2512
rect 1002 2503 1006 2507
rect 1009 2503 1013 2507
rect 2026 2503 2030 2507
rect 2033 2503 2037 2507
rect 3050 2503 3054 2507
rect 3057 2503 3061 2507
rect 4082 2503 4086 2507
rect 4089 2503 4093 2507
rect 1974 2498 1978 2502
rect 2182 2498 2186 2502
rect 2822 2498 2826 2502
rect 2934 2498 2938 2502
rect 2998 2498 3002 2502
rect 526 2488 530 2492
rect 638 2488 642 2492
rect 758 2488 762 2492
rect 1358 2488 1362 2492
rect 1454 2488 1458 2492
rect 1646 2488 1650 2492
rect 1742 2488 1746 2492
rect 1838 2488 1842 2492
rect 2030 2488 2034 2492
rect 2054 2488 2058 2492
rect 2358 2488 2362 2492
rect 2750 2488 2754 2492
rect 3022 2488 3026 2492
rect 3038 2488 3042 2492
rect 3166 2488 3170 2492
rect 3198 2488 3202 2492
rect 3382 2488 3386 2492
rect 3478 2488 3482 2492
rect 3598 2488 3602 2492
rect 3718 2488 3722 2492
rect 3742 2488 3746 2492
rect 4094 2488 4098 2492
rect 4166 2488 4170 2492
rect 4278 2488 4282 2492
rect 6 2478 10 2482
rect 78 2478 82 2482
rect 342 2478 346 2482
rect 374 2478 378 2482
rect 478 2478 482 2482
rect 518 2478 522 2482
rect 574 2478 578 2482
rect 614 2478 618 2482
rect 694 2478 698 2482
rect 982 2478 986 2482
rect 1038 2478 1042 2482
rect 1078 2478 1082 2482
rect 1094 2478 1098 2482
rect 1102 2478 1106 2482
rect 1110 2478 1114 2482
rect 1150 2478 1154 2482
rect 1262 2478 1266 2482
rect 1518 2478 1522 2482
rect 1974 2478 1978 2482
rect 2038 2478 2042 2482
rect 2182 2478 2186 2482
rect 2294 2478 2298 2482
rect 2390 2478 2394 2482
rect 2670 2478 2674 2482
rect 2774 2478 2778 2482
rect 2822 2478 2826 2482
rect 2854 2478 2858 2482
rect 2926 2478 2930 2482
rect 2934 2478 2938 2482
rect 2982 2478 2986 2482
rect 2998 2478 3002 2482
rect 3102 2478 3106 2482
rect 3222 2478 3226 2482
rect 3238 2478 3242 2482
rect 3254 2478 3258 2482
rect 3406 2478 3410 2482
rect 3486 2478 3490 2482
rect 3558 2478 3562 2482
rect 3566 2478 3570 2482
rect 3622 2478 3626 2482
rect 3630 2478 3634 2482
rect 3686 2478 3690 2482
rect 3750 2478 3754 2482
rect 3830 2478 3834 2482
rect 3886 2478 3890 2482
rect 3902 2478 3906 2482
rect 3942 2478 3946 2482
rect 4078 2478 4082 2482
rect 4110 2478 4114 2482
rect 4134 2478 4138 2482
rect 4174 2478 4178 2482
rect 4254 2478 4258 2482
rect 4278 2478 4282 2482
rect 4518 2478 4522 2482
rect 4542 2478 4546 2482
rect 4582 2478 4586 2482
rect 22 2468 26 2472
rect 62 2468 66 2472
rect 110 2468 114 2472
rect 190 2468 194 2472
rect 326 2468 330 2472
rect 406 2468 410 2472
rect 582 2468 586 2472
rect 622 2468 626 2472
rect 830 2468 834 2472
rect 846 2468 850 2472
rect 862 2468 866 2472
rect 886 2468 890 2472
rect 902 2468 906 2472
rect 918 2468 922 2472
rect 942 2468 946 2472
rect 982 2468 986 2472
rect 1006 2468 1010 2472
rect 1070 2468 1074 2472
rect 1086 2468 1090 2472
rect 1118 2468 1122 2472
rect 1190 2468 1194 2472
rect 1302 2468 1306 2472
rect 1374 2468 1378 2472
rect 1470 2468 1474 2472
rect 1574 2468 1578 2472
rect 2126 2468 2130 2472
rect 2142 2468 2146 2472
rect 2182 2468 2186 2472
rect 2462 2468 2466 2472
rect 2510 2468 2514 2472
rect 2518 2468 2522 2472
rect 2582 2468 2586 2472
rect 2590 2468 2594 2472
rect 2638 2468 2642 2472
rect 2726 2468 2730 2472
rect 2758 2468 2762 2472
rect 2910 2468 2914 2472
rect 2934 2468 2938 2472
rect 2966 2468 2970 2472
rect 3006 2468 3010 2472
rect 3054 2468 3058 2472
rect 3078 2468 3082 2472
rect 3126 2468 3130 2472
rect 3182 2468 3186 2472
rect 3190 2468 3194 2472
rect 3286 2468 3290 2472
rect 3294 2468 3298 2472
rect 3318 2468 3322 2472
rect 3342 2468 3346 2472
rect 3438 2468 3442 2472
rect 3470 2468 3474 2472
rect 3518 2468 3522 2472
rect 3550 2468 3554 2472
rect 3590 2468 3594 2472
rect 3646 2468 3650 2472
rect 3662 2468 3666 2472
rect 3694 2468 3698 2472
rect 3726 2468 3730 2472
rect 3766 2468 3770 2472
rect 3782 2468 3786 2472
rect 3838 2468 3842 2472
rect 3862 2468 3866 2472
rect 3942 2468 3946 2472
rect 3990 2468 3994 2472
rect 4054 2468 4058 2472
rect 4142 2468 4146 2472
rect 4198 2468 4202 2472
rect 4214 2468 4218 2472
rect 4230 2468 4234 2472
rect 4262 2468 4266 2472
rect 4326 2468 4330 2472
rect 4342 2468 4346 2472
rect 4358 2468 4362 2472
rect 4390 2468 4394 2472
rect 4438 2468 4442 2472
rect 4446 2468 4450 2472
rect 4574 2468 4578 2472
rect 54 2458 58 2462
rect 118 2458 122 2462
rect 206 2459 210 2463
rect 342 2458 346 2462
rect 414 2458 418 2462
rect 478 2458 482 2462
rect 510 2458 514 2462
rect 630 2458 634 2462
rect 694 2459 698 2463
rect 726 2458 730 2462
rect 766 2458 770 2462
rect 838 2458 842 2462
rect 870 2458 874 2462
rect 878 2458 882 2462
rect 910 2458 914 2462
rect 934 2458 938 2462
rect 1046 2458 1050 2462
rect 1126 2458 1130 2462
rect 1142 2458 1146 2462
rect 1182 2459 1186 2463
rect 1294 2459 1298 2463
rect 1390 2459 1394 2463
rect 1502 2458 1506 2462
rect 1638 2458 1642 2462
rect 1678 2458 1682 2462
rect 1686 2458 1690 2462
rect 1774 2458 1778 2462
rect 1806 2459 1810 2463
rect 1870 2458 1874 2462
rect 1902 2459 1906 2463
rect 1942 2458 1946 2462
rect 1950 2458 1954 2462
rect 1998 2458 2002 2462
rect 2078 2458 2082 2462
rect 2110 2459 2114 2463
rect 2150 2458 2154 2462
rect 2182 2458 2186 2462
rect 2206 2458 2210 2462
rect 2262 2458 2266 2462
rect 2302 2458 2306 2462
rect 2390 2459 2394 2463
rect 2502 2458 2506 2462
rect 2574 2458 2578 2462
rect 2638 2458 2642 2462
rect 2678 2458 2682 2462
rect 2790 2458 2794 2462
rect 2798 2458 2802 2462
rect 2854 2459 2858 2463
rect 2958 2458 2962 2462
rect 2966 2458 2970 2462
rect 2982 2458 2986 2462
rect 3126 2458 3130 2462
rect 3262 2458 3266 2462
rect 3366 2458 3370 2462
rect 3430 2458 3434 2462
rect 3462 2458 3466 2462
rect 3510 2458 3514 2462
rect 3526 2458 3530 2462
rect 3646 2458 3650 2462
rect 3670 2458 3674 2462
rect 3702 2458 3706 2462
rect 3790 2458 3794 2462
rect 3814 2458 3818 2462
rect 3918 2458 3922 2462
rect 3958 2458 3962 2462
rect 3974 2458 3978 2462
rect 4006 2458 4010 2462
rect 4062 2458 4066 2462
rect 4078 2458 4082 2462
rect 4118 2458 4122 2462
rect 4150 2458 4154 2462
rect 4190 2458 4194 2462
rect 4198 2458 4202 2462
rect 4222 2458 4226 2462
rect 4238 2458 4242 2462
rect 4254 2458 4258 2462
rect 4286 2458 4290 2462
rect 4334 2458 4338 2462
rect 4350 2458 4354 2462
rect 4430 2458 4434 2462
rect 4454 2458 4458 2462
rect 4486 2458 4490 2462
rect 38 2449 42 2453
rect 902 2448 906 2452
rect 918 2448 922 2452
rect 974 2448 978 2452
rect 1934 2448 1938 2452
rect 1982 2448 1986 2452
rect 2166 2448 2170 2452
rect 2190 2448 2194 2452
rect 2246 2448 2250 2452
rect 2478 2448 2482 2452
rect 2534 2448 2538 2452
rect 2606 2448 2610 2452
rect 2742 2448 2746 2452
rect 2758 2448 2762 2452
rect 2782 2448 2786 2452
rect 2942 2448 2946 2452
rect 3030 2448 3034 2452
rect 3166 2448 3170 2452
rect 3206 2448 3210 2452
rect 3310 2448 3314 2452
rect 3334 2448 3338 2452
rect 3342 2448 3346 2452
rect 3358 2448 3362 2452
rect 3414 2448 3418 2452
rect 3446 2448 3450 2452
rect 3494 2448 3498 2452
rect 3662 2448 3666 2452
rect 3718 2448 3722 2452
rect 3742 2448 3746 2452
rect 3782 2448 3786 2452
rect 3798 2448 3802 2452
rect 3854 2448 3858 2452
rect 3910 2448 3914 2452
rect 3966 2448 3970 2452
rect 3998 2448 4002 2452
rect 4030 2448 4034 2452
rect 4350 2448 4354 2452
rect 4406 2448 4410 2452
rect 4414 2448 4418 2452
rect 4478 2448 4482 2452
rect 982 2438 986 2442
rect 1246 2438 1250 2442
rect 3222 2438 3226 2442
rect 3318 2438 3322 2442
rect 3926 2438 3930 2442
rect 3982 2438 3986 2442
rect 4014 2438 4018 2442
rect 4190 2438 4194 2442
rect 4366 2438 4370 2442
rect 270 2428 274 2432
rect 3302 2428 3306 2432
rect 4486 2428 4490 2432
rect 174 2418 178 2422
rect 598 2418 602 2422
rect 758 2418 762 2422
rect 862 2418 866 2422
rect 998 2418 1002 2422
rect 1030 2418 1034 2422
rect 1062 2418 1066 2422
rect 1254 2418 1258 2422
rect 1550 2418 1554 2422
rect 1998 2418 2002 2422
rect 2150 2418 2154 2422
rect 2454 2418 2458 2422
rect 3230 2418 3234 2422
rect 3246 2418 3250 2422
rect 3398 2418 3402 2422
rect 3918 2418 3922 2422
rect 4006 2418 4010 2422
rect 4046 2418 4050 2422
rect 4118 2418 4122 2422
rect 4430 2418 4434 2422
rect 4566 2418 4570 2422
rect 4590 2418 4594 2422
rect 498 2403 502 2407
rect 505 2403 509 2407
rect 1522 2403 1526 2407
rect 1529 2403 1533 2407
rect 2546 2403 2550 2407
rect 2553 2403 2557 2407
rect 3570 2403 3574 2407
rect 3577 2403 3581 2407
rect 342 2388 346 2392
rect 478 2388 482 2392
rect 558 2388 562 2392
rect 862 2388 866 2392
rect 1126 2388 1130 2392
rect 1222 2388 1226 2392
rect 1542 2388 1546 2392
rect 1662 2388 1666 2392
rect 1758 2388 1762 2392
rect 3142 2388 3146 2392
rect 3342 2388 3346 2392
rect 3358 2388 3362 2392
rect 3926 2388 3930 2392
rect 4214 2388 4218 2392
rect 4318 2388 4322 2392
rect 46 2378 50 2382
rect 3542 2378 3546 2382
rect 3630 2378 3634 2382
rect 3870 2378 3874 2382
rect 326 2368 330 2372
rect 990 2368 994 2372
rect 1302 2368 1306 2372
rect 1318 2368 1322 2372
rect 1398 2368 1402 2372
rect 1414 2368 1418 2372
rect 1654 2368 1658 2372
rect 2918 2368 2922 2372
rect 3486 2368 3490 2372
rect 3878 2368 3882 2372
rect 4222 2368 4226 2372
rect 4270 2368 4274 2372
rect 4326 2368 4330 2372
rect 4518 2368 4522 2372
rect 4542 2368 4546 2372
rect 726 2358 730 2362
rect 926 2358 930 2362
rect 1950 2358 1954 2362
rect 1966 2358 1970 2362
rect 2110 2358 2114 2362
rect 2158 2358 2162 2362
rect 2246 2358 2250 2362
rect 2254 2358 2258 2362
rect 2302 2358 2306 2362
rect 2326 2358 2330 2362
rect 2374 2358 2378 2362
rect 2414 2358 2418 2362
rect 142 2348 146 2352
rect 206 2348 210 2352
rect 270 2348 274 2352
rect 358 2348 362 2352
rect 398 2348 402 2352
rect 462 2348 466 2352
rect 510 2348 514 2352
rect 614 2348 618 2352
rect 654 2348 658 2352
rect 678 2348 682 2352
rect 718 2348 722 2352
rect 742 2348 746 2352
rect 798 2347 802 2351
rect 902 2348 906 2352
rect 958 2348 962 2352
rect 966 2348 970 2352
rect 998 2348 1002 2352
rect 1014 2348 1018 2352
rect 1062 2347 1066 2351
rect 1094 2348 1098 2352
rect 1158 2347 1162 2351
rect 1190 2348 1194 2352
rect 1254 2347 1258 2351
rect 1358 2348 1362 2352
rect 1382 2348 1386 2352
rect 1422 2348 1426 2352
rect 1478 2347 1482 2351
rect 1486 2348 1490 2352
rect 1510 2348 1514 2352
rect 1606 2348 1610 2352
rect 1694 2348 1698 2352
rect 1702 2348 1706 2352
rect 1790 2348 1794 2352
rect 1822 2347 1826 2351
rect 1918 2347 1922 2351
rect 1974 2348 1978 2352
rect 2078 2347 2082 2351
rect 2110 2348 2114 2352
rect 2126 2348 2130 2352
rect 2174 2348 2178 2352
rect 2222 2348 2226 2352
rect 2398 2348 2402 2352
rect 2710 2358 2714 2362
rect 2758 2358 2762 2362
rect 2470 2348 2474 2352
rect 2582 2347 2586 2351
rect 2654 2348 2658 2352
rect 2678 2347 2682 2351
rect 2734 2348 2738 2352
rect 2750 2348 2754 2352
rect 30 2338 34 2342
rect 118 2338 122 2342
rect 150 2338 154 2342
rect 214 2338 218 2342
rect 262 2338 266 2342
rect 390 2338 394 2342
rect 534 2338 538 2342
rect 734 2338 738 2342
rect 782 2338 786 2342
rect 926 2338 930 2342
rect 1006 2338 1010 2342
rect 1142 2338 1146 2342
rect 1262 2338 1266 2342
rect 1446 2338 1450 2342
rect 1550 2338 1554 2342
rect 1726 2338 1730 2342
rect 2070 2338 2074 2342
rect 2278 2338 2282 2342
rect 2318 2338 2322 2342
rect 2342 2338 2346 2342
rect 2398 2338 2402 2342
rect 2446 2338 2450 2342
rect 2494 2338 2498 2342
rect 2510 2338 2514 2342
rect 2534 2338 2538 2342
rect 2566 2338 2570 2342
rect 2598 2338 2602 2342
rect 2750 2338 2754 2342
rect 2782 2358 2786 2362
rect 2814 2358 2818 2362
rect 2854 2358 2858 2362
rect 2894 2358 2898 2362
rect 2926 2358 2930 2362
rect 2958 2358 2962 2362
rect 3062 2358 3066 2362
rect 3134 2358 3138 2362
rect 2830 2348 2834 2352
rect 2870 2348 2874 2352
rect 2894 2348 2898 2352
rect 2950 2348 2954 2352
rect 2974 2348 2978 2352
rect 2990 2348 2994 2352
rect 3038 2348 3042 2352
rect 3086 2348 3090 2352
rect 3158 2348 3162 2352
rect 3198 2358 3202 2362
rect 3214 2358 3218 2362
rect 3238 2358 3242 2362
rect 3302 2358 3306 2362
rect 3406 2358 3410 2362
rect 3470 2358 3474 2362
rect 3526 2358 3530 2362
rect 3558 2358 3562 2362
rect 3638 2358 3642 2362
rect 3670 2358 3674 2362
rect 3718 2358 3722 2362
rect 3774 2358 3778 2362
rect 3830 2358 3834 2362
rect 3862 2358 3866 2362
rect 3910 2358 3914 2362
rect 3958 2358 3962 2362
rect 3974 2358 3978 2362
rect 4062 2358 4066 2362
rect 4142 2358 4146 2362
rect 4182 2358 4186 2362
rect 4206 2358 4210 2362
rect 4238 2358 4242 2362
rect 4342 2358 4346 2362
rect 4358 2358 4362 2362
rect 4374 2358 4378 2362
rect 4430 2358 4434 2362
rect 4462 2358 4466 2362
rect 4502 2358 4506 2362
rect 3254 2348 3258 2352
rect 3302 2348 3306 2352
rect 3374 2348 3378 2352
rect 3478 2348 3482 2352
rect 3510 2348 3514 2352
rect 3526 2348 3530 2352
rect 3542 2348 3546 2352
rect 3614 2348 3618 2352
rect 3654 2348 3658 2352
rect 3686 2348 3690 2352
rect 3694 2348 3698 2352
rect 3750 2348 3754 2352
rect 3766 2348 3770 2352
rect 3806 2348 3810 2352
rect 3822 2348 3826 2352
rect 3846 2348 3850 2352
rect 3870 2348 3874 2352
rect 3918 2348 3922 2352
rect 4014 2348 4018 2352
rect 4046 2348 4050 2352
rect 4126 2348 4130 2352
rect 4230 2348 4234 2352
rect 4270 2348 4274 2352
rect 4294 2348 4298 2352
rect 4334 2348 4338 2352
rect 4358 2348 4362 2352
rect 4406 2348 4410 2352
rect 4430 2348 4434 2352
rect 4518 2348 4522 2352
rect 4542 2348 4546 2352
rect 4582 2348 4586 2352
rect 2798 2338 2802 2342
rect 2838 2338 2842 2342
rect 2878 2338 2882 2342
rect 2918 2338 2922 2342
rect 2950 2338 2954 2342
rect 2982 2338 2986 2342
rect 3014 2338 3018 2342
rect 3030 2338 3034 2342
rect 3046 2338 3050 2342
rect 3094 2338 3098 2342
rect 3102 2338 3106 2342
rect 3118 2338 3122 2342
rect 3206 2338 3210 2342
rect 3230 2338 3234 2342
rect 3262 2338 3266 2342
rect 3310 2338 3314 2342
rect 3318 2340 3322 2344
rect 3350 2338 3354 2342
rect 3382 2338 3386 2342
rect 3430 2338 3434 2342
rect 3454 2338 3458 2342
rect 3502 2338 3506 2342
rect 3534 2338 3538 2342
rect 3614 2338 3618 2342
rect 3662 2338 3666 2342
rect 3686 2338 3690 2342
rect 3734 2338 3738 2342
rect 3790 2338 3794 2342
rect 3814 2338 3818 2342
rect 3822 2338 3826 2342
rect 3854 2338 3858 2342
rect 3894 2338 3898 2342
rect 3942 2338 3946 2342
rect 3974 2338 3978 2342
rect 3998 2338 4002 2342
rect 4030 2338 4034 2342
rect 4046 2338 4050 2342
rect 4142 2338 4146 2342
rect 4150 2338 4154 2342
rect 4158 2338 4162 2342
rect 4166 2338 4170 2342
rect 4190 2338 4194 2342
rect 4246 2338 4250 2342
rect 4262 2338 4266 2342
rect 4350 2338 4354 2342
rect 4398 2338 4402 2342
rect 4414 2338 4418 2342
rect 4526 2338 4530 2342
rect 4534 2338 4538 2342
rect 6 2328 10 2332
rect 14 2328 18 2332
rect 22 2328 26 2332
rect 174 2328 178 2332
rect 214 2328 218 2332
rect 574 2328 578 2332
rect 606 2328 610 2332
rect 766 2328 770 2332
rect 798 2328 802 2332
rect 870 2328 874 2332
rect 878 2328 882 2332
rect 886 2328 890 2332
rect 934 2328 938 2332
rect 950 2328 954 2332
rect 974 2328 978 2332
rect 990 2328 994 2332
rect 1886 2328 1890 2332
rect 1918 2328 1922 2332
rect 1990 2328 1994 2332
rect 2150 2328 2154 2332
rect 2198 2328 2202 2332
rect 2206 2328 2210 2332
rect 2294 2328 2298 2332
rect 2358 2328 2362 2332
rect 2462 2328 2466 2332
rect 2646 2328 2650 2332
rect 3006 2328 3010 2332
rect 3102 2328 3106 2332
rect 3150 2328 3154 2332
rect 3174 2328 3178 2332
rect 3278 2328 3282 2332
rect 3366 2328 3370 2332
rect 3398 2328 3402 2332
rect 3438 2328 3442 2332
rect 3582 2328 3586 2332
rect 3694 2328 3698 2332
rect 3782 2328 3786 2332
rect 3798 2328 3802 2332
rect 4006 2328 4010 2332
rect 4014 2328 4018 2332
rect 4310 2328 4314 2332
rect 4382 2328 4386 2332
rect 4422 2328 4426 2332
rect 4454 2328 4458 2332
rect 4494 2328 4498 2332
rect 4566 2328 4570 2332
rect 150 2318 154 2322
rect 214 2318 218 2322
rect 454 2318 458 2322
rect 478 2318 482 2322
rect 606 2318 610 2322
rect 942 2318 946 2322
rect 1438 2318 1442 2322
rect 1998 2318 2002 2322
rect 2158 2318 2162 2322
rect 2246 2318 2250 2322
rect 2302 2318 2306 2322
rect 2334 2318 2338 2322
rect 2350 2318 2354 2322
rect 2710 2318 2714 2322
rect 2742 2318 2746 2322
rect 2806 2318 2810 2322
rect 3134 2318 3138 2322
rect 3214 2318 3218 2322
rect 3238 2318 3242 2322
rect 3334 2318 3338 2322
rect 3390 2318 3394 2322
rect 3486 2318 3490 2322
rect 3638 2318 3642 2322
rect 4078 2318 4082 2322
rect 4182 2318 4186 2322
rect 4198 2318 4202 2322
rect 4254 2318 4258 2322
rect 4390 2318 4394 2322
rect 4446 2318 4450 2322
rect 4462 2318 4466 2322
rect 1990 2308 1994 2312
rect 2150 2308 2154 2312
rect 2198 2308 2202 2312
rect 2206 2308 2210 2312
rect 1002 2303 1006 2307
rect 1009 2303 1013 2307
rect 2026 2303 2030 2307
rect 2033 2303 2037 2307
rect 3050 2303 3054 2307
rect 3057 2303 3061 2307
rect 4082 2303 4086 2307
rect 4089 2303 4093 2307
rect 302 2288 306 2292
rect 326 2288 330 2292
rect 958 2288 962 2292
rect 1262 2288 1266 2292
rect 1366 2288 1370 2292
rect 1646 2288 1650 2292
rect 1750 2288 1754 2292
rect 1846 2288 1850 2292
rect 1950 2288 1954 2292
rect 2230 2288 2234 2292
rect 2390 2288 2394 2292
rect 2766 2288 2770 2292
rect 2854 2288 2858 2292
rect 3038 2288 3042 2292
rect 3246 2288 3250 2292
rect 3302 2288 3306 2292
rect 3374 2288 3378 2292
rect 3454 2288 3458 2292
rect 3478 2288 3482 2292
rect 3622 2288 3626 2292
rect 3686 2288 3690 2292
rect 3862 2288 3866 2292
rect 4214 2288 4218 2292
rect 4302 2288 4306 2292
rect 4494 2288 4498 2292
rect 94 2278 98 2282
rect 126 2278 130 2282
rect 174 2278 178 2282
rect 198 2278 202 2282
rect 230 2278 234 2282
rect 558 2278 562 2282
rect 582 2278 586 2282
rect 686 2278 690 2282
rect 750 2278 754 2282
rect 886 2278 890 2282
rect 894 2278 898 2282
rect 902 2278 906 2282
rect 974 2278 978 2282
rect 982 2278 986 2282
rect 998 2278 1002 2282
rect 1086 2278 1090 2282
rect 1102 2278 1106 2282
rect 1470 2278 1474 2282
rect 1918 2278 1922 2282
rect 2262 2278 2266 2282
rect 2382 2278 2386 2282
rect 2398 2278 2402 2282
rect 2534 2278 2538 2282
rect 2630 2278 2634 2282
rect 2654 2278 2658 2282
rect 2750 2278 2754 2282
rect 2822 2278 2826 2282
rect 2886 2278 2890 2282
rect 2990 2278 2994 2282
rect 3062 2278 3066 2282
rect 142 2268 146 2272
rect 166 2268 170 2272
rect 182 2268 186 2272
rect 318 2268 322 2272
rect 350 2268 354 2272
rect 382 2268 386 2272
rect 454 2268 458 2272
rect 470 2268 474 2272
rect 702 2268 706 2272
rect 726 2268 730 2272
rect 742 2268 746 2272
rect 798 2268 802 2272
rect 918 2268 922 2272
rect 958 2268 962 2272
rect 1030 2268 1034 2272
rect 1142 2268 1146 2272
rect 1206 2268 1210 2272
rect 1318 2268 1322 2272
rect 1382 2268 1386 2272
rect 1486 2268 1490 2272
rect 1550 2268 1554 2272
rect 1582 2268 1586 2272
rect 1590 2268 1594 2272
rect 1670 2268 1674 2272
rect 1790 2268 1794 2272
rect 2030 2268 2034 2272
rect 2070 2268 2074 2272
rect 2158 2268 2162 2272
rect 2206 2268 2210 2272
rect 2214 2268 2218 2272
rect 2238 2268 2242 2272
rect 2278 2268 2282 2272
rect 94 2259 98 2263
rect 190 2258 194 2262
rect 230 2259 234 2263
rect 342 2258 346 2262
rect 358 2258 362 2262
rect 390 2258 394 2262
rect 486 2258 490 2262
rect 542 2258 546 2262
rect 614 2259 618 2263
rect 646 2258 650 2262
rect 686 2258 690 2262
rect 734 2258 738 2262
rect 790 2259 794 2263
rect 878 2258 882 2262
rect 950 2258 954 2262
rect 1038 2258 1042 2262
rect 1134 2259 1138 2263
rect 1310 2258 1314 2262
rect 1398 2259 1402 2263
rect 1686 2259 1690 2263
rect 1798 2258 1802 2262
rect 1886 2258 1890 2262
rect 1918 2259 1922 2263
rect 1982 2258 1986 2262
rect 2014 2259 2018 2263
rect 2366 2268 2370 2272
rect 2518 2268 2522 2272
rect 2614 2268 2618 2272
rect 2630 2268 2634 2272
rect 2662 2268 2666 2272
rect 2686 2268 2690 2272
rect 2734 2268 2738 2272
rect 2758 2268 2762 2272
rect 2782 2268 2786 2272
rect 2862 2268 2866 2272
rect 2894 2268 2898 2272
rect 2918 2268 2922 2272
rect 2998 2268 3002 2272
rect 3014 2268 3018 2272
rect 3070 2268 3074 2272
rect 3214 2278 3218 2282
rect 3254 2278 3258 2282
rect 3278 2278 3282 2282
rect 3294 2278 3298 2282
rect 3406 2278 3410 2282
rect 3438 2278 3442 2282
rect 3446 2278 3450 2282
rect 3550 2278 3554 2282
rect 3574 2278 3578 2282
rect 3590 2278 3594 2282
rect 3670 2278 3674 2282
rect 3102 2268 3106 2272
rect 3150 2268 3154 2272
rect 3166 2268 3170 2272
rect 3198 2268 3202 2272
rect 3294 2268 3298 2272
rect 3310 2268 3314 2272
rect 3358 2268 3362 2272
rect 3390 2268 3394 2272
rect 3462 2268 3466 2272
rect 3494 2266 3498 2270
rect 3502 2268 3506 2272
rect 3510 2268 3514 2272
rect 3526 2268 3530 2272
rect 3550 2268 3554 2272
rect 3606 2268 3610 2272
rect 3646 2268 3650 2272
rect 3702 2278 3706 2282
rect 3750 2278 3754 2282
rect 3790 2278 3794 2282
rect 3798 2278 3802 2282
rect 3814 2278 3818 2282
rect 3830 2278 3834 2282
rect 3838 2278 3842 2282
rect 3878 2278 3882 2282
rect 3910 2278 3914 2282
rect 3726 2268 3730 2272
rect 3742 2268 3746 2272
rect 3758 2268 3762 2272
rect 3974 2278 3978 2282
rect 4006 2278 4010 2282
rect 4110 2278 4114 2282
rect 4246 2278 4250 2282
rect 4262 2278 4266 2282
rect 4270 2278 4274 2282
rect 4374 2278 4378 2282
rect 4398 2278 4402 2282
rect 4470 2278 4474 2282
rect 3934 2268 3938 2272
rect 3966 2268 3970 2272
rect 4022 2268 4026 2272
rect 4086 2268 4090 2272
rect 4118 2268 4122 2272
rect 4246 2268 4250 2272
rect 4286 2268 4290 2272
rect 4326 2268 4330 2272
rect 4334 2268 4338 2272
rect 4350 2268 4354 2272
rect 4406 2268 4410 2272
rect 4462 2268 4466 2272
rect 4478 2268 4482 2272
rect 4582 2268 4586 2272
rect 2094 2258 2098 2262
rect 2198 2258 2202 2262
rect 2326 2258 2330 2262
rect 2334 2258 2338 2262
rect 2406 2258 2410 2262
rect 2502 2259 2506 2263
rect 2574 2258 2578 2262
rect 2590 2258 2594 2262
rect 2614 2258 2618 2262
rect 2638 2258 2642 2262
rect 2806 2258 2810 2262
rect 2822 2258 2826 2262
rect 2870 2258 2874 2262
rect 2886 2258 2890 2262
rect 2926 2258 2930 2262
rect 2950 2258 2954 2262
rect 2982 2258 2986 2262
rect 3022 2258 3026 2262
rect 3046 2258 3050 2262
rect 3126 2258 3130 2262
rect 3142 2258 3146 2262
rect 3158 2258 3162 2262
rect 3190 2258 3194 2262
rect 3230 2258 3234 2262
rect 3318 2258 3322 2262
rect 3334 2258 3338 2262
rect 3382 2258 3386 2262
rect 3422 2258 3426 2262
rect 3470 2258 3474 2262
rect 3534 2258 3538 2262
rect 3606 2258 3610 2262
rect 3654 2258 3658 2262
rect 3694 2258 3698 2262
rect 3734 2258 3738 2262
rect 3774 2258 3778 2262
rect 3814 2258 3818 2262
rect 3894 2258 3898 2262
rect 3910 2258 3914 2262
rect 3974 2258 3978 2262
rect 4038 2258 4042 2262
rect 4070 2258 4074 2262
rect 4078 2258 4082 2262
rect 4110 2258 4114 2262
rect 4134 2258 4138 2262
rect 4166 2258 4170 2262
rect 4198 2258 4202 2262
rect 4262 2258 4266 2262
rect 4294 2258 4298 2262
rect 4318 2258 4322 2262
rect 4390 2258 4394 2262
rect 4414 2258 4418 2262
rect 4438 2258 4442 2262
rect 4454 2258 4458 2262
rect 4502 2258 4506 2262
rect 4526 2258 4530 2262
rect 4574 2258 4578 2262
rect 302 2248 306 2252
rect 1070 2248 1074 2252
rect 2174 2248 2178 2252
rect 2230 2248 2234 2252
rect 2238 2248 2242 2252
rect 2254 2248 2258 2252
rect 2302 2248 2306 2252
rect 2310 2248 2314 2252
rect 2342 2248 2346 2252
rect 2598 2248 2602 2252
rect 2678 2248 2682 2252
rect 2702 2248 2706 2252
rect 2774 2248 2778 2252
rect 2782 2248 2786 2252
rect 2886 2248 2890 2252
rect 2942 2248 2946 2252
rect 3102 2248 3106 2252
rect 3118 2248 3122 2252
rect 3166 2248 3170 2252
rect 3182 2248 3186 2252
rect 3254 2248 3258 2252
rect 3270 2248 3274 2252
rect 3326 2248 3330 2252
rect 3358 2248 3362 2252
rect 3374 2248 3378 2252
rect 3438 2248 3442 2252
rect 3566 2248 3570 2252
rect 3630 2248 3634 2252
rect 3950 2248 3954 2252
rect 4030 2248 4034 2252
rect 4062 2248 4066 2252
rect 4126 2248 4130 2252
rect 4158 2248 4162 2252
rect 4190 2248 4194 2252
rect 4262 2248 4266 2252
rect 4350 2248 4354 2252
rect 4502 2248 4506 2252
rect 6 2238 10 2242
rect 1198 2238 1202 2242
rect 2814 2238 2818 2242
rect 2958 2238 2962 2242
rect 3342 2238 3346 2242
rect 4014 2238 4018 2242
rect 4046 2238 4050 2242
rect 4142 2238 4146 2242
rect 4174 2238 4178 2242
rect 4206 2238 4210 2242
rect 4222 2238 4226 2242
rect 4494 2238 4498 2242
rect 4510 2238 4514 2242
rect 4550 2248 4554 2252
rect 4534 2238 4538 2242
rect 4566 2238 4570 2242
rect 294 2228 298 2232
rect 2150 2228 2154 2232
rect 3814 2228 3818 2232
rect 4342 2228 4346 2232
rect 4526 2228 4530 2232
rect 518 2218 522 2222
rect 878 2218 882 2222
rect 990 2218 994 2222
rect 1078 2218 1082 2222
rect 1094 2218 1098 2222
rect 1462 2218 1466 2222
rect 1478 2218 1482 2222
rect 1558 2218 1562 2222
rect 1854 2218 1858 2222
rect 2422 2218 2426 2222
rect 2438 2218 2442 2222
rect 2606 2218 2610 2222
rect 2670 2218 2674 2222
rect 3262 2218 3266 2222
rect 3334 2218 3338 2222
rect 4038 2218 4042 2222
rect 4134 2218 4138 2222
rect 4166 2218 4170 2222
rect 498 2203 502 2207
rect 505 2203 509 2207
rect 1522 2203 1526 2207
rect 1529 2203 1533 2207
rect 2546 2203 2550 2207
rect 2553 2203 2557 2207
rect 3570 2203 3574 2207
rect 3577 2203 3581 2207
rect 30 2188 34 2192
rect 54 2188 58 2192
rect 78 2188 82 2192
rect 1062 2188 1066 2192
rect 2758 2188 2762 2192
rect 2902 2188 2906 2192
rect 3182 2188 3186 2192
rect 3230 2188 3234 2192
rect 3446 2188 3450 2192
rect 3750 2188 3754 2192
rect 3870 2188 3874 2192
rect 4006 2188 4010 2192
rect 4014 2188 4018 2192
rect 4302 2188 4306 2192
rect 4326 2188 4330 2192
rect 4350 2188 4354 2192
rect 4406 2188 4410 2192
rect 4478 2188 4482 2192
rect 4518 2188 4522 2192
rect 4558 2188 4562 2192
rect 326 2178 330 2182
rect 1774 2178 1778 2182
rect 2918 2178 2922 2182
rect 3134 2178 3138 2182
rect 6 2168 10 2172
rect 118 2168 122 2172
rect 790 2168 794 2172
rect 1158 2168 1162 2172
rect 1254 2168 1258 2172
rect 1438 2168 1442 2172
rect 2454 2168 2458 2172
rect 3118 2168 3122 2172
rect 3454 2168 3458 2172
rect 3518 2168 3522 2172
rect 3526 2168 3530 2172
rect 3702 2168 3706 2172
rect 3758 2168 3762 2172
rect 4038 2168 4042 2172
rect 4062 2168 4066 2172
rect 4134 2168 4138 2172
rect 4142 2168 4146 2172
rect 4254 2168 4258 2172
rect 4422 2168 4426 2172
rect 446 2158 450 2162
rect 574 2158 578 2162
rect 774 2158 778 2162
rect 830 2158 834 2162
rect 1110 2158 1114 2162
rect 1142 2158 1146 2162
rect 1206 2158 1210 2162
rect 1422 2158 1426 2162
rect 1462 2158 1466 2162
rect 2206 2158 2210 2162
rect 2222 2158 2226 2162
rect 2246 2158 2250 2162
rect 22 2148 26 2152
rect 46 2148 50 2152
rect 70 2148 74 2152
rect 94 2148 98 2152
rect 182 2147 186 2151
rect 238 2147 242 2151
rect 382 2148 386 2152
rect 430 2148 434 2152
rect 470 2148 474 2152
rect 542 2148 546 2152
rect 606 2147 610 2151
rect 678 2148 682 2152
rect 726 2147 730 2151
rect 798 2148 802 2152
rect 838 2148 842 2152
rect 870 2148 874 2152
rect 910 2148 914 2152
rect 998 2148 1002 2152
rect 1134 2148 1138 2152
rect 1182 2148 1186 2152
rect 1286 2148 1290 2152
rect 1334 2147 1338 2151
rect 1502 2148 1506 2152
rect 1670 2148 1674 2152
rect 1686 2148 1690 2152
rect 1702 2148 1706 2152
rect 1710 2148 1714 2152
rect 1726 2148 1730 2152
rect 1742 2148 1746 2152
rect 1750 2148 1754 2152
rect 1782 2148 1786 2152
rect 1830 2148 1834 2152
rect 1854 2147 1858 2151
rect 1950 2147 1954 2151
rect 2046 2147 2050 2151
rect 2126 2148 2130 2152
rect 2158 2147 2162 2151
rect 2222 2148 2226 2152
rect 2286 2158 2290 2162
rect 2318 2158 2322 2162
rect 2326 2158 2330 2162
rect 2366 2158 2370 2162
rect 2270 2148 2274 2152
rect 2302 2148 2306 2152
rect 2438 2158 2442 2162
rect 2662 2158 2666 2162
rect 2694 2158 2698 2162
rect 2742 2158 2746 2162
rect 2838 2158 2842 2162
rect 3006 2158 3010 2162
rect 3102 2158 3106 2162
rect 3198 2158 3202 2162
rect 3246 2158 3250 2162
rect 3270 2158 3274 2162
rect 3382 2158 3386 2162
rect 3510 2158 3514 2162
rect 3598 2158 3602 2162
rect 3718 2158 3722 2162
rect 3774 2158 3778 2162
rect 3790 2158 3794 2162
rect 3806 2158 3810 2162
rect 3950 2158 3954 2162
rect 4038 2158 4042 2162
rect 4046 2158 4050 2162
rect 4094 2158 4098 2162
rect 4126 2158 4130 2162
rect 4182 2158 4186 2162
rect 4230 2158 4234 2162
rect 2398 2148 2402 2152
rect 2430 2148 2434 2152
rect 2566 2148 2570 2152
rect 2598 2147 2602 2151
rect 2630 2148 2634 2152
rect 2654 2148 2658 2152
rect 2678 2148 2682 2152
rect 2758 2148 2762 2152
rect 2798 2148 2802 2152
rect 2846 2148 2850 2152
rect 318 2138 322 2142
rect 390 2138 394 2142
rect 422 2138 426 2142
rect 518 2138 522 2142
rect 534 2138 538 2142
rect 558 2138 562 2142
rect 590 2138 594 2142
rect 678 2138 682 2142
rect 830 2138 834 2142
rect 846 2138 850 2142
rect 990 2138 994 2142
rect 1038 2138 1042 2142
rect 1086 2138 1090 2142
rect 1094 2138 1098 2142
rect 1158 2138 1162 2142
rect 1206 2138 1210 2142
rect 1222 2138 1226 2142
rect 1230 2138 1234 2142
rect 1438 2138 1442 2142
rect 1462 2138 1466 2142
rect 1478 2138 1482 2142
rect 1590 2138 1594 2142
rect 1678 2138 1682 2142
rect 1694 2138 1698 2142
rect 1718 2138 1722 2142
rect 1734 2138 1738 2142
rect 1758 2138 1762 2142
rect 1774 2138 1778 2142
rect 1934 2138 1938 2142
rect 2030 2138 2034 2142
rect 2190 2138 2194 2142
rect 2206 2138 2210 2142
rect 2230 2138 2234 2142
rect 2278 2138 2282 2142
rect 2310 2138 2314 2142
rect 2350 2138 2354 2142
rect 2398 2138 2402 2142
rect 2454 2138 2458 2142
rect 2462 2138 2466 2142
rect 2510 2138 2514 2142
rect 2686 2138 2690 2142
rect 2718 2138 2722 2142
rect 2766 2138 2770 2142
rect 2782 2138 2786 2142
rect 2822 2138 2826 2142
rect 2870 2138 2874 2142
rect 3006 2148 3010 2152
rect 3030 2148 3034 2152
rect 3070 2148 3074 2152
rect 3078 2148 3082 2152
rect 3110 2148 3114 2152
rect 3150 2148 3154 2152
rect 3182 2148 3186 2152
rect 3230 2148 3234 2152
rect 3302 2148 3306 2152
rect 3318 2148 3322 2152
rect 3334 2148 3338 2152
rect 3350 2148 3354 2152
rect 3374 2148 3378 2152
rect 3422 2148 3426 2152
rect 3438 2148 3442 2152
rect 3462 2148 3466 2152
rect 3518 2148 3522 2152
rect 3646 2148 3650 2152
rect 3662 2148 3666 2152
rect 3670 2148 3674 2152
rect 3718 2148 3722 2152
rect 3734 2148 3738 2152
rect 3766 2148 3770 2152
rect 3790 2148 3794 2152
rect 3814 2148 3818 2152
rect 3830 2148 3834 2152
rect 3902 2148 3906 2152
rect 3918 2148 3922 2152
rect 3934 2148 3938 2152
rect 3982 2148 3986 2152
rect 4006 2148 4010 2152
rect 4030 2148 4034 2152
rect 4054 2148 4058 2152
rect 4086 2148 4090 2152
rect 4110 2148 4114 2152
rect 4134 2148 4138 2152
rect 4158 2148 4162 2152
rect 4198 2148 4202 2152
rect 4214 2148 4218 2152
rect 4286 2158 4290 2162
rect 4342 2158 4346 2162
rect 4462 2158 4466 2162
rect 4254 2148 4258 2152
rect 4286 2148 4290 2152
rect 4302 2148 4306 2152
rect 4326 2148 4330 2152
rect 4382 2148 4386 2152
rect 4430 2148 4434 2152
rect 4454 2148 4458 2152
rect 4478 2148 4482 2152
rect 4494 2148 4498 2152
rect 2966 2138 2970 2142
rect 2990 2138 2994 2142
rect 3022 2138 3026 2142
rect 3038 2138 3042 2142
rect 3062 2138 3066 2142
rect 3166 2138 3170 2142
rect 3222 2138 3226 2142
rect 3254 2138 3258 2142
rect 3270 2138 3274 2142
rect 3326 2138 3330 2142
rect 3358 2138 3362 2142
rect 3398 2138 3402 2142
rect 3414 2138 3418 2142
rect 3430 2138 3434 2142
rect 3494 2138 3498 2142
rect 3542 2138 3546 2142
rect 3558 2138 3562 2142
rect 3606 2138 3610 2142
rect 3678 2138 3682 2142
rect 3742 2138 3746 2142
rect 3782 2138 3786 2142
rect 3822 2138 3826 2142
rect 3846 2138 3850 2142
rect 3862 2138 3866 2142
rect 3902 2138 3906 2142
rect 3974 2138 3978 2142
rect 4118 2138 4122 2142
rect 4174 2138 4178 2142
rect 4198 2138 4202 2142
rect 4206 2138 4210 2142
rect 4262 2138 4266 2142
rect 4278 2138 4282 2142
rect 4310 2138 4314 2142
rect 4318 2138 4322 2142
rect 4390 2138 4394 2142
rect 4438 2138 4442 2142
rect 4486 2138 4490 2142
rect 4502 2138 4506 2142
rect 4566 2138 4570 2142
rect 102 2128 106 2132
rect 110 2128 114 2132
rect 182 2128 186 2132
rect 310 2128 314 2132
rect 694 2128 698 2132
rect 726 2128 730 2132
rect 918 2128 922 2132
rect 966 2128 970 2132
rect 998 2128 1002 2132
rect 1118 2128 1122 2132
rect 1134 2128 1138 2132
rect 1198 2128 1202 2132
rect 1334 2128 1338 2132
rect 1414 2128 1418 2132
rect 1454 2128 1458 2132
rect 1502 2128 1506 2132
rect 1806 2128 1810 2132
rect 1998 2128 2002 2132
rect 2326 2128 2330 2132
rect 2342 2128 2346 2132
rect 2734 2128 2738 2132
rect 2774 2128 2778 2132
rect 2806 2128 2810 2132
rect 2894 2128 2898 2132
rect 2910 2128 2914 2132
rect 2926 2128 2930 2132
rect 2934 2128 2938 2132
rect 2950 2128 2954 2132
rect 2958 2128 2962 2132
rect 2982 2128 2986 2132
rect 3126 2128 3130 2132
rect 3166 2128 3170 2132
rect 3206 2128 3210 2132
rect 3278 2128 3282 2132
rect 3318 2128 3322 2132
rect 3374 2128 3378 2132
rect 3502 2128 3506 2132
rect 3566 2128 3570 2132
rect 3574 2128 3578 2132
rect 3590 2128 3594 2132
rect 3622 2128 3626 2132
rect 3638 2128 3642 2132
rect 3646 2128 3650 2132
rect 3694 2128 3698 2132
rect 3702 2128 3706 2132
rect 3838 2128 3842 2132
rect 3878 2128 3882 2132
rect 3918 2128 3922 2132
rect 3990 2128 3994 2132
rect 4054 2128 4058 2132
rect 4174 2128 4178 2132
rect 4270 2128 4274 2132
rect 4350 2128 4354 2132
rect 4406 2128 4410 2132
rect 4414 2128 4418 2132
rect 4430 2128 4434 2132
rect 4518 2128 4522 2132
rect 4590 2128 4594 2132
rect 302 2118 306 2122
rect 446 2118 450 2122
rect 574 2118 578 2122
rect 686 2118 690 2122
rect 918 2118 922 2122
rect 982 2118 986 2122
rect 1110 2118 1114 2122
rect 1126 2118 1130 2122
rect 1398 2118 1402 2122
rect 1406 2118 1410 2122
rect 1422 2118 1426 2122
rect 1534 2118 1538 2122
rect 1654 2118 1658 2122
rect 1886 2118 1890 2122
rect 2094 2118 2098 2122
rect 2478 2118 2482 2122
rect 2534 2118 2538 2122
rect 2814 2118 2818 2122
rect 2862 2118 2866 2122
rect 3006 2118 3010 2122
rect 3094 2118 3098 2122
rect 3158 2118 3162 2122
rect 3214 2118 3218 2122
rect 3630 2118 3634 2122
rect 3710 2118 3714 2122
rect 3966 2118 3970 2122
rect 3998 2118 4002 2122
rect 4510 2118 4514 2122
rect 1002 2103 1006 2107
rect 1009 2103 1013 2107
rect 2026 2103 2030 2107
rect 2033 2103 2037 2107
rect 3050 2103 3054 2107
rect 3057 2103 3061 2107
rect 4082 2103 4086 2107
rect 4089 2103 4093 2107
rect 302 2088 306 2092
rect 774 2088 778 2092
rect 854 2088 858 2092
rect 1038 2088 1042 2092
rect 1398 2088 1402 2092
rect 1518 2088 1522 2092
rect 1622 2088 1626 2092
rect 1846 2088 1850 2092
rect 2446 2088 2450 2092
rect 2486 2088 2490 2092
rect 2582 2088 2586 2092
rect 2734 2088 2738 2092
rect 2782 2088 2786 2092
rect 2966 2088 2970 2092
rect 3038 2088 3042 2092
rect 3070 2088 3074 2092
rect 3118 2088 3122 2092
rect 3198 2088 3202 2092
rect 3246 2088 3250 2092
rect 3294 2088 3298 2092
rect 3310 2088 3314 2092
rect 3398 2088 3402 2092
rect 3502 2088 3506 2092
rect 3526 2088 3530 2092
rect 3550 2088 3554 2092
rect 3862 2088 3866 2092
rect 3878 2088 3882 2092
rect 4062 2088 4066 2092
rect 4254 2088 4258 2092
rect 4294 2088 4298 2092
rect 4334 2088 4338 2092
rect 4398 2088 4402 2092
rect 4414 2088 4418 2092
rect 4438 2088 4442 2092
rect 4470 2088 4474 2092
rect 4486 2088 4490 2092
rect 4518 2088 4522 2092
rect 4590 2088 4594 2092
rect 246 2078 250 2082
rect 262 2078 266 2082
rect 294 2078 298 2082
rect 782 2078 786 2082
rect 814 2078 818 2082
rect 974 2078 978 2082
rect 1006 2078 1010 2082
rect 1046 2078 1050 2082
rect 1078 2078 1082 2082
rect 1102 2078 1106 2082
rect 1158 2078 1162 2082
rect 1238 2078 1242 2082
rect 1278 2078 1282 2082
rect 1406 2078 1410 2082
rect 1510 2078 1514 2082
rect 1566 2078 1570 2082
rect 1598 2078 1602 2082
rect 1982 2078 1986 2082
rect 2126 2078 2130 2082
rect 2158 2078 2162 2082
rect 2246 2078 2250 2082
rect 2294 2078 2298 2082
rect 2366 2078 2370 2082
rect 2390 2078 2394 2082
rect 30 2068 34 2072
rect 134 2068 138 2072
rect 182 2068 186 2072
rect 230 2068 234 2072
rect 278 2068 282 2072
rect 310 2068 314 2072
rect 342 2068 346 2072
rect 358 2068 362 2072
rect 390 2068 394 2072
rect 414 2068 418 2072
rect 438 2068 442 2072
rect 542 2068 546 2072
rect 590 2068 594 2072
rect 662 2068 666 2072
rect 678 2068 682 2072
rect 694 2068 698 2072
rect 726 2068 730 2072
rect 830 2068 834 2072
rect 910 2068 914 2072
rect 982 2068 986 2072
rect 1030 2068 1034 2072
rect 1046 2068 1050 2072
rect 1126 2068 1130 2072
rect 22 2058 26 2062
rect 118 2059 122 2063
rect 214 2059 218 2063
rect 270 2058 274 2062
rect 286 2058 290 2062
rect 318 2058 322 2062
rect 326 2058 330 2062
rect 334 2058 338 2062
rect 366 2058 370 2062
rect 422 2058 426 2062
rect 470 2058 474 2062
rect 494 2058 498 2062
rect 518 2058 522 2062
rect 558 2059 562 2063
rect 654 2058 658 2062
rect 710 2059 714 2063
rect 814 2058 818 2062
rect 838 2058 842 2062
rect 886 2058 890 2062
rect 982 2058 986 2062
rect 1022 2058 1026 2062
rect 1070 2058 1074 2062
rect 1094 2058 1098 2062
rect 1198 2068 1202 2072
rect 1246 2068 1250 2072
rect 1262 2068 1266 2072
rect 1294 2068 1298 2072
rect 1326 2068 1330 2072
rect 1342 2068 1346 2072
rect 1358 2068 1362 2072
rect 1382 2068 1386 2072
rect 1454 2068 1458 2072
rect 1590 2068 1594 2072
rect 1630 2068 1634 2072
rect 1638 2068 1642 2072
rect 1646 2068 1650 2072
rect 1662 2068 1666 2072
rect 1678 2068 1682 2072
rect 1686 2068 1690 2072
rect 1694 2068 1698 2072
rect 1726 2068 1730 2072
rect 1750 2068 1754 2072
rect 1766 2068 1770 2072
rect 1934 2068 1938 2072
rect 2174 2068 2178 2072
rect 2222 2068 2226 2072
rect 2278 2068 2282 2072
rect 2302 2068 2306 2072
rect 2334 2068 2338 2072
rect 2590 2078 2594 2082
rect 2598 2078 2602 2082
rect 2694 2078 2698 2082
rect 2758 2078 2762 2082
rect 2790 2078 2794 2082
rect 2838 2078 2842 2082
rect 2878 2078 2882 2082
rect 2934 2078 2938 2082
rect 2974 2078 2978 2082
rect 3046 2078 3050 2082
rect 3078 2078 3082 2082
rect 3102 2078 3106 2082
rect 3134 2078 3138 2082
rect 3206 2078 3210 2082
rect 3214 2078 3218 2082
rect 3238 2078 3242 2082
rect 3278 2078 3282 2082
rect 3438 2078 3442 2082
rect 3486 2078 3490 2082
rect 3494 2078 3498 2082
rect 3534 2078 3538 2082
rect 3694 2078 3698 2082
rect 3718 2078 3722 2082
rect 3830 2078 3834 2082
rect 3870 2078 3874 2082
rect 3974 2078 3978 2082
rect 4070 2078 4074 2082
rect 4118 2078 4122 2082
rect 4166 2078 4170 2082
rect 4206 2078 4210 2082
rect 4222 2078 4226 2082
rect 2414 2068 2418 2072
rect 2462 2068 2466 2072
rect 2510 2068 2514 2072
rect 2518 2068 2522 2072
rect 2574 2068 2578 2072
rect 2606 2068 2610 2072
rect 2630 2068 2634 2072
rect 2678 2068 2682 2072
rect 2726 2068 2730 2072
rect 2750 2068 2754 2072
rect 2774 2068 2778 2072
rect 2798 2068 2802 2072
rect 2894 2068 2898 2072
rect 2990 2068 2994 2072
rect 3102 2068 3106 2072
rect 3150 2068 3154 2072
rect 3174 2068 3178 2072
rect 3190 2068 3194 2072
rect 3254 2068 3258 2072
rect 3302 2068 3306 2072
rect 3334 2068 3338 2072
rect 3390 2068 3394 2072
rect 3574 2068 3578 2072
rect 3606 2068 3610 2072
rect 3638 2068 3642 2072
rect 3654 2068 3658 2072
rect 3678 2068 3682 2072
rect 3694 2068 3698 2072
rect 3750 2068 3754 2072
rect 3766 2068 3770 2072
rect 3782 2068 3786 2072
rect 3814 2068 3818 2072
rect 1134 2058 1138 2062
rect 1174 2058 1178 2062
rect 1222 2058 1226 2062
rect 1238 2058 1242 2062
rect 1254 2058 1258 2062
rect 1302 2058 1306 2062
rect 1342 2058 1346 2062
rect 1366 2058 1370 2062
rect 1390 2058 1394 2062
rect 1438 2059 1442 2063
rect 1470 2058 1474 2062
rect 1550 2058 1554 2062
rect 1574 2058 1578 2062
rect 1670 2058 1674 2062
rect 1782 2059 1786 2063
rect 1886 2058 1890 2062
rect 1918 2059 1922 2063
rect 1982 2058 1986 2062
rect 2014 2059 2018 2063
rect 2094 2058 2098 2062
rect 2126 2059 2130 2063
rect 2222 2058 2226 2062
rect 2350 2058 2354 2062
rect 2406 2058 2410 2062
rect 2422 2058 2426 2062
rect 2446 2058 2450 2062
rect 2486 2058 2490 2062
rect 2502 2058 2506 2062
rect 2526 2058 2530 2062
rect 2654 2058 2658 2062
rect 2686 2058 2690 2062
rect 2710 2058 2714 2062
rect 2766 2058 2770 2062
rect 2814 2058 2818 2062
rect 2854 2058 2858 2062
rect 2878 2058 2882 2062
rect 2894 2058 2898 2062
rect 2918 2058 2922 2062
rect 2950 2058 2954 2062
rect 3022 2058 3026 2062
rect 3102 2058 3106 2062
rect 3182 2058 3186 2062
rect 3214 2058 3218 2062
rect 3230 2058 3234 2062
rect 3262 2058 3266 2062
rect 3326 2058 3330 2062
rect 3350 2058 3354 2062
rect 3374 2058 3378 2062
rect 3414 2058 3418 2062
rect 3454 2058 3458 2062
rect 3462 2058 3466 2062
rect 3510 2058 3514 2062
rect 3518 2058 3522 2062
rect 3558 2058 3562 2062
rect 3598 2058 3602 2062
rect 3630 2058 3634 2062
rect 3678 2058 3682 2062
rect 3694 2058 3698 2062
rect 3718 2058 3722 2062
rect 3758 2058 3762 2062
rect 3774 2058 3778 2062
rect 3790 2058 3794 2062
rect 3814 2058 3818 2062
rect 3846 2058 3850 2062
rect 3854 2058 3858 2062
rect 3894 2058 3898 2062
rect 3934 2068 3938 2072
rect 3958 2068 3962 2072
rect 3998 2068 4002 2072
rect 4014 2068 4018 2072
rect 4110 2068 4114 2072
rect 4126 2068 4130 2072
rect 4142 2068 4146 2072
rect 4166 2068 4170 2072
rect 4302 2078 4306 2082
rect 4342 2078 4346 2082
rect 4358 2078 4362 2082
rect 4366 2078 4370 2082
rect 4422 2078 4426 2082
rect 4430 2078 4434 2082
rect 4598 2078 4602 2082
rect 4270 2068 4274 2072
rect 4318 2068 4322 2072
rect 4446 2068 4450 2072
rect 4462 2068 4466 2072
rect 4478 2068 4482 2072
rect 4494 2068 4498 2072
rect 4542 2068 4546 2072
rect 4574 2068 4578 2072
rect 3926 2058 3930 2062
rect 3950 2058 3954 2062
rect 4022 2058 4026 2062
rect 4038 2058 4042 2062
rect 4046 2058 4050 2062
rect 4150 2058 4154 2062
rect 4190 2058 4194 2062
rect 4206 2058 4210 2062
rect 4262 2058 4266 2062
rect 4278 2058 4282 2062
rect 4382 2058 4386 2062
rect 4390 2058 4394 2062
rect 4406 2058 4410 2062
rect 4454 2058 4458 2062
rect 4510 2058 4514 2062
rect 4534 2058 4538 2062
rect 4566 2058 4570 2062
rect 4582 2058 4586 2062
rect 254 2048 258 2052
rect 382 2048 386 2052
rect 446 2048 450 2052
rect 678 2048 682 2052
rect 822 2048 826 2052
rect 878 2048 882 2052
rect 966 2048 970 2052
rect 1054 2048 1058 2052
rect 1150 2048 1154 2052
rect 1270 2048 1274 2052
rect 1318 2048 1322 2052
rect 1326 2048 1330 2052
rect 1366 2048 1370 2052
rect 1574 2048 1578 2052
rect 1662 2048 1666 2052
rect 1710 2048 1714 2052
rect 1734 2048 1738 2052
rect 1742 2048 1746 2052
rect 2158 2048 2162 2052
rect 2206 2048 2210 2052
rect 2318 2048 2322 2052
rect 2326 2048 2330 2052
rect 2462 2048 2466 2052
rect 2478 2048 2482 2052
rect 2486 2048 2490 2052
rect 2630 2048 2634 2052
rect 2646 2048 2650 2052
rect 2678 2048 2682 2052
rect 2710 2048 2714 2052
rect 2814 2048 2818 2052
rect 2854 2048 2858 2052
rect 2870 2048 2874 2052
rect 2942 2048 2946 2052
rect 3014 2048 3018 2052
rect 3286 2048 3290 2052
rect 3334 2048 3338 2052
rect 3374 2048 3378 2052
rect 3382 2048 3386 2052
rect 3398 2048 3402 2052
rect 3446 2048 3450 2052
rect 3542 2048 3546 2052
rect 3582 2048 3586 2052
rect 3614 2048 3618 2052
rect 3806 2048 3810 2052
rect 3878 2048 3882 2052
rect 3966 2048 3970 2052
rect 4030 2048 4034 2052
rect 4142 2048 4146 2052
rect 4198 2048 4202 2052
rect 4230 2048 4234 2052
rect 4294 2048 4298 2052
rect 4358 2048 4362 2052
rect 4518 2048 4522 2052
rect 4550 2048 4554 2052
rect 6 2038 10 2042
rect 150 2038 154 2042
rect 342 2038 346 2042
rect 462 2038 466 2042
rect 510 2038 514 2042
rect 526 2038 530 2042
rect 622 2038 626 2042
rect 758 2038 762 2042
rect 782 2038 786 2042
rect 806 2038 810 2042
rect 894 2038 898 2042
rect 1302 2038 1306 2042
rect 1830 2038 1834 2042
rect 2254 2038 2258 2042
rect 2438 2038 2442 2042
rect 2910 2038 2914 2042
rect 2934 2038 2938 2042
rect 3342 2038 3346 2042
rect 3846 2038 3850 2042
rect 4014 2038 4018 2042
rect 4182 2038 4186 2042
rect 886 2028 890 2032
rect 1718 2028 1722 2032
rect 2270 2028 2274 2032
rect 2806 2028 2810 2032
rect 470 2018 474 2022
rect 518 2018 522 2022
rect 638 2018 642 2022
rect 934 2018 938 2022
rect 1118 2018 1122 2022
rect 1134 2018 1138 2022
rect 1222 2018 1226 2022
rect 1286 2018 1290 2022
rect 1502 2018 1506 2022
rect 1854 2018 1858 2022
rect 1950 2018 1954 2022
rect 2054 2018 2058 2022
rect 2310 2018 2314 2022
rect 2702 2018 2706 2022
rect 3270 2018 3274 2022
rect 3622 2018 3626 2022
rect 3790 2018 3794 2022
rect 4078 2018 4082 2022
rect 4190 2018 4194 2022
rect 4398 2018 4402 2022
rect 4406 2018 4410 2022
rect 4566 2018 4570 2022
rect 498 2003 502 2007
rect 505 2003 509 2007
rect 1522 2003 1526 2007
rect 1529 2003 1533 2007
rect 2546 2003 2550 2007
rect 2553 2003 2557 2007
rect 3570 2003 3574 2007
rect 3577 2003 3581 2007
rect 150 1988 154 1992
rect 310 1988 314 1992
rect 414 1988 418 1992
rect 894 1988 898 1992
rect 1398 1988 1402 1992
rect 1430 1988 1434 1992
rect 1758 1988 1762 1992
rect 1822 1988 1826 1992
rect 2046 1988 2050 1992
rect 2350 1988 2354 1992
rect 2526 1988 2530 1992
rect 2798 1988 2802 1992
rect 2886 1988 2890 1992
rect 3006 1988 3010 1992
rect 3086 1988 3090 1992
rect 3182 1988 3186 1992
rect 3694 1988 3698 1992
rect 3782 1988 3786 1992
rect 3830 1988 3834 1992
rect 4094 1988 4098 1992
rect 4182 1988 4186 1992
rect 4254 1988 4258 1992
rect 4326 1988 4330 1992
rect 2630 1978 2634 1982
rect 2750 1978 2754 1982
rect 30 1968 34 1972
rect 54 1968 58 1972
rect 318 1968 322 1972
rect 398 1968 402 1972
rect 534 1968 538 1972
rect 630 1968 634 1972
rect 654 1968 658 1972
rect 686 1968 690 1972
rect 798 1968 802 1972
rect 998 1968 1002 1972
rect 1614 1968 1618 1972
rect 1998 1968 2002 1972
rect 2086 1968 2090 1972
rect 3534 1968 3538 1972
rect 3702 1968 3706 1972
rect 3966 1968 3970 1972
rect 4398 1968 4402 1972
rect 4494 1968 4498 1972
rect 22 1948 26 1952
rect 46 1948 50 1952
rect 118 1947 122 1951
rect 214 1947 218 1951
rect 254 1948 258 1952
rect 278 1958 282 1962
rect 334 1958 338 1962
rect 374 1958 378 1962
rect 382 1958 386 1962
rect 550 1958 554 1962
rect 582 1958 586 1962
rect 606 1958 610 1962
rect 614 1958 618 1962
rect 670 1958 674 1962
rect 702 1958 706 1962
rect 1174 1958 1178 1962
rect 1230 1958 1234 1962
rect 1510 1958 1514 1962
rect 302 1948 306 1952
rect 310 1948 314 1952
rect 398 1948 402 1952
rect 454 1948 458 1952
rect 478 1947 482 1951
rect 542 1948 546 1952
rect 566 1948 570 1952
rect 582 1948 586 1952
rect 630 1948 634 1952
rect 662 1948 666 1952
rect 678 1948 682 1952
rect 694 1948 698 1952
rect 734 1947 738 1951
rect 758 1948 762 1952
rect 830 1947 834 1951
rect 1062 1948 1066 1952
rect 1086 1948 1090 1952
rect 1110 1948 1114 1952
rect 1198 1948 1202 1952
rect 1214 1948 1218 1952
rect 1254 1948 1258 1952
rect 1334 1947 1338 1951
rect 1366 1948 1370 1952
rect 1462 1948 1466 1952
rect 1518 1948 1522 1952
rect 1550 1948 1554 1952
rect 1646 1958 1650 1962
rect 1678 1958 1682 1962
rect 1894 1958 1898 1962
rect 1982 1958 1986 1962
rect 2062 1958 2066 1962
rect 2070 1958 2074 1962
rect 2118 1958 2122 1962
rect 2286 1958 2290 1962
rect 2382 1958 2386 1962
rect 2446 1958 2450 1962
rect 2510 1958 2514 1962
rect 2542 1958 2546 1962
rect 2638 1958 2642 1962
rect 2678 1958 2682 1962
rect 2918 1958 2922 1962
rect 3054 1958 3058 1962
rect 3166 1958 3170 1962
rect 3222 1958 3226 1962
rect 3302 1958 3306 1962
rect 1638 1948 1642 1952
rect 1646 1948 1650 1952
rect 1694 1948 1698 1952
rect 1726 1948 1730 1952
rect 1742 1948 1746 1952
rect 1774 1948 1778 1952
rect 1814 1948 1818 1952
rect 1846 1948 1850 1952
rect 1854 1948 1858 1952
rect 1886 1948 1890 1952
rect 1934 1948 1938 1952
rect 1958 1948 1962 1952
rect 2046 1948 2050 1952
rect 2086 1948 2090 1952
rect 2158 1948 2162 1952
rect 2230 1948 2234 1952
rect 2286 1948 2290 1952
rect 2342 1948 2346 1952
rect 2374 1948 2378 1952
rect 2398 1948 2402 1952
rect 2470 1948 2474 1952
rect 2526 1948 2530 1952
rect 2678 1948 2682 1952
rect 2694 1948 2698 1952
rect 2742 1948 2746 1952
rect 2798 1948 2802 1952
rect 2838 1948 2842 1952
rect 2862 1948 2866 1952
rect 2982 1948 2986 1952
rect 3014 1948 3018 1952
rect 3078 1948 3082 1952
rect 3110 1948 3114 1952
rect 3198 1948 3202 1952
rect 3222 1948 3226 1952
rect 3238 1948 3242 1952
rect 3254 1948 3258 1952
rect 3454 1958 3458 1962
rect 3494 1958 3498 1962
rect 3518 1958 3522 1962
rect 3326 1948 3330 1952
rect 3374 1948 3378 1952
rect 3422 1948 3426 1952
rect 3590 1948 3594 1952
rect 3614 1958 3618 1962
rect 3718 1958 3722 1962
rect 3766 1958 3770 1962
rect 3822 1958 3826 1962
rect 3870 1958 3874 1962
rect 3902 1958 3906 1962
rect 3982 1958 3986 1962
rect 4014 1958 4018 1962
rect 4046 1958 4050 1962
rect 4166 1958 4170 1962
rect 4190 1958 4194 1962
rect 4294 1958 4298 1962
rect 3654 1948 3658 1952
rect 3662 1948 3666 1952
rect 3710 1948 3714 1952
rect 3742 1948 3746 1952
rect 3806 1948 3810 1952
rect 3822 1948 3826 1952
rect 3846 1948 3850 1952
rect 3854 1948 3858 1952
rect 3862 1948 3866 1952
rect 3878 1948 3882 1952
rect 3894 1948 3898 1952
rect 3918 1948 3922 1952
rect 3966 1948 3970 1952
rect 3998 1948 4002 1952
rect 4054 1948 4058 1952
rect 4118 1948 4122 1952
rect 4142 1948 4146 1952
rect 4198 1948 4202 1952
rect 4222 1948 4226 1952
rect 4238 1948 4242 1952
rect 4246 1948 4250 1952
rect 4326 1948 4330 1952
rect 4374 1948 4378 1952
rect 4398 1948 4402 1952
rect 4414 1948 4418 1952
rect 4566 1958 4570 1962
rect 4462 1948 4466 1952
rect 4494 1948 4498 1952
rect 4550 1948 4554 1952
rect 6 1938 10 1942
rect 134 1938 138 1942
rect 230 1938 234 1942
rect 246 1938 250 1942
rect 270 1938 274 1942
rect 294 1938 298 1942
rect 358 1938 362 1942
rect 406 1938 410 1942
rect 510 1938 514 1942
rect 558 1938 562 1942
rect 590 1938 594 1942
rect 638 1938 642 1942
rect 814 1938 818 1942
rect 902 1938 906 1942
rect 974 1938 978 1942
rect 1022 1938 1026 1942
rect 1078 1938 1082 1942
rect 1142 1938 1146 1942
rect 1158 1938 1162 1942
rect 1190 1938 1194 1942
rect 1222 1938 1226 1942
rect 1230 1938 1234 1942
rect 1246 1938 1250 1942
rect 1406 1938 1410 1942
rect 1470 1938 1474 1942
rect 1494 1938 1498 1942
rect 1510 1938 1514 1942
rect 1574 1938 1578 1942
rect 1614 1938 1618 1942
rect 1622 1940 1626 1944
rect 1670 1938 1674 1942
rect 1734 1938 1738 1942
rect 1782 1938 1786 1942
rect 1798 1938 1802 1942
rect 1822 1938 1826 1942
rect 1838 1938 1842 1942
rect 1862 1938 1866 1942
rect 1878 1938 1882 1942
rect 1910 1938 1914 1942
rect 1942 1938 1946 1942
rect 1998 1938 2002 1942
rect 2134 1938 2138 1942
rect 2214 1938 2218 1942
rect 2302 1938 2306 1942
rect 2318 1938 2322 1942
rect 2398 1938 2402 1942
rect 2422 1938 2426 1942
rect 2454 1938 2458 1942
rect 2494 1938 2498 1942
rect 2518 1938 2522 1942
rect 2614 1940 2618 1944
rect 2654 1938 2658 1942
rect 2670 1938 2674 1942
rect 2702 1938 2706 1942
rect 2710 1938 2714 1942
rect 2718 1940 2722 1944
rect 2766 1938 2770 1942
rect 2886 1938 2890 1942
rect 2902 1938 2906 1942
rect 2934 1938 2938 1942
rect 3038 1938 3042 1942
rect 3134 1938 3138 1942
rect 3150 1938 3154 1942
rect 3190 1938 3194 1942
rect 3246 1938 3250 1942
rect 3278 1938 3282 1942
rect 3286 1938 3290 1942
rect 3318 1938 3322 1942
rect 3334 1938 3338 1942
rect 3350 1938 3354 1942
rect 3430 1938 3434 1942
rect 3470 1938 3474 1942
rect 3502 1938 3506 1942
rect 3518 1938 3522 1942
rect 3542 1938 3546 1942
rect 3558 1938 3562 1942
rect 3582 1938 3586 1942
rect 3670 1938 3674 1942
rect 3750 1938 3754 1942
rect 3798 1938 3802 1942
rect 3838 1938 3842 1942
rect 3902 1938 3906 1942
rect 3934 1938 3938 1942
rect 3958 1938 3962 1942
rect 3990 1938 3994 1942
rect 4022 1938 4026 1942
rect 4062 1938 4066 1942
rect 4086 1938 4090 1942
rect 4150 1938 4154 1942
rect 4166 1938 4170 1942
rect 4254 1938 4258 1942
rect 4278 1938 4282 1942
rect 4366 1938 4370 1942
rect 4406 1938 4410 1942
rect 4486 1938 4490 1942
rect 4534 1938 4538 1942
rect 4542 1938 4546 1942
rect 4582 1938 4586 1942
rect 1046 1928 1050 1932
rect 1054 1928 1058 1932
rect 1070 1928 1074 1932
rect 1126 1928 1130 1932
rect 1142 1928 1146 1932
rect 1270 1928 1274 1932
rect 1278 1928 1282 1932
rect 1294 1928 1298 1932
rect 1486 1928 1490 1932
rect 1534 1928 1538 1932
rect 1582 1928 1586 1932
rect 1790 1928 1794 1932
rect 1862 1928 1866 1932
rect 2006 1928 2010 1932
rect 2110 1928 2114 1932
rect 2182 1928 2186 1932
rect 2278 1928 2282 1932
rect 2310 1928 2314 1932
rect 2430 1928 2434 1932
rect 2470 1928 2474 1932
rect 2566 1928 2570 1932
rect 2598 1928 2602 1932
rect 2662 1928 2666 1932
rect 2742 1928 2746 1932
rect 2846 1928 2850 1932
rect 2854 1928 2858 1932
rect 2878 1928 2882 1932
rect 2886 1928 2890 1932
rect 2942 1928 2946 1932
rect 2974 1928 2978 1932
rect 3030 1928 3034 1932
rect 3158 1928 3162 1932
rect 3174 1928 3178 1932
rect 3366 1928 3370 1932
rect 3406 1928 3410 1932
rect 3414 1928 3418 1932
rect 3638 1928 3642 1932
rect 3686 1928 3690 1932
rect 3726 1928 3730 1932
rect 3758 1928 3762 1932
rect 3774 1928 3778 1932
rect 3918 1928 3922 1932
rect 3950 1928 3954 1932
rect 4046 1928 4050 1932
rect 4078 1928 4082 1932
rect 4102 1928 4106 1932
rect 4126 1928 4130 1932
rect 4214 1928 4218 1932
rect 4294 1928 4298 1932
rect 4310 1928 4314 1932
rect 4350 1928 4354 1932
rect 4430 1928 4434 1932
rect 4478 1928 4482 1932
rect 4518 1928 4522 1932
rect 334 1918 338 1922
rect 374 1918 378 1922
rect 598 1918 602 1922
rect 662 1918 666 1922
rect 958 1918 962 1922
rect 1094 1918 1098 1922
rect 1150 1918 1154 1922
rect 1174 1918 1178 1922
rect 1286 1918 1290 1922
rect 1302 1918 1306 1922
rect 1478 1918 1482 1922
rect 1558 1918 1562 1922
rect 1894 1918 1898 1922
rect 1918 1918 1922 1922
rect 1974 1918 1978 1922
rect 2142 1918 2146 1922
rect 2462 1918 2466 1922
rect 2510 1918 2514 1922
rect 2638 1918 2642 1922
rect 3222 1918 3226 1922
rect 3358 1918 3362 1922
rect 3438 1918 3442 1922
rect 3454 1918 3458 1922
rect 3494 1918 3498 1922
rect 3518 1918 3522 1922
rect 3606 1918 3610 1922
rect 3646 1918 3650 1922
rect 3678 1918 3682 1922
rect 3734 1918 3738 1922
rect 3942 1918 3946 1922
rect 4158 1918 4162 1922
rect 4206 1918 4210 1922
rect 4438 1918 4442 1922
rect 4470 1918 4474 1922
rect 4558 1918 4562 1922
rect 4574 1918 4578 1922
rect 1002 1903 1006 1907
rect 1009 1903 1013 1907
rect 2026 1903 2030 1907
rect 2033 1903 2037 1907
rect 3050 1903 3054 1907
rect 3057 1903 3061 1907
rect 4082 1903 4086 1907
rect 4089 1903 4093 1907
rect 310 1888 314 1892
rect 534 1888 538 1892
rect 774 1888 778 1892
rect 902 1888 906 1892
rect 1110 1888 1114 1892
rect 1182 1888 1186 1892
rect 1534 1888 1538 1892
rect 1630 1888 1634 1892
rect 1694 1888 1698 1892
rect 1726 1888 1730 1892
rect 1934 1888 1938 1892
rect 1982 1888 1986 1892
rect 2198 1888 2202 1892
rect 2502 1888 2506 1892
rect 2542 1888 2546 1892
rect 2734 1888 2738 1892
rect 2862 1888 2866 1892
rect 2982 1888 2986 1892
rect 3030 1888 3034 1892
rect 3118 1888 3122 1892
rect 3830 1888 3834 1892
rect 3846 1888 3850 1892
rect 3918 1888 3922 1892
rect 3958 1888 3962 1892
rect 3982 1888 3986 1892
rect 4054 1888 4058 1892
rect 4142 1888 4146 1892
rect 4246 1888 4250 1892
rect 4310 1888 4314 1892
rect 4406 1888 4410 1892
rect 4438 1888 4442 1892
rect 4510 1888 4514 1892
rect 326 1878 330 1882
rect 342 1878 346 1882
rect 1118 1878 1122 1882
rect 6 1868 10 1872
rect 30 1868 34 1872
rect 134 1868 138 1872
rect 150 1868 154 1872
rect 214 1868 218 1872
rect 230 1868 234 1872
rect 350 1868 354 1872
rect 382 1868 386 1872
rect 446 1868 450 1872
rect 486 1868 490 1872
rect 550 1868 554 1872
rect 558 1868 562 1872
rect 614 1868 618 1872
rect 822 1868 826 1872
rect 918 1868 922 1872
rect 1030 1868 1034 1872
rect 1158 1878 1162 1882
rect 1206 1878 1210 1882
rect 1294 1878 1298 1882
rect 1326 1878 1330 1882
rect 1374 1878 1378 1882
rect 1382 1878 1386 1882
rect 1454 1878 1458 1882
rect 1190 1868 1194 1872
rect 1254 1868 1258 1872
rect 1262 1868 1266 1872
rect 1310 1868 1314 1872
rect 1382 1868 1386 1872
rect 1422 1868 1426 1872
rect 1550 1868 1554 1872
rect 1638 1868 1642 1872
rect 1686 1868 1690 1872
rect 1718 1868 1722 1872
rect 22 1858 26 1862
rect 118 1859 122 1863
rect 246 1859 250 1863
rect 358 1858 362 1862
rect 382 1858 386 1862
rect 438 1858 442 1862
rect 470 1858 474 1862
rect 534 1858 538 1862
rect 566 1858 570 1862
rect 598 1858 602 1862
rect 606 1858 610 1862
rect 638 1858 642 1862
rect 646 1858 650 1862
rect 678 1858 682 1862
rect 710 1859 714 1863
rect 742 1858 746 1862
rect 790 1858 794 1862
rect 806 1858 810 1862
rect 838 1859 842 1863
rect 870 1858 874 1862
rect 934 1859 938 1863
rect 958 1858 962 1862
rect 1046 1859 1050 1863
rect 1198 1858 1202 1862
rect 1246 1858 1250 1862
rect 1270 1858 1274 1862
rect 1342 1858 1346 1862
rect 1406 1858 1410 1862
rect 1462 1858 1466 1862
rect 1566 1859 1570 1863
rect 1638 1858 1642 1862
rect 1710 1858 1714 1862
rect 374 1848 378 1852
rect 478 1848 482 1852
rect 582 1848 586 1852
rect 782 1848 786 1852
rect 1230 1848 1234 1852
rect 1286 1848 1290 1852
rect 1334 1848 1338 1852
rect 1406 1848 1410 1852
rect 1422 1848 1426 1852
rect 1870 1878 1874 1882
rect 1886 1878 1890 1882
rect 1950 1878 1954 1882
rect 2054 1878 2058 1882
rect 2070 1878 2074 1882
rect 2102 1878 2106 1882
rect 2134 1878 2138 1882
rect 2334 1878 2338 1882
rect 2398 1878 2402 1882
rect 2406 1878 2410 1882
rect 2494 1878 2498 1882
rect 2566 1878 2570 1882
rect 2606 1878 2610 1882
rect 2622 1878 2626 1882
rect 2630 1878 2634 1882
rect 2662 1878 2666 1882
rect 2774 1878 2778 1882
rect 2902 1878 2906 1882
rect 2918 1878 2922 1882
rect 2934 1878 2938 1882
rect 2998 1878 3002 1882
rect 3046 1878 3050 1882
rect 3086 1878 3090 1882
rect 3238 1878 3242 1882
rect 3294 1878 3298 1882
rect 3318 1878 3322 1882
rect 3614 1878 3618 1882
rect 3718 1878 3722 1882
rect 1750 1868 1754 1872
rect 1766 1868 1770 1872
rect 1790 1868 1794 1872
rect 1806 1868 1810 1872
rect 1878 1868 1882 1872
rect 1918 1868 1922 1872
rect 1942 1868 1946 1872
rect 1974 1868 1978 1872
rect 2078 1868 2082 1872
rect 2142 1868 2146 1872
rect 2182 1868 2186 1872
rect 2206 1868 2210 1872
rect 2238 1868 2242 1872
rect 1742 1858 1746 1862
rect 1758 1858 1762 1862
rect 1774 1858 1778 1862
rect 1782 1858 1786 1862
rect 1798 1858 1802 1862
rect 1814 1858 1818 1862
rect 1854 1858 1858 1862
rect 1870 1858 1874 1862
rect 1990 1858 1994 1862
rect 2022 1858 2026 1862
rect 2078 1858 2082 1862
rect 2126 1858 2130 1862
rect 2230 1858 2234 1862
rect 2254 1858 2258 1862
rect 2374 1868 2378 1872
rect 2422 1868 2426 1872
rect 2510 1868 2514 1872
rect 2518 1868 2522 1872
rect 2742 1868 2746 1872
rect 2766 1868 2770 1872
rect 2798 1868 2802 1872
rect 2318 1858 2322 1862
rect 2350 1858 2354 1862
rect 2454 1858 2458 1862
rect 2478 1858 2482 1862
rect 2486 1858 2490 1862
rect 2606 1858 2610 1862
rect 2686 1858 2690 1862
rect 2710 1858 2714 1862
rect 2782 1858 2786 1862
rect 2830 1868 2834 1872
rect 2878 1868 2882 1872
rect 2886 1868 2890 1872
rect 2902 1868 2906 1872
rect 2934 1868 2938 1872
rect 2974 1868 2978 1872
rect 3014 1868 3018 1872
rect 3166 1868 3170 1872
rect 3198 1868 3202 1872
rect 3294 1868 3298 1872
rect 3358 1868 3362 1872
rect 3398 1868 3402 1872
rect 3422 1868 3426 1872
rect 3486 1868 3490 1872
rect 3550 1868 3554 1872
rect 3630 1868 3634 1872
rect 3710 1868 3714 1872
rect 3870 1878 3874 1882
rect 3926 1878 3930 1882
rect 4014 1878 4018 1882
rect 4078 1878 4082 1882
rect 4118 1878 4122 1882
rect 4150 1878 4154 1882
rect 4206 1878 4210 1882
rect 4278 1878 4282 1882
rect 4318 1878 4322 1882
rect 4446 1878 4450 1882
rect 3758 1868 3762 1872
rect 3814 1868 3818 1872
rect 3838 1868 3842 1872
rect 3862 1868 3866 1872
rect 3886 1868 3890 1872
rect 3934 1868 3938 1872
rect 3974 1868 3978 1872
rect 4014 1868 4018 1872
rect 4046 1868 4050 1872
rect 4134 1868 4138 1872
rect 4198 1868 4202 1872
rect 4230 1868 4234 1872
rect 4262 1868 4266 1872
rect 4270 1868 4274 1872
rect 4286 1868 4290 1872
rect 4358 1868 4362 1872
rect 4398 1868 4402 1872
rect 4414 1868 4418 1872
rect 4430 1868 4434 1872
rect 4446 1868 4450 1872
rect 4502 1878 4506 1882
rect 4518 1878 4522 1882
rect 4542 1878 4546 1882
rect 4582 1878 4586 1882
rect 4470 1868 4474 1872
rect 4486 1868 4490 1872
rect 4550 1868 4554 1872
rect 2822 1858 2826 1862
rect 2918 1858 2922 1862
rect 2958 1858 2962 1862
rect 3070 1858 3074 1862
rect 3102 1858 3106 1862
rect 3190 1858 3194 1862
rect 3230 1858 3234 1862
rect 3254 1858 3258 1862
rect 3270 1858 3274 1862
rect 3310 1858 3314 1862
rect 3342 1858 3346 1862
rect 3350 1858 3354 1862
rect 3374 1858 3378 1862
rect 3390 1858 3394 1862
rect 3414 1858 3418 1862
rect 3470 1858 3474 1862
rect 3534 1858 3538 1862
rect 3566 1858 3570 1862
rect 3574 1858 3578 1862
rect 3598 1858 3602 1862
rect 3638 1858 3642 1862
rect 3678 1858 3682 1862
rect 3734 1858 3738 1862
rect 3766 1858 3770 1862
rect 3806 1858 3810 1862
rect 3822 1858 3826 1862
rect 3942 1858 3946 1862
rect 3966 1858 3970 1862
rect 3998 1858 4002 1862
rect 4038 1858 4042 1862
rect 4102 1858 4106 1862
rect 4126 1858 4130 1862
rect 4174 1858 4178 1862
rect 4206 1858 4210 1862
rect 4222 1858 4226 1862
rect 4254 1858 4258 1862
rect 4294 1858 4298 1862
rect 4350 1858 4354 1862
rect 4374 1858 4378 1862
rect 4422 1858 4426 1862
rect 4478 1858 4482 1862
rect 4526 1858 4530 1862
rect 4542 1858 4546 1862
rect 4598 1858 4602 1862
rect 1838 1849 1842 1853
rect 1902 1848 1906 1852
rect 1926 1848 1930 1852
rect 2062 1848 2066 1852
rect 2166 1848 2170 1852
rect 2174 1848 2178 1852
rect 2190 1848 2194 1852
rect 2214 1848 2218 1852
rect 2230 1848 2234 1852
rect 2246 1848 2250 1852
rect 2278 1848 2282 1852
rect 2294 1848 2298 1852
rect 2438 1848 2442 1852
rect 2550 1848 2554 1852
rect 2590 1848 2594 1852
rect 2702 1848 2706 1852
rect 2750 1848 2754 1852
rect 2790 1848 2794 1852
rect 2822 1848 2826 1852
rect 2838 1848 2842 1852
rect 2854 1848 2858 1852
rect 2862 1848 2866 1852
rect 2966 1848 2970 1852
rect 3174 1848 3178 1852
rect 3206 1848 3210 1852
rect 3286 1848 3290 1852
rect 3334 1848 3338 1852
rect 3414 1848 3418 1852
rect 3454 1848 3458 1852
rect 3510 1848 3514 1852
rect 3654 1848 3658 1852
rect 3750 1848 3754 1852
rect 3782 1848 3786 1852
rect 3846 1848 3850 1852
rect 3886 1848 3890 1852
rect 3902 1848 3906 1852
rect 4022 1848 4026 1852
rect 4246 1848 4250 1852
rect 4310 1848 4314 1852
rect 4350 1848 4354 1852
rect 4366 1848 4370 1852
rect 4414 1848 4418 1852
rect 4558 1848 4562 1852
rect 4574 1848 4578 1852
rect 422 1838 426 1842
rect 438 1838 442 1842
rect 462 1838 466 1842
rect 622 1838 626 1842
rect 638 1838 642 1842
rect 798 1838 802 1842
rect 1350 1838 1354 1842
rect 1502 1838 1506 1842
rect 1734 1838 1738 1842
rect 2262 1838 2266 1842
rect 2294 1838 2298 1842
rect 2654 1838 2658 1842
rect 2678 1838 2682 1842
rect 2718 1838 2722 1842
rect 2950 1838 2954 1842
rect 3470 1838 3474 1842
rect 4110 1838 4114 1842
rect 4166 1838 4170 1842
rect 4382 1838 4386 1842
rect 4398 1838 4402 1842
rect 1214 1828 1218 1832
rect 318 1818 322 1822
rect 334 1818 338 1822
rect 390 1818 394 1822
rect 454 1818 458 1822
rect 998 1818 1002 1822
rect 1134 1818 1138 1822
rect 1270 1818 1274 1822
rect 1342 1818 1346 1822
rect 1366 1818 1370 1822
rect 1910 1818 1914 1822
rect 2254 1818 2258 1822
rect 2390 1818 2394 1822
rect 2414 1818 2418 1822
rect 2430 1818 2434 1822
rect 2470 1818 2474 1822
rect 2614 1818 2618 1822
rect 2686 1818 2690 1822
rect 2710 1818 2714 1822
rect 2814 1818 2818 1822
rect 2910 1818 2914 1822
rect 2942 1818 2946 1822
rect 3158 1818 3162 1822
rect 3190 1818 3194 1822
rect 3222 1818 3226 1822
rect 3302 1818 3306 1822
rect 3326 1818 3330 1822
rect 3430 1818 3434 1822
rect 3494 1818 3498 1822
rect 3534 1818 3538 1822
rect 3590 1818 3594 1822
rect 3622 1818 3626 1822
rect 3678 1818 3682 1822
rect 3734 1818 3738 1822
rect 3766 1818 3770 1822
rect 3806 1818 3810 1822
rect 3854 1818 3858 1822
rect 3878 1818 3882 1822
rect 4054 1818 4058 1822
rect 4174 1818 4178 1822
rect 4222 1818 4226 1822
rect 4454 1818 4458 1822
rect 4534 1818 4538 1822
rect 4590 1818 4594 1822
rect 498 1803 502 1807
rect 505 1803 509 1807
rect 1522 1803 1526 1807
rect 1529 1803 1533 1807
rect 2546 1803 2550 1807
rect 2553 1803 2557 1807
rect 3570 1803 3574 1807
rect 3577 1803 3581 1807
rect 30 1788 34 1792
rect 166 1788 170 1792
rect 206 1788 210 1792
rect 350 1788 354 1792
rect 782 1788 786 1792
rect 838 1788 842 1792
rect 958 1788 962 1792
rect 1182 1788 1186 1792
rect 1454 1788 1458 1792
rect 1566 1788 1570 1792
rect 1702 1788 1706 1792
rect 1942 1788 1946 1792
rect 1958 1788 1962 1792
rect 2094 1788 2098 1792
rect 2270 1788 2274 1792
rect 2526 1788 2530 1792
rect 2766 1788 2770 1792
rect 2806 1788 2810 1792
rect 2918 1788 2922 1792
rect 3134 1788 3138 1792
rect 3358 1788 3362 1792
rect 3550 1788 3554 1792
rect 3998 1788 4002 1792
rect 4030 1788 4034 1792
rect 4438 1788 4442 1792
rect 4558 1788 4562 1792
rect 590 1778 594 1782
rect 718 1778 722 1782
rect 6 1768 10 1772
rect 54 1768 58 1772
rect 374 1768 378 1772
rect 486 1768 490 1772
rect 598 1768 602 1772
rect 246 1758 250 1762
rect 310 1758 314 1762
rect 582 1758 586 1762
rect 718 1768 722 1772
rect 726 1768 730 1772
rect 758 1768 762 1772
rect 846 1768 850 1772
rect 1598 1768 1602 1772
rect 1638 1768 1642 1772
rect 1758 1768 1762 1772
rect 1894 1768 1898 1772
rect 1934 1768 1938 1772
rect 2142 1768 2146 1772
rect 2230 1768 2234 1772
rect 2662 1768 2666 1772
rect 3126 1768 3130 1772
rect 4390 1768 4394 1772
rect 4446 1768 4450 1772
rect 4454 1768 4458 1772
rect 862 1758 866 1762
rect 1030 1758 1034 1762
rect 1118 1758 1122 1762
rect 1166 1758 1170 1762
rect 1278 1758 1282 1762
rect 22 1748 26 1752
rect 46 1748 50 1752
rect 70 1748 74 1752
rect 102 1747 106 1751
rect 254 1748 258 1752
rect 302 1748 306 1752
rect 438 1747 442 1751
rect 550 1747 554 1751
rect 590 1748 594 1752
rect 638 1747 642 1751
rect 670 1748 674 1752
rect 718 1748 722 1752
rect 742 1748 746 1752
rect 798 1748 802 1752
rect 806 1748 810 1752
rect 854 1748 858 1752
rect 894 1747 898 1751
rect 918 1748 922 1752
rect 86 1738 90 1742
rect 222 1738 226 1742
rect 230 1738 234 1742
rect 246 1738 250 1742
rect 262 1738 266 1742
rect 286 1738 290 1742
rect 318 1738 322 1742
rect 366 1738 370 1742
rect 454 1738 458 1742
rect 534 1738 538 1742
rect 622 1738 626 1742
rect 830 1738 834 1742
rect 990 1748 994 1752
rect 1014 1748 1018 1752
rect 1094 1748 1098 1752
rect 1110 1748 1114 1752
rect 1182 1748 1186 1752
rect 1262 1748 1266 1752
rect 1358 1758 1362 1762
rect 1582 1758 1586 1762
rect 1614 1758 1618 1762
rect 1742 1758 1746 1762
rect 1926 1758 1930 1762
rect 1046 1738 1050 1742
rect 1086 1738 1090 1742
rect 1390 1747 1394 1751
rect 1422 1748 1426 1752
rect 1494 1748 1498 1752
rect 1606 1748 1610 1752
rect 1622 1748 1626 1752
rect 1654 1748 1658 1752
rect 1686 1748 1690 1752
rect 1718 1748 1722 1752
rect 1734 1748 1738 1752
rect 1750 1748 1754 1752
rect 1790 1748 1794 1752
rect 1798 1748 1802 1752
rect 1830 1748 1834 1752
rect 1894 1748 1898 1752
rect 1926 1748 1930 1752
rect 2174 1758 2178 1762
rect 2198 1758 2202 1762
rect 2382 1758 2386 1762
rect 2390 1758 2394 1762
rect 2438 1758 2442 1762
rect 2446 1758 2450 1762
rect 2534 1758 2538 1762
rect 2846 1758 2850 1762
rect 2862 1758 2866 1762
rect 2942 1758 2946 1762
rect 3142 1758 3146 1762
rect 3166 1758 3170 1762
rect 2078 1748 2082 1752
rect 2134 1748 2138 1752
rect 2214 1748 2218 1752
rect 2238 1748 2242 1752
rect 2278 1748 2282 1752
rect 2318 1748 2322 1752
rect 2342 1748 2346 1752
rect 2422 1748 2426 1752
rect 2486 1748 2490 1752
rect 2582 1748 2586 1752
rect 2614 1748 2618 1752
rect 2646 1748 2650 1752
rect 2654 1748 2658 1752
rect 2686 1748 2690 1752
rect 2694 1748 2698 1752
rect 2726 1748 2730 1752
rect 2774 1748 2778 1752
rect 2814 1748 2818 1752
rect 2822 1748 2826 1752
rect 2854 1748 2858 1752
rect 2990 1748 2994 1752
rect 3006 1748 3010 1752
rect 3046 1748 3050 1752
rect 3094 1748 3098 1752
rect 3134 1748 3138 1752
rect 3230 1758 3234 1762
rect 3262 1758 3266 1762
rect 3294 1758 3298 1762
rect 3302 1758 3306 1762
rect 3318 1758 3322 1762
rect 3326 1758 3330 1762
rect 3390 1758 3394 1762
rect 3190 1748 3194 1752
rect 3206 1748 3210 1752
rect 3246 1748 3250 1752
rect 3262 1748 3266 1752
rect 3278 1748 3282 1752
rect 3302 1748 3306 1752
rect 3342 1748 3346 1752
rect 3406 1748 3410 1752
rect 3446 1758 3450 1762
rect 3470 1758 3474 1762
rect 3526 1758 3530 1762
rect 3622 1758 3626 1762
rect 3750 1758 3754 1762
rect 3782 1758 3786 1762
rect 3814 1758 3818 1762
rect 3862 1758 3866 1762
rect 3910 1758 3914 1762
rect 3918 1758 3922 1762
rect 4094 1758 4098 1762
rect 4334 1758 4338 1762
rect 3510 1748 3514 1752
rect 3566 1748 3570 1752
rect 3606 1748 3610 1752
rect 3630 1748 3634 1752
rect 3646 1748 3650 1752
rect 3678 1748 3682 1752
rect 3702 1748 3706 1752
rect 3798 1748 3802 1752
rect 3838 1748 3842 1752
rect 3862 1748 3866 1752
rect 3934 1748 3938 1752
rect 3974 1748 3978 1752
rect 3982 1748 3986 1752
rect 4014 1748 4018 1752
rect 4110 1748 4114 1752
rect 4142 1748 4146 1752
rect 4166 1748 4170 1752
rect 4206 1748 4210 1752
rect 4246 1748 4250 1752
rect 4262 1748 4266 1752
rect 4278 1748 4282 1752
rect 4310 1748 4314 1752
rect 4350 1748 4354 1752
rect 4366 1748 4370 1752
rect 4390 1748 4394 1752
rect 4414 1758 4418 1762
rect 4502 1758 4506 1762
rect 4454 1748 4458 1752
rect 4486 1748 4490 1752
rect 4542 1748 4546 1752
rect 4590 1748 4594 1752
rect 1142 1738 1146 1742
rect 1190 1738 1194 1742
rect 1198 1738 1202 1742
rect 1246 1738 1250 1742
rect 1254 1738 1258 1742
rect 1302 1738 1306 1742
rect 1326 1738 1330 1742
rect 1502 1738 1506 1742
rect 1662 1738 1666 1742
rect 1686 1738 1690 1742
rect 1822 1738 1826 1742
rect 1894 1738 1898 1742
rect 1974 1738 1978 1742
rect 2070 1738 2074 1742
rect 2118 1738 2122 1742
rect 2158 1738 2162 1742
rect 2174 1738 2178 1742
rect 2182 1738 2186 1742
rect 2190 1738 2194 1742
rect 2198 1738 2202 1742
rect 2310 1738 2314 1742
rect 2366 1738 2370 1742
rect 2406 1738 2410 1742
rect 2414 1738 2418 1742
rect 2462 1738 2466 1742
rect 2494 1738 2498 1742
rect 2590 1738 2594 1742
rect 2606 1738 2610 1742
rect 2630 1738 2634 1742
rect 2638 1738 2642 1742
rect 2662 1738 2666 1742
rect 2678 1738 2682 1742
rect 2702 1738 2706 1742
rect 2734 1738 2738 1742
rect 2790 1738 2794 1742
rect 2822 1738 2826 1742
rect 2926 1738 2930 1742
rect 2942 1738 2946 1742
rect 2958 1740 2962 1744
rect 2982 1738 2986 1742
rect 3014 1738 3018 1742
rect 3150 1738 3154 1742
rect 3182 1738 3186 1742
rect 3198 1738 3202 1742
rect 3206 1738 3210 1742
rect 3238 1738 3242 1742
rect 3270 1738 3274 1742
rect 3318 1738 3322 1742
rect 3334 1738 3338 1742
rect 3366 1738 3370 1742
rect 3414 1738 3418 1742
rect 3470 1738 3474 1742
rect 3486 1738 3490 1742
rect 3518 1738 3522 1742
rect 3542 1738 3546 1742
rect 3574 1738 3578 1742
rect 3598 1738 3602 1742
rect 3630 1738 3634 1742
rect 3686 1738 3690 1742
rect 3694 1738 3698 1742
rect 3726 1738 3730 1742
rect 3742 1738 3746 1742
rect 3758 1740 3762 1744
rect 3806 1738 3810 1742
rect 3830 1738 3834 1742
rect 3862 1738 3866 1742
rect 3878 1738 3882 1742
rect 3886 1738 3890 1742
rect 3926 1738 3930 1742
rect 3942 1738 3946 1742
rect 3966 1738 3970 1742
rect 4046 1738 4050 1742
rect 4054 1740 4058 1744
rect 4118 1738 4122 1742
rect 4166 1738 4170 1742
rect 4182 1738 4186 1742
rect 4198 1738 4202 1742
rect 4222 1738 4226 1742
rect 4238 1738 4242 1742
rect 4254 1738 4258 1742
rect 4286 1738 4290 1742
rect 4318 1738 4322 1742
rect 4342 1738 4346 1742
rect 4374 1738 4378 1742
rect 4430 1738 4434 1742
rect 4494 1738 4498 1742
rect 4518 1738 4522 1742
rect 4534 1738 4538 1742
rect 4566 1738 4570 1742
rect 278 1728 282 1732
rect 966 1728 970 1732
rect 1022 1728 1026 1732
rect 1054 1728 1058 1732
rect 1078 1728 1082 1732
rect 1110 1728 1114 1732
rect 1158 1728 1162 1732
rect 1334 1728 1338 1732
rect 1582 1728 1586 1732
rect 1726 1728 1730 1732
rect 1774 1728 1778 1732
rect 1790 1728 1794 1732
rect 1854 1728 1858 1732
rect 1886 1728 1890 1732
rect 1950 1728 1954 1732
rect 2006 1728 2010 1732
rect 2030 1728 2034 1732
rect 2078 1728 2082 1732
rect 2126 1728 2130 1732
rect 2150 1728 2154 1732
rect 2238 1728 2242 1732
rect 2254 1728 2258 1732
rect 2262 1728 2266 1732
rect 2302 1728 2306 1732
rect 2334 1728 2338 1732
rect 2358 1728 2362 1732
rect 2502 1728 2506 1732
rect 2510 1728 2514 1732
rect 2574 1728 2578 1732
rect 2598 1728 2602 1732
rect 2622 1728 2626 1732
rect 2718 1728 2722 1732
rect 2750 1728 2754 1732
rect 2758 1728 2762 1732
rect 2798 1728 2802 1732
rect 2870 1728 2874 1732
rect 2878 1728 2882 1732
rect 2902 1728 2906 1732
rect 2910 1728 2914 1732
rect 3022 1728 3026 1732
rect 3070 1728 3074 1732
rect 3110 1728 3114 1732
rect 3374 1728 3378 1732
rect 3534 1728 3538 1732
rect 3646 1728 3650 1732
rect 3854 1728 3858 1732
rect 3950 1728 3954 1732
rect 4278 1728 4282 1732
rect 4294 1728 4298 1732
rect 4574 1728 4578 1732
rect 238 1718 242 1722
rect 974 1718 978 1722
rect 1222 1718 1226 1722
rect 1286 1718 1290 1722
rect 1310 1718 1314 1722
rect 1350 1718 1354 1722
rect 1606 1718 1610 1722
rect 1670 1718 1674 1722
rect 1758 1718 1762 1722
rect 1782 1718 1786 1722
rect 1846 1718 1850 1722
rect 1862 1718 1866 1722
rect 1990 1718 1994 1722
rect 2286 1718 2290 1722
rect 2326 1718 2330 1722
rect 2350 1718 2354 1722
rect 2382 1718 2386 1722
rect 2390 1718 2394 1722
rect 2438 1718 2442 1722
rect 2454 1718 2458 1722
rect 2470 1718 2474 1722
rect 2742 1718 2746 1722
rect 2782 1718 2786 1722
rect 2846 1718 2850 1722
rect 2942 1718 2946 1722
rect 2974 1718 2978 1722
rect 3006 1718 3010 1722
rect 3030 1718 3034 1722
rect 3230 1718 3234 1722
rect 3382 1718 3386 1722
rect 3398 1718 3402 1722
rect 3438 1718 3442 1722
rect 3494 1718 3498 1722
rect 3678 1718 3682 1722
rect 3718 1718 3722 1722
rect 3774 1718 3778 1722
rect 3782 1718 3786 1722
rect 3822 1718 3826 1722
rect 3910 1718 3914 1722
rect 3958 1718 3962 1722
rect 4070 1718 4074 1722
rect 4086 1718 4090 1722
rect 4190 1718 4194 1722
rect 4230 1718 4234 1722
rect 4302 1718 4306 1722
rect 4326 1718 4330 1722
rect 4366 1718 4370 1722
rect 1002 1703 1006 1707
rect 1009 1703 1013 1707
rect 2026 1703 2030 1707
rect 2033 1703 2037 1707
rect 3050 1703 3054 1707
rect 3057 1703 3061 1707
rect 4082 1703 4086 1707
rect 4089 1703 4093 1707
rect 54 1688 58 1692
rect 278 1688 282 1692
rect 366 1688 370 1692
rect 438 1688 442 1692
rect 670 1688 674 1692
rect 910 1688 914 1692
rect 1022 1688 1026 1692
rect 1134 1688 1138 1692
rect 1158 1688 1162 1692
rect 1198 1688 1202 1692
rect 1278 1688 1282 1692
rect 1886 1688 1890 1692
rect 2038 1688 2042 1692
rect 2174 1688 2178 1692
rect 2342 1688 2346 1692
rect 2830 1688 2834 1692
rect 2854 1688 2858 1692
rect 2870 1688 2874 1692
rect 2966 1688 2970 1692
rect 3006 1688 3010 1692
rect 3326 1688 3330 1692
rect 3614 1688 3618 1692
rect 4590 1688 4594 1692
rect 214 1678 218 1682
rect 222 1678 226 1682
rect 270 1678 274 1682
rect 302 1678 306 1682
rect 382 1678 386 1682
rect 766 1678 770 1682
rect 1166 1678 1170 1682
rect 1174 1678 1178 1682
rect 1222 1678 1226 1682
rect 1238 1678 1242 1682
rect 1270 1678 1274 1682
rect 1302 1678 1306 1682
rect 1318 1678 1322 1682
rect 1446 1678 1450 1682
rect 1798 1678 1802 1682
rect 1974 1678 1978 1682
rect 2118 1678 2122 1682
rect 2150 1678 2154 1682
rect 2166 1678 2170 1682
rect 2430 1678 2434 1682
rect 2446 1678 2450 1682
rect 2494 1678 2498 1682
rect 2502 1678 2506 1682
rect 2614 1678 2618 1682
rect 2622 1678 2626 1682
rect 2678 1678 2682 1682
rect 2766 1678 2770 1682
rect 2798 1678 2802 1682
rect 2926 1678 2930 1682
rect 2934 1678 2938 1682
rect 2974 1678 2978 1682
rect 3070 1678 3074 1682
rect 3142 1678 3146 1682
rect 3254 1678 3258 1682
rect 3270 1678 3274 1682
rect 3398 1678 3402 1682
rect 3462 1678 3466 1682
rect 3478 1678 3482 1682
rect 3710 1678 3714 1682
rect 3766 1678 3770 1682
rect 3854 1678 3858 1682
rect 3926 1678 3930 1682
rect 4198 1678 4202 1682
rect 4246 1678 4250 1682
rect 4254 1678 4258 1682
rect 4318 1678 4322 1682
rect 4358 1678 4362 1682
rect 4414 1678 4418 1682
rect 4430 1678 4434 1682
rect 30 1668 34 1672
rect 150 1668 154 1672
rect 198 1668 202 1672
rect 286 1668 290 1672
rect 342 1668 346 1672
rect 406 1668 410 1672
rect 534 1668 538 1672
rect 622 1668 626 1672
rect 966 1668 970 1672
rect 1054 1668 1058 1672
rect 1150 1668 1154 1672
rect 1206 1668 1210 1672
rect 1262 1668 1266 1672
rect 1342 1668 1346 1672
rect 1350 1668 1354 1672
rect 1366 1668 1370 1672
rect 1414 1668 1418 1672
rect 1534 1668 1538 1672
rect 1550 1668 1554 1672
rect 1598 1668 1602 1672
rect 1638 1668 1642 1672
rect 1694 1668 1698 1672
rect 1702 1668 1706 1672
rect 1718 1668 1722 1672
rect 1758 1668 1762 1672
rect 1814 1668 1818 1672
rect 1846 1668 1850 1672
rect 1854 1668 1858 1672
rect 1902 1668 1906 1672
rect 1926 1668 1930 1672
rect 1982 1668 1986 1672
rect 2006 1668 2010 1672
rect 2054 1668 2058 1672
rect 2182 1668 2186 1672
rect 22 1658 26 1662
rect 46 1658 50 1662
rect 86 1658 90 1662
rect 118 1659 122 1663
rect 190 1658 194 1662
rect 246 1658 250 1662
rect 286 1658 290 1662
rect 326 1658 330 1662
rect 350 1658 354 1662
rect 478 1658 482 1662
rect 502 1659 506 1663
rect 542 1658 546 1662
rect 566 1658 570 1662
rect 606 1659 610 1663
rect 686 1658 690 1662
rect 718 1658 722 1662
rect 766 1659 770 1663
rect 854 1658 858 1662
rect 862 1658 866 1662
rect 886 1658 890 1662
rect 926 1658 930 1662
rect 958 1659 962 1663
rect 1070 1659 1074 1663
rect 1142 1658 1146 1662
rect 1214 1658 1218 1662
rect 1254 1658 1258 1662
rect 1270 1658 1274 1662
rect 1286 1658 1290 1662
rect 1446 1659 1450 1663
rect 1550 1658 1554 1662
rect 1582 1658 1586 1662
rect 1614 1658 1618 1662
rect 1686 1658 1690 1662
rect 1726 1658 1730 1662
rect 1742 1658 1746 1662
rect 1750 1658 1754 1662
rect 1782 1658 1786 1662
rect 1950 1658 1954 1662
rect 2094 1658 2098 1662
rect 2102 1658 2106 1662
rect 2126 1658 2130 1662
rect 2142 1658 2146 1662
rect 2222 1666 2226 1670
rect 2246 1668 2250 1672
rect 2262 1668 2266 1672
rect 2350 1668 2354 1672
rect 2374 1668 2378 1672
rect 2510 1668 2514 1672
rect 2534 1668 2538 1672
rect 2638 1668 2642 1672
rect 2718 1668 2722 1672
rect 2742 1668 2746 1672
rect 2790 1668 2794 1672
rect 2806 1668 2810 1672
rect 2894 1668 2898 1672
rect 2918 1668 2922 1672
rect 2950 1668 2954 1672
rect 2990 1668 2994 1672
rect 3006 1668 3010 1672
rect 3086 1668 3090 1672
rect 3118 1668 3122 1672
rect 3166 1668 3170 1672
rect 3190 1668 3194 1672
rect 3342 1668 3346 1672
rect 3406 1668 3410 1672
rect 3438 1668 3442 1672
rect 3454 1668 3458 1672
rect 3646 1668 3650 1672
rect 3670 1668 3674 1672
rect 3814 1668 3818 1672
rect 3846 1668 3850 1672
rect 3870 1668 3874 1672
rect 3902 1668 3906 1672
rect 3958 1668 3962 1672
rect 3966 1668 3970 1672
rect 4022 1668 4026 1672
rect 4046 1668 4050 1672
rect 4054 1668 4058 1672
rect 4102 1668 4106 1672
rect 4134 1668 4138 1672
rect 4142 1668 4146 1672
rect 4206 1668 4210 1672
rect 4246 1668 4250 1672
rect 4262 1668 4266 1672
rect 4318 1668 4322 1672
rect 4366 1668 4370 1672
rect 4574 1678 4578 1682
rect 4598 1678 4602 1682
rect 4454 1668 4458 1672
rect 4502 1668 4506 1672
rect 2278 1658 2282 1662
rect 2302 1658 2306 1662
rect 2310 1658 2314 1662
rect 2398 1658 2402 1662
rect 2430 1658 2434 1662
rect 2478 1658 2482 1662
rect 2590 1658 2594 1662
rect 2622 1658 2626 1662
rect 2654 1658 2658 1662
rect 2694 1658 2698 1662
rect 2750 1658 2754 1662
rect 2814 1658 2818 1662
rect 2838 1658 2842 1662
rect 2886 1658 2890 1662
rect 2982 1658 2986 1662
rect 3014 1658 3018 1662
rect 3022 1658 3026 1662
rect 3046 1658 3050 1662
rect 3094 1658 3098 1662
rect 3110 1658 3114 1662
rect 3158 1658 3162 1662
rect 3198 1658 3202 1662
rect 3230 1658 3234 1662
rect 3270 1658 3274 1662
rect 3310 1658 3314 1662
rect 3318 1658 3322 1662
rect 3342 1658 3346 1662
rect 3358 1658 3362 1662
rect 3390 1658 3394 1662
rect 3430 1658 3434 1662
rect 3446 1658 3450 1662
rect 3494 1658 3498 1662
rect 3518 1658 3522 1662
rect 3526 1658 3530 1662
rect 3534 1658 3538 1662
rect 3542 1658 3546 1662
rect 3574 1658 3578 1662
rect 3590 1658 3594 1662
rect 3646 1658 3650 1662
rect 3670 1658 3674 1662
rect 3686 1658 3690 1662
rect 3742 1658 3746 1662
rect 3774 1658 3778 1662
rect 3782 1658 3786 1662
rect 3806 1658 3810 1662
rect 3838 1658 3842 1662
rect 3878 1658 3882 1662
rect 3894 1658 3898 1662
rect 3902 1658 3906 1662
rect 3950 1658 3954 1662
rect 3974 1658 3978 1662
rect 4014 1658 4018 1662
rect 4062 1658 4066 1662
rect 4126 1658 4130 1662
rect 4174 1658 4178 1662
rect 4302 1658 4306 1662
rect 4374 1658 4378 1662
rect 4382 1658 4386 1662
rect 4414 1658 4418 1662
rect 4462 1658 4466 1662
rect 4486 1658 4490 1662
rect 4526 1658 4530 1662
rect 4534 1658 4538 1662
rect 4558 1658 4562 1662
rect 4582 1658 4586 1662
rect 166 1648 170 1652
rect 310 1648 314 1652
rect 366 1648 370 1652
rect 390 1648 394 1652
rect 430 1648 434 1652
rect 574 1648 578 1652
rect 6 1638 10 1642
rect 174 1638 178 1642
rect 238 1638 242 1642
rect 326 1638 330 1642
rect 454 1638 458 1642
rect 558 1638 562 1642
rect 718 1648 722 1652
rect 894 1648 898 1652
rect 1326 1648 1330 1652
rect 1518 1648 1522 1652
rect 1734 1648 1738 1652
rect 1790 1648 1794 1652
rect 1830 1648 1834 1652
rect 1878 1648 1882 1652
rect 1886 1648 1890 1652
rect 1910 1648 1914 1652
rect 1998 1648 2002 1652
rect 2070 1648 2074 1652
rect 2078 1648 2082 1652
rect 2094 1648 2098 1652
rect 2206 1648 2210 1652
rect 2246 1648 2250 1652
rect 2358 1648 2362 1652
rect 2454 1648 2458 1652
rect 2534 1648 2538 1652
rect 2550 1648 2554 1652
rect 2670 1648 2674 1652
rect 2702 1648 2706 1652
rect 2718 1648 2722 1652
rect 2870 1648 2874 1652
rect 3094 1648 3098 1652
rect 3134 1648 3138 1652
rect 3182 1648 3186 1652
rect 3214 1648 3218 1652
rect 3326 1648 3330 1652
rect 3430 1648 3434 1652
rect 3630 1648 3634 1652
rect 3654 1648 3658 1652
rect 3678 1648 3682 1652
rect 3726 1648 3730 1652
rect 3822 1648 3826 1652
rect 3838 1648 3842 1652
rect 3894 1648 3898 1652
rect 3926 1648 3930 1652
rect 3934 1648 3938 1652
rect 3950 1648 3954 1652
rect 3990 1648 3994 1652
rect 4078 1648 4082 1652
rect 4158 1648 4162 1652
rect 4406 1648 4410 1652
rect 4526 1648 4530 1652
rect 694 1638 698 1642
rect 726 1638 730 1642
rect 846 1638 850 1642
rect 878 1638 882 1642
rect 1622 1638 1626 1642
rect 1654 1638 1658 1642
rect 1766 1638 1770 1642
rect 1774 1638 1778 1642
rect 1782 1638 1786 1642
rect 1982 1638 1986 1642
rect 2262 1638 2266 1642
rect 2422 1638 2426 1642
rect 2694 1638 2698 1642
rect 2718 1638 2722 1642
rect 3110 1638 3114 1642
rect 3238 1638 3242 1642
rect 3694 1638 3698 1642
rect 3854 1638 3858 1642
rect 4182 1638 4186 1642
rect 4302 1638 4306 1642
rect 4534 1638 4538 1642
rect 686 1628 690 1632
rect 1390 1628 1394 1632
rect 214 1618 218 1622
rect 246 1618 250 1622
rect 374 1618 378 1622
rect 398 1618 402 1622
rect 422 1618 426 1622
rect 718 1618 722 1622
rect 830 1618 834 1622
rect 838 1618 842 1622
rect 870 1618 874 1622
rect 910 1618 914 1622
rect 1294 1618 1298 1622
rect 1310 1618 1314 1622
rect 1334 1618 1338 1622
rect 1358 1618 1362 1622
rect 1614 1618 1618 1622
rect 1702 1618 1706 1622
rect 1862 1618 1866 1622
rect 1950 1618 1954 1622
rect 2126 1618 2130 1622
rect 2150 1618 2154 1622
rect 2198 1618 2202 1622
rect 2238 1618 2242 1622
rect 2286 1618 2290 1622
rect 2326 1618 2330 1622
rect 2398 1618 2402 1622
rect 2462 1618 2466 1622
rect 2582 1618 2586 1622
rect 2638 1618 2642 1622
rect 2654 1618 2658 1622
rect 2734 1618 2738 1622
rect 2750 1618 2754 1622
rect 2774 1618 2778 1622
rect 2854 1618 2858 1622
rect 2902 1618 2906 1622
rect 3022 1618 3026 1622
rect 3150 1618 3154 1622
rect 3174 1618 3178 1622
rect 3302 1618 3306 1622
rect 3366 1618 3370 1622
rect 3502 1618 3506 1622
rect 3550 1618 3554 1622
rect 3686 1618 3690 1622
rect 3718 1618 3722 1622
rect 3742 1618 3746 1622
rect 4014 1618 4018 1622
rect 4038 1618 4042 1622
rect 4126 1618 4130 1622
rect 4174 1618 4178 1622
rect 4238 1618 4242 1622
rect 4294 1618 4298 1622
rect 4486 1618 4490 1622
rect 498 1603 502 1607
rect 505 1603 509 1607
rect 1522 1603 1526 1607
rect 1529 1603 1533 1607
rect 2546 1603 2550 1607
rect 2553 1603 2557 1607
rect 3570 1603 3574 1607
rect 3577 1603 3581 1607
rect 254 1588 258 1592
rect 558 1588 562 1592
rect 726 1588 730 1592
rect 750 1588 754 1592
rect 982 1588 986 1592
rect 1694 1588 1698 1592
rect 1798 1588 1802 1592
rect 1886 1588 1890 1592
rect 2814 1588 2818 1592
rect 2838 1588 2842 1592
rect 3022 1588 3026 1592
rect 3046 1588 3050 1592
rect 3094 1588 3098 1592
rect 3294 1588 3298 1592
rect 3414 1588 3418 1592
rect 3470 1588 3474 1592
rect 3710 1588 3714 1592
rect 4070 1588 4074 1592
rect 4198 1588 4202 1592
rect 4286 1588 4290 1592
rect 518 1578 522 1582
rect 590 1578 594 1582
rect 614 1578 618 1582
rect 1406 1578 1410 1582
rect 3446 1578 3450 1582
rect 126 1568 130 1572
rect 230 1568 234 1572
rect 742 1568 746 1572
rect 782 1568 786 1572
rect 886 1568 890 1572
rect 966 1568 970 1572
rect 1894 1568 1898 1572
rect 1958 1568 1962 1572
rect 2278 1568 2282 1572
rect 2846 1568 2850 1572
rect 4166 1568 4170 1572
rect 4206 1568 4210 1572
rect 4238 1568 4242 1572
rect 4374 1568 4378 1572
rect 238 1558 242 1562
rect 294 1558 298 1562
rect 390 1558 394 1562
rect 446 1558 450 1562
rect 454 1558 458 1562
rect 486 1558 490 1562
rect 542 1558 546 1562
rect 574 1558 578 1562
rect 766 1558 770 1562
rect 990 1558 994 1562
rect 1078 1558 1082 1562
rect 1118 1558 1122 1562
rect 1142 1558 1146 1562
rect 1198 1558 1202 1562
rect 1366 1558 1370 1562
rect 1494 1558 1498 1562
rect 1574 1558 1578 1562
rect 1766 1558 1770 1562
rect 1814 1558 1818 1562
rect 1838 1558 1842 1562
rect 1878 1558 1882 1562
rect 1942 1558 1946 1562
rect 2046 1558 2050 1562
rect 2134 1558 2138 1562
rect 22 1548 26 1552
rect 62 1548 66 1552
rect 94 1547 98 1551
rect 150 1548 154 1552
rect 182 1548 186 1552
rect 254 1548 258 1552
rect 270 1548 274 1552
rect 294 1548 298 1552
rect 334 1548 338 1552
rect 374 1548 378 1552
rect 398 1548 402 1552
rect 462 1548 466 1552
rect 470 1548 474 1552
rect 558 1548 562 1552
rect 590 1548 594 1552
rect 630 1548 634 1552
rect 6 1538 10 1542
rect 86 1538 90 1542
rect 662 1547 666 1551
rect 750 1548 754 1552
rect 774 1548 778 1552
rect 790 1548 794 1552
rect 822 1547 826 1551
rect 918 1547 922 1551
rect 1158 1548 1162 1552
rect 1342 1548 1346 1552
rect 1350 1548 1354 1552
rect 1366 1548 1370 1552
rect 1390 1548 1394 1552
rect 1486 1548 1490 1552
rect 1558 1548 1562 1552
rect 1614 1548 1618 1552
rect 1638 1548 1642 1552
rect 1662 1548 1666 1552
rect 1678 1548 1682 1552
rect 1710 1548 1714 1552
rect 1758 1548 1762 1552
rect 1830 1548 1834 1552
rect 1886 1548 1890 1552
rect 1934 1548 1938 1552
rect 1958 1548 1962 1552
rect 206 1538 210 1542
rect 262 1538 266 1542
rect 270 1538 274 1542
rect 342 1538 346 1542
rect 366 1538 370 1542
rect 422 1538 426 1542
rect 502 1538 506 1542
rect 566 1538 570 1542
rect 598 1538 602 1542
rect 670 1538 674 1542
rect 806 1538 810 1542
rect 902 1538 906 1542
rect 1006 1538 1010 1542
rect 1046 1538 1050 1542
rect 1054 1538 1058 1542
rect 1118 1538 1122 1542
rect 1158 1538 1162 1542
rect 1182 1538 1186 1542
rect 1198 1538 1202 1542
rect 1214 1538 1218 1542
rect 1222 1538 1226 1542
rect 1270 1538 1274 1542
rect 1318 1538 1322 1542
rect 1342 1538 1346 1542
rect 1414 1538 1418 1542
rect 1430 1538 1434 1542
rect 1478 1538 1482 1542
rect 1510 1538 1514 1542
rect 1550 1538 1554 1542
rect 1606 1538 1610 1542
rect 1654 1538 1658 1542
rect 1670 1538 1674 1542
rect 1750 1538 1754 1542
rect 1790 1538 1794 1542
rect 1862 1538 1866 1542
rect 1926 1538 1930 1542
rect 1966 1538 1970 1542
rect 1990 1538 1994 1542
rect 2006 1548 2010 1552
rect 2022 1548 2026 1552
rect 2078 1548 2082 1552
rect 2166 1548 2170 1552
rect 2198 1548 2202 1552
rect 2294 1558 2298 1562
rect 2382 1558 2386 1562
rect 2414 1558 2418 1562
rect 2438 1558 2442 1562
rect 2478 1558 2482 1562
rect 2222 1548 2226 1552
rect 2278 1548 2282 1552
rect 2294 1548 2298 1552
rect 2318 1548 2322 1552
rect 2350 1548 2354 1552
rect 2366 1548 2370 1552
rect 2390 1548 2394 1552
rect 2470 1548 2474 1552
rect 2486 1548 2490 1552
rect 2494 1548 2498 1552
rect 2526 1558 2530 1562
rect 2590 1558 2594 1562
rect 2654 1558 2658 1562
rect 2830 1558 2834 1562
rect 2862 1558 2866 1562
rect 2574 1548 2578 1552
rect 2622 1548 2626 1552
rect 2638 1548 2642 1552
rect 2670 1548 2674 1552
rect 2726 1548 2730 1552
rect 2766 1548 2770 1552
rect 2814 1548 2818 1552
rect 2854 1548 2858 1552
rect 2886 1548 2890 1552
rect 2942 1558 2946 1562
rect 3030 1558 3034 1562
rect 3078 1558 3082 1562
rect 3150 1558 3154 1562
rect 3174 1558 3178 1562
rect 3190 1558 3194 1562
rect 2070 1538 2074 1542
rect 2102 1538 2106 1542
rect 2110 1538 2114 1542
rect 2142 1538 2146 1542
rect 2166 1538 2170 1542
rect 2190 1538 2194 1542
rect 2222 1538 2226 1542
rect 2238 1538 2242 1542
rect 2310 1538 2314 1542
rect 2318 1538 2322 1542
rect 2342 1538 2346 1542
rect 2358 1538 2362 1542
rect 2390 1538 2394 1542
rect 2454 1538 2458 1542
rect 2502 1538 2506 1542
rect 2526 1538 2530 1542
rect 2542 1538 2546 1542
rect 2606 1538 2610 1542
rect 2630 1538 2634 1542
rect 2694 1538 2698 1542
rect 2742 1538 2746 1542
rect 2790 1538 2794 1542
rect 2958 1548 2962 1552
rect 2974 1548 2978 1552
rect 3006 1548 3010 1552
rect 3046 1548 3050 1552
rect 3094 1548 3098 1552
rect 3126 1548 3130 1552
rect 3158 1548 3162 1552
rect 3166 1548 3170 1552
rect 3286 1558 3290 1562
rect 3318 1558 3322 1562
rect 3406 1558 3410 1562
rect 3422 1558 3426 1562
rect 3494 1558 3498 1562
rect 3574 1558 3578 1562
rect 3222 1548 3226 1552
rect 3238 1548 3242 1552
rect 3278 1548 3282 1552
rect 3350 1548 3354 1552
rect 3366 1548 3370 1552
rect 3390 1548 3394 1552
rect 3398 1548 3402 1552
rect 3446 1548 3450 1552
rect 3486 1548 3490 1552
rect 3526 1548 3530 1552
rect 3630 1558 3634 1562
rect 3614 1548 3618 1552
rect 3646 1548 3650 1552
rect 3662 1548 3666 1552
rect 3686 1548 3690 1552
rect 3790 1548 3794 1552
rect 3894 1558 3898 1562
rect 3926 1558 3930 1562
rect 4030 1558 4034 1562
rect 4222 1558 4226 1562
rect 4254 1558 4258 1562
rect 4294 1558 4298 1562
rect 4350 1558 4354 1562
rect 4398 1558 4402 1562
rect 4430 1558 4434 1562
rect 4470 1558 4474 1562
rect 4510 1558 4514 1562
rect 3854 1548 3858 1552
rect 3950 1548 3954 1552
rect 3982 1548 3986 1552
rect 3998 1548 4002 1552
rect 4014 1548 4018 1552
rect 4030 1548 4034 1552
rect 4078 1548 4082 1552
rect 4094 1548 4098 1552
rect 4118 1548 4122 1552
rect 4158 1548 4162 1552
rect 4190 1548 4194 1552
rect 4214 1548 4218 1552
rect 4238 1548 4242 1552
rect 4262 1548 4266 1552
rect 4310 1548 4314 1552
rect 4326 1548 4330 1552
rect 4414 1548 4418 1552
rect 4462 1548 4466 1552
rect 4470 1548 4474 1552
rect 4526 1548 4530 1552
rect 4550 1548 4554 1552
rect 4566 1548 4570 1552
rect 2910 1538 2914 1542
rect 2998 1538 3002 1542
rect 3054 1538 3058 1542
rect 3102 1538 3106 1542
rect 3134 1538 3138 1542
rect 3166 1538 3170 1542
rect 3214 1538 3218 1542
rect 3246 1538 3250 1542
rect 3270 1538 3274 1542
rect 3302 1538 3306 1542
rect 3310 1538 3314 1542
rect 3334 1538 3338 1542
rect 3422 1538 3426 1542
rect 3454 1538 3458 1542
rect 3510 1538 3514 1542
rect 3550 1538 3554 1542
rect 3558 1538 3562 1542
rect 3622 1538 3626 1542
rect 3638 1538 3642 1542
rect 3662 1538 3666 1542
rect 3710 1538 3714 1542
rect 3726 1538 3730 1542
rect 3734 1540 3738 1544
rect 3790 1538 3794 1542
rect 3806 1538 3810 1542
rect 3870 1538 3874 1542
rect 3878 1538 3882 1542
rect 3942 1538 3946 1542
rect 3974 1538 3978 1542
rect 4006 1538 4010 1542
rect 4038 1538 4042 1542
rect 4046 1538 4050 1542
rect 4134 1538 4138 1542
rect 4150 1538 4154 1542
rect 4182 1538 4186 1542
rect 4230 1538 4234 1542
rect 4270 1538 4274 1542
rect 4286 1538 4290 1542
rect 4366 1538 4370 1542
rect 4390 1538 4394 1542
rect 4406 1538 4410 1542
rect 4454 1538 4458 1542
rect 4462 1538 4466 1542
rect 4494 1538 4498 1542
rect 4510 1538 4514 1542
rect 4558 1538 4562 1542
rect 182 1528 186 1532
rect 350 1528 354 1532
rect 398 1528 402 1532
rect 414 1528 418 1532
rect 446 1528 450 1532
rect 534 1528 538 1532
rect 998 1528 1002 1532
rect 1054 1528 1058 1532
rect 1086 1528 1090 1532
rect 1134 1528 1138 1532
rect 1198 1528 1202 1532
rect 1326 1528 1330 1532
rect 1374 1528 1378 1532
rect 1398 1528 1402 1532
rect 1462 1528 1466 1532
rect 1534 1528 1538 1532
rect 1550 1528 1554 1532
rect 1694 1528 1698 1532
rect 1718 1528 1722 1532
rect 1870 1528 1874 1532
rect 1910 1528 1914 1532
rect 1974 1528 1978 1532
rect 2006 1528 2010 1532
rect 2030 1528 2034 1532
rect 2262 1528 2266 1532
rect 2278 1528 2282 1532
rect 2726 1528 2730 1532
rect 2750 1528 2754 1532
rect 2870 1528 2874 1532
rect 2910 1528 2914 1532
rect 2990 1528 2994 1532
rect 3142 1528 3146 1532
rect 3254 1528 3258 1532
rect 3262 1528 3266 1532
rect 3334 1528 3338 1532
rect 3670 1528 3674 1532
rect 3830 1528 3834 1532
rect 3918 1528 3922 1532
rect 3998 1528 4002 1532
rect 4062 1528 4066 1532
rect 4134 1528 4138 1532
rect 4166 1528 4170 1532
rect 4286 1528 4290 1532
rect 4342 1528 4346 1532
rect 4574 1528 4578 1532
rect 30 1518 34 1522
rect 190 1518 194 1522
rect 222 1518 226 1522
rect 342 1518 346 1522
rect 1030 1518 1034 1522
rect 1078 1518 1082 1522
rect 1110 1518 1114 1522
rect 1142 1518 1146 1522
rect 1246 1518 1250 1522
rect 1318 1518 1322 1522
rect 1470 1518 1474 1522
rect 1502 1518 1506 1522
rect 1630 1518 1634 1522
rect 1742 1518 1746 1522
rect 1774 1518 1778 1522
rect 1798 1518 1802 1522
rect 1918 1518 1922 1522
rect 1982 1518 1986 1522
rect 2086 1518 2090 1522
rect 2150 1518 2154 1522
rect 2174 1518 2178 1522
rect 2206 1518 2210 1522
rect 2246 1518 2250 1522
rect 2286 1518 2290 1522
rect 2342 1518 2346 1522
rect 2382 1518 2386 1522
rect 2438 1518 2442 1522
rect 2510 1518 2514 1522
rect 2590 1518 2594 1522
rect 2686 1518 2690 1522
rect 2742 1518 2746 1522
rect 2758 1518 2762 1522
rect 3022 1518 3026 1522
rect 3110 1518 3114 1522
rect 3374 1518 3378 1522
rect 3494 1518 3498 1522
rect 3598 1518 3602 1522
rect 3750 1518 3754 1522
rect 3766 1518 3770 1522
rect 3798 1518 3802 1522
rect 3822 1518 3826 1522
rect 3862 1518 3866 1522
rect 3894 1518 3898 1522
rect 3910 1518 3914 1522
rect 3926 1518 3930 1522
rect 4142 1518 4146 1522
rect 4382 1518 4386 1522
rect 4542 1518 4546 1522
rect 1002 1503 1006 1507
rect 1009 1503 1013 1507
rect 2026 1503 2030 1507
rect 2033 1503 2037 1507
rect 3050 1503 3054 1507
rect 3057 1503 3061 1507
rect 4082 1503 4086 1507
rect 4089 1503 4093 1507
rect 62 1488 66 1492
rect 166 1488 170 1492
rect 262 1488 266 1492
rect 278 1488 282 1492
rect 366 1488 370 1492
rect 382 1488 386 1492
rect 438 1488 442 1492
rect 718 1488 722 1492
rect 1126 1488 1130 1492
rect 1350 1488 1354 1492
rect 1606 1488 1610 1492
rect 1694 1488 1698 1492
rect 1886 1488 1890 1492
rect 2046 1488 2050 1492
rect 2190 1488 2194 1492
rect 2574 1488 2578 1492
rect 2622 1488 2626 1492
rect 2654 1488 2658 1492
rect 2710 1488 2714 1492
rect 2886 1488 2890 1492
rect 2966 1488 2970 1492
rect 3150 1488 3154 1492
rect 3374 1488 3378 1492
rect 3502 1488 3506 1492
rect 3646 1488 3650 1492
rect 3662 1488 3666 1492
rect 3838 1488 3842 1492
rect 4126 1488 4130 1492
rect 4198 1488 4202 1492
rect 4278 1488 4282 1492
rect 4310 1488 4314 1492
rect 4398 1488 4402 1492
rect 4534 1488 4538 1492
rect 166 1478 170 1482
rect 182 1478 186 1482
rect 30 1468 34 1472
rect 118 1468 122 1472
rect 206 1478 210 1482
rect 222 1478 226 1482
rect 310 1478 314 1482
rect 334 1478 338 1482
rect 390 1478 394 1482
rect 918 1478 922 1482
rect 926 1478 930 1482
rect 1134 1478 1138 1482
rect 1214 1478 1218 1482
rect 1222 1478 1226 1482
rect 1438 1478 1442 1482
rect 1534 1478 1538 1482
rect 1662 1478 1666 1482
rect 1742 1478 1746 1482
rect 1790 1478 1794 1482
rect 1966 1478 1970 1482
rect 2054 1478 2058 1482
rect 2126 1478 2130 1482
rect 2246 1478 2250 1482
rect 2294 1478 2298 1482
rect 2846 1478 2850 1482
rect 2934 1478 2938 1482
rect 2950 1478 2954 1482
rect 3062 1478 3066 1482
rect 3094 1478 3098 1482
rect 3110 1478 3114 1482
rect 3566 1478 3570 1482
rect 3670 1478 3674 1482
rect 3710 1478 3714 1482
rect 3718 1478 3722 1482
rect 3886 1478 3890 1482
rect 3990 1478 3994 1482
rect 3998 1478 4002 1482
rect 4006 1478 4010 1482
rect 286 1468 290 1472
rect 350 1468 354 1472
rect 398 1468 402 1472
rect 430 1468 434 1472
rect 550 1468 554 1472
rect 670 1468 674 1472
rect 758 1468 762 1472
rect 806 1468 810 1472
rect 814 1468 818 1472
rect 22 1458 26 1462
rect 46 1458 50 1462
rect 158 1458 162 1462
rect 206 1458 210 1462
rect 230 1458 234 1462
rect 286 1458 290 1462
rect 318 1458 322 1462
rect 422 1458 426 1462
rect 534 1459 538 1463
rect 566 1458 570 1462
rect 582 1458 586 1462
rect 598 1458 602 1462
rect 622 1458 626 1462
rect 654 1459 658 1463
rect 734 1458 738 1462
rect 870 1468 874 1472
rect 886 1468 890 1472
rect 958 1468 962 1472
rect 990 1468 994 1472
rect 998 1468 1002 1472
rect 1014 1468 1018 1472
rect 1070 1468 1074 1472
rect 1150 1468 1154 1472
rect 1174 1468 1178 1472
rect 1270 1468 1274 1472
rect 1286 1468 1290 1472
rect 1318 1468 1322 1472
rect 1326 1468 1330 1472
rect 1374 1468 1378 1472
rect 1382 1468 1386 1472
rect 1430 1468 1434 1472
rect 1502 1468 1506 1472
rect 1518 1468 1522 1472
rect 1550 1468 1554 1472
rect 1582 1468 1586 1472
rect 1598 1468 1602 1472
rect 1622 1468 1626 1472
rect 1654 1468 1658 1472
rect 1694 1468 1698 1472
rect 1854 1468 1858 1472
rect 1862 1468 1866 1472
rect 1942 1468 1946 1472
rect 2006 1468 2010 1472
rect 2094 1466 2098 1470
rect 2102 1468 2106 1472
rect 2158 1468 2162 1472
rect 2174 1468 2178 1472
rect 2214 1468 2218 1472
rect 2262 1468 2266 1472
rect 2302 1468 2306 1472
rect 2350 1468 2354 1472
rect 2470 1468 2474 1472
rect 878 1458 882 1462
rect 902 1458 906 1462
rect 982 1458 986 1462
rect 1046 1458 1050 1462
rect 1078 1458 1082 1462
rect 1094 1458 1098 1462
rect 1110 1458 1114 1462
rect 1182 1458 1186 1462
rect 1198 1458 1202 1462
rect 1246 1458 1250 1462
rect 1294 1458 1298 1462
rect 1310 1458 1314 1462
rect 1462 1458 1466 1462
rect 1486 1458 1490 1462
rect 1526 1458 1530 1462
rect 1558 1458 1562 1462
rect 1590 1458 1594 1462
rect 1630 1458 1634 1462
rect 1646 1458 1650 1462
rect 1686 1458 1690 1462
rect 1702 1458 1706 1462
rect 1766 1458 1770 1462
rect 1814 1458 1818 1462
rect 1902 1458 1906 1462
rect 1918 1458 1922 1462
rect 1934 1458 1938 1462
rect 1950 1458 1954 1462
rect 1966 1458 1970 1462
rect 2014 1458 2018 1462
rect 2054 1458 2058 1462
rect 2070 1458 2074 1462
rect 2078 1458 2082 1462
rect 2110 1458 2114 1462
rect 2150 1458 2154 1462
rect 2198 1458 2202 1462
rect 2222 1458 2226 1462
rect 2270 1458 2274 1462
rect 2278 1458 2282 1462
rect 2318 1458 2322 1462
rect 2342 1458 2346 1462
rect 2366 1458 2370 1462
rect 2390 1458 2394 1462
rect 2430 1458 2434 1462
rect 2454 1458 2458 1462
rect 2462 1458 2466 1462
rect 2478 1458 2482 1462
rect 2550 1468 2554 1472
rect 2598 1468 2602 1472
rect 2630 1468 2634 1472
rect 2742 1468 2746 1472
rect 2750 1468 2754 1472
rect 2766 1468 2770 1472
rect 2806 1468 2810 1472
rect 2862 1468 2866 1472
rect 2894 1468 2898 1472
rect 2950 1468 2954 1472
rect 2982 1468 2986 1472
rect 3054 1468 3058 1472
rect 3078 1468 3082 1472
rect 3118 1468 3122 1472
rect 3166 1468 3170 1472
rect 3174 1468 3178 1472
rect 3230 1468 3234 1472
rect 3246 1468 3250 1472
rect 3398 1468 3402 1472
rect 3430 1468 3434 1472
rect 3462 1468 3466 1472
rect 3510 1468 3514 1472
rect 3542 1468 3546 1472
rect 3590 1468 3594 1472
rect 3614 1468 3618 1472
rect 3622 1468 3626 1472
rect 3702 1468 3706 1472
rect 3726 1468 3730 1472
rect 3790 1468 3794 1472
rect 3798 1468 3802 1472
rect 3870 1468 3874 1472
rect 3902 1468 3906 1472
rect 3918 1468 3922 1472
rect 3950 1468 3954 1472
rect 4022 1468 4026 1472
rect 4270 1478 4274 1482
rect 4118 1468 4122 1472
rect 4134 1468 4138 1472
rect 4230 1468 4234 1472
rect 4246 1468 4250 1472
rect 4262 1468 4266 1472
rect 4286 1468 4290 1472
rect 4406 1478 4410 1482
rect 4446 1478 4450 1482
rect 4462 1478 4466 1482
rect 4326 1468 4330 1472
rect 4342 1468 4346 1472
rect 4374 1468 4378 1472
rect 4390 1468 4394 1472
rect 4414 1468 4418 1472
rect 4430 1468 4434 1472
rect 4494 1468 4498 1472
rect 4502 1468 4506 1472
rect 4526 1468 4530 1472
rect 4558 1468 4562 1472
rect 4590 1468 4594 1472
rect 2510 1458 2514 1462
rect 2654 1458 2658 1462
rect 2670 1458 2674 1462
rect 2710 1458 2714 1462
rect 2774 1458 2778 1462
rect 2798 1458 2802 1462
rect 2822 1458 2826 1462
rect 2870 1458 2874 1462
rect 2902 1458 2906 1462
rect 2926 1458 2930 1462
rect 2958 1458 2962 1462
rect 2990 1458 2994 1462
rect 3030 1458 3034 1462
rect 3086 1458 3090 1462
rect 3094 1458 3098 1462
rect 3118 1458 3122 1462
rect 3182 1458 3186 1462
rect 3198 1458 3202 1462
rect 3230 1458 3234 1462
rect 3262 1458 3266 1462
rect 3270 1458 3274 1462
rect 3278 1458 3282 1462
rect 3302 1458 3306 1462
rect 3318 1458 3322 1462
rect 3326 1458 3330 1462
rect 3350 1458 3354 1462
rect 3390 1458 3394 1462
rect 3406 1458 3410 1462
rect 3438 1458 3442 1462
rect 3454 1458 3458 1462
rect 3470 1458 3474 1462
rect 3534 1458 3538 1462
rect 3582 1458 3586 1462
rect 3630 1458 3634 1462
rect 3654 1458 3658 1462
rect 3678 1458 3682 1462
rect 3694 1458 3698 1462
rect 3734 1458 3738 1462
rect 3742 1458 3746 1462
rect 3774 1458 3778 1462
rect 3806 1458 3810 1462
rect 3862 1458 3866 1462
rect 3910 1458 3914 1462
rect 3942 1458 3946 1462
rect 3974 1458 3978 1462
rect 4014 1458 4018 1462
rect 4030 1458 4034 1462
rect 4038 1458 4042 1462
rect 4054 1458 4058 1462
rect 4062 1458 4066 1462
rect 4150 1458 4154 1462
rect 4158 1458 4162 1462
rect 4182 1458 4186 1462
rect 4230 1458 4234 1462
rect 4254 1458 4258 1462
rect 4294 1458 4298 1462
rect 4302 1458 4306 1462
rect 4334 1458 4338 1462
rect 4382 1458 4386 1462
rect 4422 1458 4426 1462
rect 4462 1458 4466 1462
rect 4478 1458 4482 1462
rect 4486 1458 4490 1462
rect 4534 1458 4538 1462
rect 4550 1458 4554 1462
rect 262 1448 266 1452
rect 270 1448 274 1452
rect 366 1448 370 1452
rect 446 1448 450 1452
rect 590 1448 594 1452
rect 614 1448 618 1452
rect 6 1438 10 1442
rect 286 1438 290 1442
rect 574 1438 578 1442
rect 894 1448 898 1452
rect 934 1448 938 1452
rect 942 1448 946 1452
rect 966 1448 970 1452
rect 982 1448 986 1452
rect 998 1448 1002 1452
rect 1038 1448 1042 1452
rect 1102 1448 1106 1452
rect 1150 1448 1154 1452
rect 1166 1448 1170 1452
rect 1182 1448 1186 1452
rect 1198 1448 1202 1452
rect 1270 1448 1274 1452
rect 1294 1448 1298 1452
rect 1486 1448 1490 1452
rect 1566 1448 1570 1452
rect 1630 1448 1634 1452
rect 1782 1448 1786 1452
rect 1838 1448 1842 1452
rect 1878 1448 1882 1452
rect 1910 1448 1914 1452
rect 1918 1448 1922 1452
rect 1974 1448 1978 1452
rect 2030 1448 2034 1452
rect 2150 1448 2154 1452
rect 2206 1448 2210 1452
rect 2318 1448 2322 1452
rect 2326 1448 2330 1452
rect 2342 1448 2346 1452
rect 2358 1448 2362 1452
rect 2534 1448 2538 1452
rect 2574 1448 2578 1452
rect 2662 1448 2666 1452
rect 2718 1448 2722 1452
rect 2726 1448 2730 1452
rect 2782 1448 2786 1452
rect 2814 1448 2818 1452
rect 2878 1448 2882 1452
rect 2974 1448 2978 1452
rect 3014 1448 3018 1452
rect 3142 1448 3146 1452
rect 3150 1448 3154 1452
rect 3198 1448 3202 1452
rect 3206 1448 3210 1452
rect 3222 1448 3226 1452
rect 3454 1448 3458 1452
rect 3486 1448 3490 1452
rect 3518 1448 3522 1452
rect 3614 1448 3618 1452
rect 3678 1448 3682 1452
rect 3774 1448 3778 1452
rect 3822 1448 3826 1452
rect 3894 1448 3898 1452
rect 3926 1448 3930 1452
rect 3958 1448 3962 1452
rect 3982 1448 3986 1452
rect 4134 1448 4138 1452
rect 4166 1448 4170 1452
rect 4174 1448 4178 1452
rect 4206 1448 4210 1452
rect 4238 1448 4242 1452
rect 4358 1448 4362 1452
rect 4438 1448 4442 1452
rect 4470 1448 4474 1452
rect 4502 1448 4506 1452
rect 4518 1448 4522 1452
rect 4566 1448 4570 1452
rect 742 1438 746 1442
rect 1046 1438 1050 1442
rect 1118 1438 1122 1442
rect 1254 1438 1258 1442
rect 1470 1438 1474 1442
rect 1582 1438 1586 1442
rect 1862 1438 1866 1442
rect 1894 1438 1898 1442
rect 2190 1438 2194 1442
rect 2222 1438 2226 1442
rect 2374 1438 2378 1442
rect 2646 1438 2650 1442
rect 2678 1438 2682 1442
rect 2702 1438 2706 1442
rect 2742 1438 2746 1442
rect 2830 1438 2834 1442
rect 2846 1438 2850 1442
rect 2990 1438 2994 1442
rect 3294 1438 3298 1442
rect 3494 1438 3498 1442
rect 3982 1438 3986 1442
rect 4190 1438 4194 1442
rect 4222 1438 4226 1442
rect 1646 1428 1650 1432
rect 2406 1428 2410 1432
rect 62 1418 66 1422
rect 462 1418 466 1422
rect 734 1418 738 1422
rect 782 1418 786 1422
rect 838 1418 842 1422
rect 910 1418 914 1422
rect 950 1418 954 1422
rect 1046 1418 1050 1422
rect 1158 1418 1162 1422
rect 1246 1418 1250 1422
rect 1398 1418 1402 1422
rect 1462 1418 1466 1422
rect 1766 1418 1770 1422
rect 1798 1418 1802 1422
rect 1814 1418 1818 1422
rect 1990 1418 1994 1422
rect 2278 1418 2282 1422
rect 2366 1418 2370 1422
rect 2446 1418 2450 1422
rect 2510 1418 2514 1422
rect 2734 1418 2738 1422
rect 2798 1418 2802 1422
rect 2822 1418 2826 1422
rect 3062 1418 3066 1422
rect 3126 1418 3130 1422
rect 3342 1418 3346 1422
rect 3406 1418 3410 1422
rect 3534 1418 3538 1422
rect 3558 1418 3562 1422
rect 3758 1418 3762 1422
rect 3782 1418 3786 1422
rect 3806 1418 3810 1422
rect 3942 1418 3946 1422
rect 4070 1418 4074 1422
rect 4574 1418 4578 1422
rect 498 1403 502 1407
rect 505 1403 509 1407
rect 1522 1403 1526 1407
rect 1529 1403 1533 1407
rect 2546 1403 2550 1407
rect 2553 1403 2557 1407
rect 3570 1403 3574 1407
rect 3577 1403 3581 1407
rect 54 1388 58 1392
rect 222 1388 226 1392
rect 438 1388 442 1392
rect 558 1388 562 1392
rect 982 1388 986 1392
rect 1326 1388 1330 1392
rect 1646 1388 1650 1392
rect 1870 1388 1874 1392
rect 1894 1388 1898 1392
rect 1974 1388 1978 1392
rect 2174 1388 2178 1392
rect 2526 1388 2530 1392
rect 2590 1388 2594 1392
rect 2646 1388 2650 1392
rect 2774 1388 2778 1392
rect 2806 1388 2810 1392
rect 2886 1388 2890 1392
rect 3014 1388 3018 1392
rect 3094 1388 3098 1392
rect 3142 1388 3146 1392
rect 3230 1388 3234 1392
rect 3430 1388 3434 1392
rect 3470 1388 3474 1392
rect 3510 1388 3514 1392
rect 3726 1388 3730 1392
rect 3814 1388 3818 1392
rect 3982 1388 3986 1392
rect 4006 1388 4010 1392
rect 4086 1388 4090 1392
rect 4198 1388 4202 1392
rect 4230 1388 4234 1392
rect 4334 1388 4338 1392
rect 4462 1388 4466 1392
rect 4526 1388 4530 1392
rect 30 1378 34 1382
rect 598 1378 602 1382
rect 3198 1378 3202 1382
rect 78 1368 82 1372
rect 214 1368 218 1372
rect 230 1368 234 1372
rect 718 1368 722 1372
rect 1174 1368 1178 1372
rect 1862 1368 1866 1372
rect 2166 1368 2170 1372
rect 2462 1368 2466 1372
rect 2582 1368 2586 1372
rect 2606 1368 2610 1372
rect 2638 1368 2642 1372
rect 2766 1368 2770 1372
rect 3134 1368 3138 1372
rect 4574 1368 4578 1372
rect 190 1358 194 1362
rect 198 1358 202 1362
rect 350 1358 354 1362
rect 22 1348 26 1352
rect 46 1348 50 1352
rect 70 1348 74 1352
rect 142 1347 146 1351
rect 206 1348 210 1352
rect 262 1348 266 1352
rect 294 1347 298 1351
rect 326 1348 330 1352
rect 374 1348 378 1352
rect 390 1358 394 1362
rect 430 1358 434 1362
rect 574 1358 578 1362
rect 582 1358 586 1362
rect 734 1358 738 1362
rect 942 1358 946 1362
rect 974 1358 978 1362
rect 1038 1358 1042 1362
rect 1102 1358 1106 1362
rect 1134 1358 1138 1362
rect 1182 1358 1186 1362
rect 1214 1358 1218 1362
rect 1238 1358 1242 1362
rect 1294 1358 1298 1362
rect 1342 1358 1346 1362
rect 1382 1358 1386 1362
rect 1390 1358 1394 1362
rect 1494 1358 1498 1362
rect 1718 1358 1722 1362
rect 1742 1358 1746 1362
rect 1798 1358 1802 1362
rect 1846 1358 1850 1362
rect 1878 1358 1882 1362
rect 470 1348 474 1352
rect 478 1348 482 1352
rect 542 1348 546 1352
rect 598 1348 602 1352
rect 678 1347 682 1351
rect 710 1348 714 1352
rect 726 1348 730 1352
rect 766 1348 770 1352
rect 926 1348 930 1352
rect 966 1348 970 1352
rect 1022 1348 1026 1352
rect 1054 1348 1058 1352
rect 1070 1348 1074 1352
rect 1086 1348 1090 1352
rect 1110 1348 1114 1352
rect 1126 1348 1130 1352
rect 1150 1348 1154 1352
rect 1182 1348 1186 1352
rect 1198 1348 1202 1352
rect 1254 1348 1258 1352
rect 1430 1348 1434 1352
rect 1494 1348 1498 1352
rect 1510 1348 1514 1352
rect 1542 1348 1546 1352
rect 1590 1348 1594 1352
rect 1662 1348 1666 1352
rect 1678 1348 1682 1352
rect 1766 1348 1770 1352
rect 1774 1348 1778 1352
rect 1830 1348 1834 1352
rect 1862 1348 1866 1352
rect 1894 1348 1898 1352
rect 1918 1358 1922 1362
rect 1990 1358 1994 1362
rect 2062 1358 2066 1362
rect 2070 1358 2074 1362
rect 2102 1358 2106 1362
rect 2110 1358 2114 1362
rect 2150 1358 2154 1362
rect 2198 1358 2202 1362
rect 1918 1348 1922 1352
rect 1934 1348 1938 1352
rect 1974 1348 1978 1352
rect 2014 1348 2018 1352
rect 2046 1348 2050 1352
rect 2142 1348 2146 1352
rect 2158 1348 2162 1352
rect 2214 1348 2218 1352
rect 2262 1358 2266 1362
rect 2334 1358 2338 1362
rect 2438 1358 2442 1362
rect 2478 1358 2482 1362
rect 2494 1358 2498 1362
rect 2566 1358 2570 1362
rect 2622 1358 2626 1362
rect 2662 1358 2666 1362
rect 2734 1358 2738 1362
rect 2782 1358 2786 1362
rect 2790 1358 2794 1362
rect 2838 1358 2842 1362
rect 2846 1358 2850 1362
rect 3062 1358 3066 1362
rect 3118 1358 3122 1362
rect 3166 1358 3170 1362
rect 3182 1358 3186 1362
rect 3262 1358 3266 1362
rect 3318 1358 3322 1362
rect 3374 1358 3378 1362
rect 3422 1358 3426 1362
rect 3566 1358 3570 1362
rect 3614 1358 3618 1362
rect 3678 1358 3682 1362
rect 3710 1358 3714 1362
rect 3758 1358 3762 1362
rect 3782 1358 3786 1362
rect 3990 1358 3994 1362
rect 4014 1358 4018 1362
rect 4142 1358 4146 1362
rect 4166 1358 4170 1362
rect 4246 1358 4250 1362
rect 4262 1358 4266 1362
rect 4374 1358 4378 1362
rect 4414 1358 4418 1362
rect 4494 1358 4498 1362
rect 2238 1348 2242 1352
rect 6 1338 10 1342
rect 134 1338 138 1342
rect 174 1338 178 1342
rect 310 1338 314 1342
rect 326 1338 330 1342
rect 358 1338 362 1342
rect 414 1338 418 1342
rect 550 1338 554 1342
rect 606 1338 610 1342
rect 670 1338 674 1342
rect 694 1338 698 1342
rect 742 1338 746 1342
rect 774 1338 778 1342
rect 838 1338 842 1342
rect 846 1338 850 1342
rect 894 1338 898 1342
rect 934 1338 938 1342
rect 990 1338 994 1342
rect 1014 1338 1018 1342
rect 1030 1338 1034 1342
rect 1062 1338 1066 1342
rect 1078 1338 1082 1342
rect 1094 1338 1098 1342
rect 1158 1338 1162 1342
rect 1230 1338 1234 1342
rect 1254 1338 1258 1342
rect 1278 1338 1282 1342
rect 1310 1338 1314 1342
rect 1358 1338 1362 1342
rect 1366 1338 1370 1342
rect 1406 1338 1410 1342
rect 1446 1338 1450 1342
rect 1502 1338 1506 1342
rect 1518 1338 1522 1342
rect 1550 1338 1554 1342
rect 1598 1338 1602 1342
rect 1670 1338 1674 1342
rect 1702 1338 1706 1342
rect 1726 1338 1730 1342
rect 1814 1338 1818 1342
rect 1822 1338 1826 1342
rect 1886 1338 1890 1342
rect 1966 1338 1970 1342
rect 2126 1338 2130 1342
rect 2142 1338 2146 1342
rect 2182 1338 2186 1342
rect 2206 1338 2210 1342
rect 2246 1338 2250 1342
rect 2262 1338 2266 1342
rect 2278 1348 2282 1352
rect 2326 1348 2330 1352
rect 2358 1348 2362 1352
rect 2390 1348 2394 1352
rect 2406 1348 2410 1352
rect 2422 1348 2426 1352
rect 2438 1348 2442 1352
rect 2470 1348 2474 1352
rect 2502 1348 2506 1352
rect 2526 1348 2530 1352
rect 2582 1348 2586 1352
rect 2614 1348 2618 1352
rect 2630 1348 2634 1352
rect 2670 1348 2674 1352
rect 2702 1348 2706 1352
rect 2710 1348 2714 1352
rect 2774 1348 2778 1352
rect 2862 1348 2866 1352
rect 2910 1348 2914 1352
rect 2942 1348 2946 1352
rect 2998 1348 3002 1352
rect 3030 1348 3034 1352
rect 3046 1348 3050 1352
rect 3110 1348 3114 1352
rect 3134 1348 3138 1352
rect 3190 1348 3194 1352
rect 3230 1348 3234 1352
rect 3254 1348 3258 1352
rect 3310 1348 3314 1352
rect 3358 1348 3362 1352
rect 3374 1348 3378 1352
rect 3414 1348 3418 1352
rect 3430 1348 3434 1352
rect 3454 1348 3458 1352
rect 3494 1348 3498 1352
rect 3518 1348 3522 1352
rect 3526 1348 3530 1352
rect 3534 1348 3538 1352
rect 3614 1348 3618 1352
rect 3638 1348 3642 1352
rect 3702 1348 3706 1352
rect 3726 1348 3730 1352
rect 3838 1348 3842 1352
rect 3846 1348 3850 1352
rect 3854 1348 3858 1352
rect 3870 1348 3874 1352
rect 3878 1348 3882 1352
rect 3894 1348 3898 1352
rect 3926 1348 3930 1352
rect 3950 1348 3954 1352
rect 3966 1348 3970 1352
rect 4022 1348 4026 1352
rect 4038 1348 4042 1352
rect 4062 1348 4066 1352
rect 4118 1348 4122 1352
rect 4174 1348 4178 1352
rect 4182 1348 4186 1352
rect 4214 1348 4218 1352
rect 4230 1348 4234 1352
rect 4254 1348 4258 1352
rect 4286 1348 4290 1352
rect 4318 1348 4322 1352
rect 4342 1348 4346 1352
rect 4350 1348 4354 1352
rect 4358 1348 4362 1352
rect 4398 1348 4402 1352
rect 4430 1348 4434 1352
rect 4454 1348 4458 1352
rect 4478 1348 4482 1352
rect 4502 1348 4506 1352
rect 4510 1348 4514 1352
rect 4518 1348 4522 1352
rect 4566 1348 4570 1352
rect 4590 1348 4594 1352
rect 4598 1348 4602 1352
rect 2318 1338 2322 1342
rect 2350 1338 2354 1342
rect 2366 1338 2370 1342
rect 2414 1338 2418 1342
rect 2446 1338 2450 1342
rect 2694 1338 2698 1342
rect 2750 1338 2754 1342
rect 2814 1338 2818 1342
rect 2822 1338 2826 1342
rect 2854 1338 2858 1342
rect 2886 1338 2890 1342
rect 2918 1338 2922 1342
rect 2950 1338 2954 1342
rect 2974 1338 2978 1342
rect 3038 1338 3042 1342
rect 3150 1338 3154 1342
rect 3262 1338 3266 1342
rect 3278 1338 3282 1342
rect 3334 1338 3338 1342
rect 3366 1338 3370 1342
rect 3390 1338 3394 1342
rect 3398 1338 3402 1342
rect 3542 1338 3546 1342
rect 3558 1338 3562 1342
rect 3606 1338 3610 1342
rect 3630 1338 3634 1342
rect 3662 1338 3666 1342
rect 3734 1338 3738 1342
rect 3742 1338 3746 1342
rect 3766 1338 3770 1342
rect 3806 1338 3810 1342
rect 3830 1338 3834 1342
rect 3974 1338 3978 1342
rect 3998 1338 4002 1342
rect 4046 1338 4050 1342
rect 4054 1338 4058 1342
rect 4150 1338 4154 1342
rect 4222 1338 4226 1342
rect 4278 1338 4282 1342
rect 4390 1338 4394 1342
rect 902 1328 906 1332
rect 950 1328 954 1332
rect 1046 1328 1050 1332
rect 1110 1328 1114 1332
rect 1126 1328 1130 1332
rect 1286 1328 1290 1332
rect 1318 1328 1322 1332
rect 1414 1328 1418 1332
rect 1582 1328 1586 1332
rect 1630 1328 1634 1332
rect 1750 1328 1754 1332
rect 1774 1328 1778 1332
rect 1790 1328 1794 1332
rect 1918 1328 1922 1332
rect 1958 1328 1962 1332
rect 1998 1328 2002 1332
rect 2014 1328 2018 1332
rect 2294 1328 2298 1332
rect 2382 1328 2386 1332
rect 2390 1328 2394 1332
rect 2406 1328 2410 1332
rect 2470 1328 2474 1332
rect 2486 1328 2490 1332
rect 2518 1328 2522 1332
rect 2542 1328 2546 1332
rect 2598 1328 2602 1332
rect 2654 1328 2658 1332
rect 2678 1328 2682 1332
rect 2726 1328 2730 1332
rect 2926 1328 2930 1332
rect 2966 1328 2970 1332
rect 3174 1328 3178 1332
rect 3206 1328 3210 1332
rect 3214 1328 3218 1332
rect 3286 1328 3290 1332
rect 3294 1328 3298 1332
rect 3446 1328 3450 1332
rect 3558 1328 3562 1332
rect 3654 1328 3658 1332
rect 3686 1328 3690 1332
rect 3694 1328 3698 1332
rect 3790 1328 3794 1332
rect 3910 1328 3914 1332
rect 3942 1328 3946 1332
rect 3966 1328 3970 1332
rect 4102 1328 4106 1332
rect 4270 1328 4274 1332
rect 4486 1328 4490 1332
rect 190 1318 194 1322
rect 430 1318 434 1322
rect 614 1318 618 1322
rect 870 1318 874 1322
rect 958 1318 962 1322
rect 1214 1318 1218 1322
rect 1238 1318 1242 1322
rect 1302 1318 1306 1322
rect 1382 1318 1386 1322
rect 1398 1318 1402 1322
rect 1558 1318 1562 1322
rect 1606 1318 1610 1322
rect 1694 1318 1698 1322
rect 1742 1318 1746 1322
rect 1758 1318 1762 1322
rect 1806 1318 1810 1322
rect 1846 1318 1850 1322
rect 1950 1318 1954 1322
rect 2062 1318 2066 1322
rect 2102 1318 2106 1322
rect 2110 1318 2114 1322
rect 2190 1318 2194 1322
rect 2230 1318 2234 1322
rect 2310 1318 2314 1322
rect 2334 1318 2338 1322
rect 2510 1318 2514 1322
rect 2686 1318 2690 1322
rect 2718 1318 2722 1322
rect 2734 1318 2738 1322
rect 2830 1318 2834 1322
rect 2958 1318 2962 1322
rect 3070 1318 3074 1322
rect 3158 1318 3162 1322
rect 3182 1318 3186 1322
rect 3246 1318 3250 1322
rect 3342 1318 3346 1322
rect 3550 1318 3554 1322
rect 3614 1318 3618 1322
rect 3646 1318 3650 1322
rect 3678 1318 3682 1322
rect 3750 1318 3754 1322
rect 3782 1318 3786 1322
rect 3934 1318 3938 1322
rect 4142 1318 4146 1322
rect 4166 1318 4170 1322
rect 4302 1318 4306 1322
rect 4446 1318 4450 1322
rect 1002 1303 1006 1307
rect 1009 1303 1013 1307
rect 2026 1303 2030 1307
rect 2033 1303 2037 1307
rect 3050 1303 3054 1307
rect 3057 1303 3061 1307
rect 4082 1303 4086 1307
rect 4089 1303 4093 1307
rect 158 1288 162 1292
rect 198 1288 202 1292
rect 294 1288 298 1292
rect 438 1288 442 1292
rect 494 1288 498 1292
rect 622 1288 626 1292
rect 862 1288 866 1292
rect 910 1288 914 1292
rect 1070 1288 1074 1292
rect 1190 1288 1194 1292
rect 1262 1288 1266 1292
rect 1414 1288 1418 1292
rect 1646 1288 1650 1292
rect 1814 1288 1818 1292
rect 1822 1288 1826 1292
rect 2150 1288 2154 1292
rect 2262 1288 2266 1292
rect 2350 1288 2354 1292
rect 2478 1288 2482 1292
rect 2526 1288 2530 1292
rect 2574 1288 2578 1292
rect 2630 1288 2634 1292
rect 2710 1288 2714 1292
rect 2758 1288 2762 1292
rect 2886 1288 2890 1292
rect 3022 1288 3026 1292
rect 3126 1288 3130 1292
rect 3190 1288 3194 1292
rect 3286 1288 3290 1292
rect 3430 1288 3434 1292
rect 3486 1288 3490 1292
rect 3702 1288 3706 1292
rect 3734 1288 3738 1292
rect 3758 1288 3762 1292
rect 3846 1288 3850 1292
rect 3998 1288 4002 1292
rect 4126 1288 4130 1292
rect 4214 1288 4218 1292
rect 4318 1288 4322 1292
rect 4550 1288 4554 1292
rect 4582 1288 4586 1292
rect 222 1278 226 1282
rect 270 1278 274 1282
rect 302 1278 306 1282
rect 326 1278 330 1282
rect 334 1278 338 1282
rect 366 1278 370 1282
rect 870 1278 874 1282
rect 942 1278 946 1282
rect 30 1268 34 1272
rect 110 1268 114 1272
rect 134 1268 138 1272
rect 150 1268 154 1272
rect 174 1268 178 1272
rect 230 1268 234 1272
rect 286 1268 290 1272
rect 326 1268 330 1272
rect 342 1268 346 1272
rect 382 1268 386 1272
rect 590 1268 594 1272
rect 702 1268 706 1272
rect 718 1268 722 1272
rect 782 1268 786 1272
rect 790 1268 794 1272
rect 838 1268 842 1272
rect 854 1268 858 1272
rect 902 1268 906 1272
rect 950 1268 954 1272
rect 1022 1268 1026 1272
rect 1046 1278 1050 1282
rect 1078 1278 1082 1282
rect 1110 1278 1114 1282
rect 1118 1278 1122 1282
rect 1286 1278 1290 1282
rect 1334 1278 1338 1282
rect 1486 1278 1490 1282
rect 1806 1278 1810 1282
rect 1870 1278 1874 1282
rect 1878 1278 1882 1282
rect 2006 1278 2010 1282
rect 2070 1278 2074 1282
rect 2110 1278 2114 1282
rect 2222 1278 2226 1282
rect 2286 1278 2290 1282
rect 2342 1278 2346 1282
rect 2390 1278 2394 1282
rect 2406 1278 2410 1282
rect 2422 1278 2426 1282
rect 2446 1278 2450 1282
rect 2622 1278 2626 1282
rect 2686 1278 2690 1282
rect 2766 1278 2770 1282
rect 2774 1278 2778 1282
rect 2862 1278 2866 1282
rect 3014 1278 3018 1282
rect 3174 1278 3178 1282
rect 3238 1278 3242 1282
rect 3278 1278 3282 1282
rect 3398 1278 3402 1282
rect 3422 1278 3426 1282
rect 1054 1268 1058 1272
rect 1078 1268 1082 1272
rect 1094 1268 1098 1272
rect 1126 1268 1130 1272
rect 1174 1268 1178 1272
rect 1198 1268 1202 1272
rect 1206 1268 1210 1272
rect 1286 1268 1290 1272
rect 1358 1268 1362 1272
rect 1366 1268 1370 1272
rect 1406 1268 1410 1272
rect 1422 1268 1426 1272
rect 1454 1268 1458 1272
rect 1462 1268 1466 1272
rect 1574 1268 1578 1272
rect 1614 1268 1618 1272
rect 1630 1268 1634 1272
rect 22 1258 26 1262
rect 118 1259 122 1263
rect 182 1258 186 1262
rect 206 1258 210 1262
rect 222 1258 226 1262
rect 254 1258 258 1262
rect 278 1258 282 1262
rect 310 1258 314 1262
rect 366 1258 370 1262
rect 422 1258 426 1262
rect 446 1258 450 1262
rect 470 1258 474 1262
rect 478 1258 482 1262
rect 542 1258 546 1262
rect 566 1258 570 1262
rect 598 1258 602 1262
rect 606 1258 610 1262
rect 678 1258 682 1262
rect 846 1258 850 1262
rect 894 1258 898 1262
rect 1022 1258 1026 1262
rect 1102 1258 1106 1262
rect 1230 1258 1234 1262
rect 1302 1258 1306 1262
rect 1310 1258 1314 1262
rect 1342 1258 1346 1262
rect 1358 1258 1362 1262
rect 1374 1258 1378 1262
rect 1398 1258 1402 1262
rect 1486 1258 1490 1262
rect 1510 1258 1514 1262
rect 1574 1258 1578 1262
rect 1606 1258 1610 1262
rect 1622 1258 1626 1262
rect 1638 1258 1642 1262
rect 1662 1258 1666 1262
rect 1710 1268 1714 1272
rect 1774 1268 1778 1272
rect 1862 1268 1866 1272
rect 1886 1268 1890 1272
rect 1918 1268 1922 1272
rect 1942 1268 1946 1272
rect 1694 1258 1698 1262
rect 1718 1258 1722 1262
rect 1734 1258 1738 1262
rect 1758 1258 1762 1262
rect 1766 1258 1770 1262
rect 1838 1258 1842 1262
rect 1854 1258 1858 1262
rect 1886 1258 1890 1262
rect 1974 1266 1978 1270
rect 2022 1268 2026 1272
rect 2102 1268 2106 1272
rect 2118 1268 2122 1272
rect 2126 1268 2130 1272
rect 2158 1268 2162 1272
rect 2190 1268 2194 1272
rect 2094 1258 2098 1262
rect 2166 1258 2170 1262
rect 2246 1266 2250 1270
rect 2254 1268 2258 1272
rect 2358 1268 2362 1272
rect 2478 1268 2482 1272
rect 2494 1268 2498 1272
rect 2542 1268 2546 1272
rect 2558 1268 2562 1272
rect 2614 1268 2618 1272
rect 2638 1268 2642 1272
rect 2686 1268 2690 1272
rect 2750 1268 2754 1272
rect 2790 1268 2794 1272
rect 2806 1268 2810 1272
rect 2870 1268 2874 1272
rect 2894 1268 2898 1272
rect 2950 1268 2954 1272
rect 2990 1268 2994 1272
rect 3006 1268 3010 1272
rect 3070 1268 3074 1272
rect 3110 1268 3114 1272
rect 3118 1268 3122 1272
rect 3166 1268 3170 1272
rect 3230 1268 3234 1272
rect 3270 1268 3274 1272
rect 3294 1268 3298 1272
rect 3334 1268 3338 1272
rect 3366 1268 3370 1272
rect 3446 1268 3450 1272
rect 3494 1268 3498 1272
rect 3798 1278 3802 1282
rect 3974 1278 3978 1282
rect 4238 1278 4242 1282
rect 4278 1278 4282 1282
rect 4542 1278 4546 1282
rect 3526 1268 3530 1272
rect 3598 1268 3602 1272
rect 3630 1268 3634 1272
rect 3662 1268 3666 1272
rect 3670 1268 3674 1272
rect 3734 1268 3738 1272
rect 3758 1268 3762 1272
rect 3774 1268 3778 1272
rect 3822 1268 3826 1272
rect 2206 1258 2210 1262
rect 2302 1258 2306 1262
rect 2318 1258 2322 1262
rect 2366 1258 2370 1262
rect 2454 1258 2458 1262
rect 2486 1258 2490 1262
rect 2646 1258 2650 1262
rect 2654 1258 2658 1262
rect 2678 1258 2682 1262
rect 2702 1258 2706 1262
rect 2726 1258 2730 1262
rect 2742 1258 2746 1262
rect 2782 1258 2786 1262
rect 2798 1258 2802 1262
rect 2806 1258 2810 1262
rect 2838 1258 2842 1262
rect 2902 1258 2906 1262
rect 2918 1258 2922 1262
rect 2950 1258 2954 1262
rect 2958 1258 2962 1262
rect 3030 1258 3034 1262
rect 3062 1258 3066 1262
rect 3102 1258 3106 1262
rect 3142 1258 3146 1262
rect 3158 1258 3162 1262
rect 3174 1258 3178 1262
rect 3222 1258 3226 1262
rect 3374 1258 3378 1262
rect 3422 1258 3426 1262
rect 3438 1258 3442 1262
rect 3470 1258 3474 1262
rect 3502 1258 3506 1262
rect 3526 1258 3530 1262
rect 3542 1258 3546 1262
rect 3590 1258 3594 1262
rect 3622 1258 3626 1262
rect 3638 1258 3642 1262
rect 3654 1258 3658 1262
rect 3678 1258 3682 1262
rect 3718 1258 3722 1262
rect 3782 1258 3786 1262
rect 3870 1268 3874 1272
rect 3878 1268 3882 1272
rect 3934 1268 3938 1272
rect 3942 1268 3946 1272
rect 4014 1266 4018 1270
rect 4022 1268 4026 1272
rect 4054 1268 4058 1272
rect 4078 1268 4082 1272
rect 4094 1268 4098 1272
rect 3902 1258 3906 1262
rect 3910 1258 3914 1262
rect 3926 1258 3930 1262
rect 3950 1258 3954 1262
rect 3974 1258 3978 1262
rect 3990 1258 3994 1262
rect 4046 1258 4050 1262
rect 4062 1258 4066 1262
rect 4110 1258 4114 1262
rect 4166 1268 4170 1272
rect 4206 1268 4210 1272
rect 4230 1268 4234 1272
rect 4310 1268 4314 1272
rect 4326 1268 4330 1272
rect 4342 1268 4346 1272
rect 4358 1268 4362 1272
rect 4374 1268 4378 1272
rect 4390 1268 4394 1272
rect 4470 1268 4474 1272
rect 4502 1268 4506 1272
rect 4518 1268 4522 1272
rect 4542 1268 4546 1272
rect 4558 1268 4562 1272
rect 4142 1258 4146 1262
rect 4270 1258 4274 1262
rect 4278 1258 4282 1262
rect 4294 1258 4298 1262
rect 4334 1258 4338 1262
rect 4382 1258 4386 1262
rect 4398 1258 4402 1262
rect 4406 1258 4410 1262
rect 4422 1258 4426 1262
rect 4430 1258 4434 1262
rect 4438 1258 4442 1262
rect 4462 1258 4466 1262
rect 4494 1258 4498 1262
rect 4534 1258 4538 1262
rect 4566 1258 4570 1262
rect 4598 1258 4602 1262
rect 166 1248 170 1252
rect 246 1248 250 1252
rect 406 1248 410 1252
rect 438 1248 442 1252
rect 550 1248 554 1252
rect 910 1248 914 1252
rect 1182 1248 1186 1252
rect 1222 1248 1226 1252
rect 1390 1248 1394 1252
rect 1438 1248 1442 1252
rect 1478 1248 1482 1252
rect 1542 1248 1546 1252
rect 1582 1248 1586 1252
rect 1646 1248 1650 1252
rect 1734 1248 1738 1252
rect 1742 1248 1746 1252
rect 1806 1248 1810 1252
rect 1822 1248 1826 1252
rect 1958 1248 1962 1252
rect 1990 1248 1994 1252
rect 2078 1248 2082 1252
rect 2094 1248 2098 1252
rect 2190 1248 2194 1252
rect 2198 1248 2202 1252
rect 2230 1248 2234 1252
rect 2262 1248 2266 1252
rect 2334 1248 2338 1252
rect 2366 1248 2370 1252
rect 2382 1248 2386 1252
rect 2510 1248 2514 1252
rect 2574 1248 2578 1252
rect 2710 1248 2714 1252
rect 2830 1248 2834 1252
rect 2862 1248 2866 1252
rect 2886 1248 2890 1252
rect 2918 1248 2922 1252
rect 2926 1248 2930 1252
rect 2942 1248 2946 1252
rect 2990 1248 2994 1252
rect 3038 1248 3042 1252
rect 3086 1248 3090 1252
rect 3134 1248 3138 1252
rect 3254 1248 3258 1252
rect 3310 1248 3314 1252
rect 3406 1248 3410 1252
rect 3478 1248 3482 1252
rect 3574 1248 3578 1252
rect 3606 1248 3610 1252
rect 3694 1248 3698 1252
rect 3734 1248 3738 1252
rect 3758 1248 3762 1252
rect 3806 1248 3810 1252
rect 3854 1248 3858 1252
rect 3910 1248 3914 1252
rect 3966 1248 3970 1252
rect 4030 1248 4034 1252
rect 4062 1248 4066 1252
rect 4158 1248 4162 1252
rect 4182 1248 4186 1252
rect 4190 1248 4194 1252
rect 4342 1248 4346 1252
rect 4446 1248 4450 1252
rect 4478 1248 4482 1252
rect 4510 1248 4514 1252
rect 6 1238 10 1242
rect 542 1238 546 1242
rect 574 1238 578 1242
rect 614 1238 618 1242
rect 878 1238 882 1242
rect 1158 1238 1162 1242
rect 1318 1238 1322 1242
rect 1454 1238 1458 1242
rect 1518 1238 1522 1242
rect 1598 1238 1602 1242
rect 1894 1238 1898 1242
rect 2214 1238 2218 1242
rect 2606 1238 2610 1242
rect 3006 1238 3010 1242
rect 3358 1238 3362 1242
rect 4494 1238 4498 1242
rect 518 1228 522 1232
rect 3622 1228 3626 1232
rect 4174 1228 4178 1232
rect 4198 1228 4202 1232
rect 566 1218 570 1222
rect 726 1218 730 1222
rect 814 1218 818 1222
rect 974 1218 978 1222
rect 1006 1218 1010 1222
rect 1326 1218 1330 1222
rect 1374 1218 1378 1222
rect 1510 1218 1514 1222
rect 1566 1218 1570 1222
rect 1758 1218 1762 1222
rect 1782 1218 1786 1222
rect 1926 1218 1930 1222
rect 2038 1218 2042 1222
rect 2134 1218 2138 1222
rect 2318 1218 2322 1222
rect 3054 1218 3058 1222
rect 3262 1218 3266 1222
rect 3382 1218 3386 1222
rect 3502 1218 3506 1222
rect 3678 1218 3682 1222
rect 3790 1218 3794 1222
rect 3950 1218 3954 1222
rect 4046 1218 4050 1222
rect 4142 1218 4146 1222
rect 4214 1218 4218 1222
rect 4254 1218 4258 1222
rect 498 1203 502 1207
rect 505 1203 509 1207
rect 1522 1203 1526 1207
rect 1529 1203 1533 1207
rect 2546 1203 2550 1207
rect 2553 1203 2557 1207
rect 3570 1203 3574 1207
rect 3577 1203 3581 1207
rect 30 1188 34 1192
rect 542 1188 546 1192
rect 710 1188 714 1192
rect 734 1188 738 1192
rect 982 1188 986 1192
rect 1142 1188 1146 1192
rect 1574 1188 1578 1192
rect 1678 1188 1682 1192
rect 1982 1188 1986 1192
rect 2118 1188 2122 1192
rect 2286 1188 2290 1192
rect 2446 1188 2450 1192
rect 2470 1188 2474 1192
rect 2518 1188 2522 1192
rect 2894 1188 2898 1192
rect 3022 1188 3026 1192
rect 3078 1188 3082 1192
rect 3166 1188 3170 1192
rect 3654 1188 3658 1192
rect 4374 1188 4378 1192
rect 4422 1188 4426 1192
rect 4510 1188 4514 1192
rect 4534 1188 4538 1192
rect 174 1178 178 1182
rect 1718 1178 1722 1182
rect 1998 1178 2002 1182
rect 4142 1178 4146 1182
rect 54 1168 58 1172
rect 78 1168 82 1172
rect 270 1168 274 1172
rect 718 1168 722 1172
rect 742 1168 746 1172
rect 886 1168 890 1172
rect 1118 1168 1122 1172
rect 1182 1168 1186 1172
rect 1270 1168 1274 1172
rect 1334 1168 1338 1172
rect 2030 1168 2034 1172
rect 2326 1168 2330 1172
rect 2470 1168 2474 1172
rect 3030 1168 3034 1172
rect 3582 1168 3586 1172
rect 3942 1168 3946 1172
rect 286 1158 290 1162
rect 294 1158 298 1162
rect 334 1158 338 1162
rect 462 1158 466 1162
rect 478 1158 482 1162
rect 558 1158 562 1162
rect 22 1148 26 1152
rect 46 1148 50 1152
rect 70 1148 74 1152
rect 110 1148 114 1152
rect 142 1147 146 1151
rect 206 1148 210 1152
rect 238 1147 242 1151
rect 406 1147 410 1151
rect 446 1148 450 1152
rect 454 1148 458 1152
rect 478 1148 482 1152
rect 542 1148 546 1152
rect 574 1148 578 1152
rect 582 1148 586 1152
rect 598 1158 602 1162
rect 646 1158 650 1162
rect 654 1158 658 1162
rect 670 1158 674 1162
rect 694 1158 698 1162
rect 758 1158 762 1162
rect 990 1158 994 1162
rect 1014 1158 1018 1162
rect 1070 1158 1074 1162
rect 1086 1158 1090 1162
rect 1102 1158 1106 1162
rect 1126 1158 1130 1162
rect 1350 1158 1354 1162
rect 1470 1158 1474 1162
rect 1478 1158 1482 1162
rect 1502 1158 1506 1162
rect 1566 1158 1570 1162
rect 1646 1158 1650 1162
rect 1774 1158 1778 1162
rect 1870 1158 1874 1162
rect 1894 1158 1898 1162
rect 1950 1158 1954 1162
rect 2134 1158 2138 1162
rect 2158 1158 2162 1162
rect 2214 1158 2218 1162
rect 2222 1158 2226 1162
rect 2254 1158 2258 1162
rect 2270 1158 2274 1162
rect 2366 1158 2370 1162
rect 2398 1158 2402 1162
rect 2438 1158 2442 1162
rect 2462 1158 2466 1162
rect 2630 1158 2634 1162
rect 2726 1158 2730 1162
rect 2862 1158 2866 1162
rect 2910 1158 2914 1162
rect 2926 1158 2930 1162
rect 3014 1158 3018 1162
rect 3054 1158 3058 1162
rect 3182 1158 3186 1162
rect 3238 1158 3242 1162
rect 3262 1158 3266 1162
rect 3294 1158 3298 1162
rect 638 1148 642 1152
rect 3398 1157 3402 1161
rect 3422 1158 3426 1162
rect 702 1148 706 1152
rect 710 1148 714 1152
rect 750 1148 754 1152
rect 790 1148 794 1152
rect 830 1148 834 1152
rect 854 1148 858 1152
rect 918 1147 922 1151
rect 1006 1148 1010 1152
rect 1038 1148 1042 1152
rect 1054 1148 1058 1152
rect 1086 1148 1090 1152
rect 1142 1148 1146 1152
rect 1238 1148 1242 1152
rect 1294 1148 1298 1152
rect 1358 1148 1362 1152
rect 1398 1148 1402 1152
rect 1422 1148 1426 1152
rect 1430 1148 1434 1152
rect 1454 1148 1458 1152
rect 1598 1148 1602 1152
rect 1670 1148 1674 1152
rect 1702 1148 1706 1152
rect 1734 1148 1738 1152
rect 1742 1148 1746 1152
rect 1766 1148 1770 1152
rect 1814 1148 1818 1152
rect 1838 1148 1842 1152
rect 1894 1148 1898 1152
rect 1910 1148 1914 1152
rect 1934 1148 1938 1152
rect 1958 1148 1962 1152
rect 3518 1158 3522 1162
rect 3550 1158 3554 1162
rect 3566 1158 3570 1162
rect 3670 1158 3674 1162
rect 3678 1158 3682 1162
rect 3694 1158 3698 1162
rect 3750 1158 3754 1162
rect 3790 1158 3794 1162
rect 3862 1158 3866 1162
rect 3902 1158 3906 1162
rect 3918 1158 3922 1162
rect 3926 1158 3930 1162
rect 3990 1158 3994 1162
rect 4070 1158 4074 1162
rect 2022 1148 2026 1152
rect 2054 1148 2058 1152
rect 6 1138 10 1142
rect 158 1138 162 1142
rect 270 1138 274 1142
rect 318 1138 322 1142
rect 398 1138 402 1142
rect 438 1138 442 1142
rect 470 1138 474 1142
rect 526 1138 530 1142
rect 566 1138 570 1142
rect 614 1138 618 1142
rect 622 1138 626 1142
rect 670 1138 674 1142
rect 766 1138 770 1142
rect 902 1138 906 1142
rect 1030 1138 1034 1142
rect 1062 1138 1066 1142
rect 1094 1138 1098 1142
rect 1118 1138 1122 1142
rect 1150 1138 1154 1142
rect 1158 1138 1162 1142
rect 1206 1138 1210 1142
rect 1214 1138 1218 1142
rect 1230 1138 1234 1142
rect 1246 1138 1250 1142
rect 1294 1138 1298 1142
rect 1318 1138 1322 1142
rect 1334 1138 1338 1142
rect 1390 1138 1394 1142
rect 1446 1138 1450 1142
rect 1494 1138 1498 1142
rect 1518 1138 1522 1142
rect 1542 1138 1546 1142
rect 1606 1138 1610 1142
rect 1662 1138 1666 1142
rect 1678 1138 1682 1142
rect 1694 1138 1698 1142
rect 1790 1138 1794 1142
rect 1806 1138 1810 1142
rect 1846 1138 1850 1142
rect 1878 1138 1882 1142
rect 1918 1138 1922 1142
rect 1926 1138 1930 1142
rect 1966 1138 1970 1142
rect 1990 1138 1994 1142
rect 2022 1138 2026 1142
rect 2086 1148 2090 1152
rect 2118 1148 2122 1152
rect 2174 1148 2178 1152
rect 2190 1148 2194 1152
rect 2214 1148 2218 1152
rect 2238 1148 2242 1152
rect 2286 1148 2290 1152
rect 2302 1148 2306 1152
rect 2334 1148 2338 1152
rect 2350 1148 2354 1152
rect 2382 1148 2386 1152
rect 2406 1148 2410 1152
rect 2430 1148 2434 1152
rect 2478 1148 2482 1152
rect 2494 1148 2498 1152
rect 2550 1148 2554 1152
rect 2582 1148 2586 1152
rect 2606 1148 2610 1152
rect 2678 1148 2682 1152
rect 2710 1148 2714 1152
rect 2790 1148 2794 1152
rect 2814 1148 2818 1152
rect 2846 1148 2850 1152
rect 2878 1148 2882 1152
rect 2926 1148 2930 1152
rect 2934 1148 2938 1152
rect 2966 1148 2970 1152
rect 2982 1148 2986 1152
rect 3038 1148 3042 1152
rect 3094 1148 3098 1152
rect 3110 1148 3114 1152
rect 3150 1148 3154 1152
rect 3230 1148 3234 1152
rect 3278 1148 3282 1152
rect 3310 1148 3314 1152
rect 3350 1148 3354 1152
rect 3382 1148 3386 1152
rect 3438 1148 3442 1152
rect 3454 1148 3458 1152
rect 3462 1148 3466 1152
rect 3470 1148 3474 1152
rect 3510 1148 3514 1152
rect 3566 1148 3570 1152
rect 3734 1148 3738 1152
rect 3758 1148 3762 1152
rect 3782 1148 3786 1152
rect 3806 1148 3810 1152
rect 3838 1148 3842 1152
rect 3870 1148 3874 1152
rect 3894 1148 3898 1152
rect 3966 1148 3970 1152
rect 4006 1148 4010 1152
rect 4014 1148 4018 1152
rect 4150 1158 4154 1162
rect 4214 1158 4218 1162
rect 4278 1158 4282 1162
rect 4310 1158 4314 1162
rect 4390 1158 4394 1162
rect 4430 1158 4434 1162
rect 4478 1158 4482 1162
rect 4526 1158 4530 1162
rect 4102 1148 4106 1152
rect 4118 1148 4122 1152
rect 4182 1148 4186 1152
rect 4198 1148 4202 1152
rect 4262 1148 4266 1152
rect 4278 1148 4282 1152
rect 4294 1148 4298 1152
rect 4318 1148 4322 1152
rect 4350 1148 4354 1152
rect 4358 1148 4362 1152
rect 4446 1148 4450 1152
rect 4462 1148 4466 1152
rect 4526 1148 4530 1152
rect 4550 1148 4554 1152
rect 4574 1148 4578 1152
rect 2110 1138 2114 1142
rect 2142 1138 2146 1142
rect 2158 1138 2162 1142
rect 2182 1138 2186 1142
rect 2198 1138 2202 1142
rect 2302 1138 2306 1142
rect 2310 1138 2314 1142
rect 2326 1138 2330 1142
rect 2342 1138 2346 1142
rect 2374 1138 2378 1142
rect 2454 1138 2458 1142
rect 2526 1138 2530 1142
rect 2646 1138 2650 1142
rect 2702 1138 2706 1142
rect 2750 1138 2754 1142
rect 2782 1138 2786 1142
rect 2886 1138 2890 1142
rect 2934 1138 2938 1142
rect 2974 1138 2978 1142
rect 2998 1138 3002 1142
rect 3070 1138 3074 1142
rect 3102 1138 3106 1142
rect 3126 1138 3130 1142
rect 3158 1138 3162 1142
rect 3182 1138 3186 1142
rect 3198 1138 3202 1142
rect 3254 1138 3258 1142
rect 3286 1138 3290 1142
rect 3302 1138 3306 1142
rect 3318 1138 3322 1142
rect 3342 1138 3346 1142
rect 3366 1138 3370 1142
rect 3414 1138 3418 1142
rect 3446 1138 3450 1142
rect 3478 1138 3482 1142
rect 3502 1138 3506 1142
rect 3534 1138 3538 1142
rect 3574 1138 3578 1142
rect 3630 1138 3634 1142
rect 3646 1138 3650 1142
rect 3678 1138 3682 1142
rect 3694 1138 3698 1142
rect 3718 1138 3722 1142
rect 3726 1138 3730 1142
rect 3846 1138 3850 1142
rect 3942 1138 3946 1142
rect 3974 1138 3978 1142
rect 4038 1138 4042 1142
rect 4078 1138 4082 1142
rect 4110 1138 4114 1142
rect 4126 1138 4130 1142
rect 4166 1138 4170 1142
rect 4174 1138 4178 1142
rect 4206 1138 4210 1142
rect 4230 1138 4234 1142
rect 4286 1138 4290 1142
rect 4318 1138 4322 1142
rect 4326 1138 4330 1142
rect 4342 1138 4346 1142
rect 4406 1138 4410 1142
rect 4438 1138 4442 1142
rect 4454 1138 4458 1142
rect 4478 1138 4482 1142
rect 4494 1138 4498 1142
rect 4502 1138 4506 1142
rect 4558 1138 4562 1142
rect 4582 1138 4586 1142
rect 526 1128 530 1132
rect 1214 1128 1218 1132
rect 1302 1128 1306 1132
rect 1358 1128 1362 1132
rect 1414 1128 1418 1132
rect 1438 1128 1442 1132
rect 1638 1128 1642 1132
rect 1838 1128 1842 1132
rect 1886 1128 1890 1132
rect 1950 1128 1954 1132
rect 1982 1128 1986 1132
rect 2062 1128 2066 1132
rect 2102 1128 2106 1132
rect 2214 1128 2218 1132
rect 2254 1128 2258 1132
rect 2414 1128 2418 1132
rect 2494 1128 2498 1132
rect 2510 1128 2514 1132
rect 2526 1128 2530 1132
rect 2598 1128 2602 1132
rect 2622 1128 2626 1132
rect 2654 1128 2658 1132
rect 2694 1128 2698 1132
rect 2726 1128 2730 1132
rect 2758 1128 2762 1132
rect 2774 1128 2778 1132
rect 2902 1128 2906 1132
rect 2942 1128 2946 1132
rect 2958 1128 2962 1132
rect 2990 1128 2994 1132
rect 3326 1128 3330 1132
rect 3334 1128 3338 1132
rect 3374 1128 3378 1132
rect 3486 1128 3490 1132
rect 3542 1128 3546 1132
rect 3622 1128 3626 1132
rect 3630 1128 3634 1132
rect 3790 1128 3794 1132
rect 3822 1128 3826 1132
rect 3886 1128 3890 1132
rect 4030 1128 4034 1132
rect 4142 1128 4146 1132
rect 4158 1128 4162 1132
rect 4238 1128 4242 1132
rect 4550 1128 4554 1132
rect 302 1118 306 1122
rect 334 1118 338 1122
rect 342 1118 346 1122
rect 654 1118 658 1122
rect 1382 1118 1386 1122
rect 1470 1118 1474 1122
rect 1478 1118 1482 1122
rect 1502 1118 1506 1122
rect 1550 1118 1554 1122
rect 1646 1118 1650 1122
rect 1870 1118 1874 1122
rect 2150 1118 2154 1122
rect 2366 1118 2370 1122
rect 2438 1118 2442 1122
rect 2566 1118 2570 1122
rect 2614 1118 2618 1122
rect 2630 1118 2634 1122
rect 2662 1118 2666 1122
rect 2734 1118 2738 1122
rect 2782 1118 2786 1122
rect 3006 1118 3010 1122
rect 3134 1118 3138 1122
rect 3238 1118 3242 1122
rect 3262 1118 3266 1122
rect 3494 1118 3498 1122
rect 3702 1118 3706 1122
rect 3750 1118 3754 1122
rect 3854 1118 3858 1122
rect 3934 1118 3938 1122
rect 4198 1118 4202 1122
rect 4214 1118 4218 1122
rect 4334 1118 4338 1122
rect 4398 1118 4402 1122
rect 4430 1118 4434 1122
rect 4486 1118 4490 1122
rect 1002 1103 1006 1107
rect 1009 1103 1013 1107
rect 2026 1103 2030 1107
rect 2033 1103 2037 1107
rect 3050 1103 3054 1107
rect 3057 1103 3061 1107
rect 4082 1103 4086 1107
rect 4089 1103 4093 1107
rect 54 1088 58 1092
rect 150 1088 154 1092
rect 414 1088 418 1092
rect 446 1088 450 1092
rect 478 1088 482 1092
rect 582 1088 586 1092
rect 678 1088 682 1092
rect 806 1088 810 1092
rect 902 1088 906 1092
rect 1038 1088 1042 1092
rect 1054 1088 1058 1092
rect 1134 1088 1138 1092
rect 1294 1088 1298 1092
rect 1302 1088 1306 1092
rect 1334 1088 1338 1092
rect 1486 1088 1490 1092
rect 1630 1088 1634 1092
rect 1758 1088 1762 1092
rect 1822 1088 1826 1092
rect 1902 1088 1906 1092
rect 1918 1088 1922 1092
rect 1974 1088 1978 1092
rect 2230 1088 2234 1092
rect 2406 1088 2410 1092
rect 2518 1088 2522 1092
rect 2558 1088 2562 1092
rect 2582 1088 2586 1092
rect 2662 1088 2666 1092
rect 2694 1088 2698 1092
rect 2702 1088 2706 1092
rect 2734 1088 2738 1092
rect 2798 1088 2802 1092
rect 2838 1088 2842 1092
rect 3086 1088 3090 1092
rect 3270 1088 3274 1092
rect 3374 1088 3378 1092
rect 3550 1088 3554 1092
rect 3686 1088 3690 1092
rect 3734 1088 3738 1092
rect 3846 1088 3850 1092
rect 3878 1088 3882 1092
rect 4126 1088 4130 1092
rect 4558 1088 4562 1092
rect 4574 1088 4578 1092
rect 270 1078 274 1082
rect 462 1078 466 1082
rect 1126 1078 1130 1082
rect 1158 1078 1162 1082
rect 1174 1078 1178 1082
rect 1262 1078 1266 1082
rect 1326 1078 1330 1082
rect 1358 1078 1362 1082
rect 1446 1078 1450 1082
rect 1526 1078 1530 1082
rect 1550 1078 1554 1082
rect 1750 1078 1754 1082
rect 1798 1078 1802 1082
rect 1870 1078 1874 1082
rect 1926 1078 1930 1082
rect 30 1068 34 1072
rect 110 1068 114 1072
rect 230 1068 234 1072
rect 254 1068 258 1072
rect 302 1068 306 1072
rect 22 1058 26 1062
rect 46 1058 50 1062
rect 118 1059 122 1063
rect 214 1059 218 1063
rect 246 1058 250 1062
rect 278 1058 282 1062
rect 294 1058 298 1062
rect 302 1058 306 1062
rect 366 1068 370 1072
rect 422 1068 426 1072
rect 486 1068 490 1072
rect 598 1068 602 1072
rect 726 1068 730 1072
rect 854 1068 858 1072
rect 910 1068 914 1072
rect 942 1068 946 1072
rect 958 1068 962 1072
rect 998 1068 1002 1072
rect 1022 1066 1026 1070
rect 1062 1068 1066 1072
rect 1070 1068 1074 1072
rect 1118 1068 1122 1072
rect 1142 1068 1146 1072
rect 1190 1068 1194 1072
rect 1222 1068 1226 1072
rect 1270 1068 1274 1072
rect 1318 1068 1322 1072
rect 1342 1068 1346 1072
rect 1406 1068 1410 1072
rect 1478 1068 1482 1072
rect 1542 1068 1546 1072
rect 1558 1068 1562 1072
rect 1582 1068 1586 1072
rect 1614 1068 1618 1072
rect 1630 1068 1634 1072
rect 1790 1068 1794 1072
rect 1894 1068 1898 1072
rect 1934 1068 1938 1072
rect 1982 1068 1986 1072
rect 318 1058 322 1062
rect 358 1058 362 1062
rect 390 1058 394 1062
rect 430 1058 434 1062
rect 526 1058 530 1062
rect 550 1058 554 1062
rect 614 1059 618 1063
rect 686 1058 690 1062
rect 694 1058 698 1062
rect 742 1059 746 1063
rect 838 1059 842 1063
rect 958 1058 962 1062
rect 990 1058 994 1062
rect 1150 1058 1154 1062
rect 1198 1058 1202 1062
rect 1230 1058 1234 1062
rect 1278 1058 1282 1062
rect 1350 1058 1354 1062
rect 1390 1058 1394 1062
rect 1446 1058 1450 1062
rect 1470 1058 1474 1062
rect 1510 1058 1514 1062
rect 1598 1058 1602 1062
rect 1606 1058 1610 1062
rect 1638 1058 1642 1062
rect 1654 1058 1658 1062
rect 1678 1058 1682 1062
rect 1686 1058 1690 1062
rect 1710 1058 1714 1062
rect 1782 1058 1786 1062
rect 1830 1058 1834 1062
rect 1854 1058 1858 1062
rect 1886 1058 1890 1062
rect 1934 1058 1938 1062
rect 2046 1078 2050 1082
rect 2174 1078 2178 1082
rect 2206 1078 2210 1082
rect 2358 1078 2362 1082
rect 2494 1078 2498 1082
rect 2638 1078 2642 1082
rect 2670 1078 2674 1082
rect 2806 1078 2810 1082
rect 2822 1078 2826 1082
rect 2910 1078 2914 1082
rect 2950 1078 2954 1082
rect 3110 1078 3114 1082
rect 3278 1078 3282 1082
rect 3310 1078 3314 1082
rect 3414 1078 3418 1082
rect 3446 1078 3450 1082
rect 3502 1078 3506 1082
rect 3526 1078 3530 1082
rect 3558 1078 3562 1082
rect 3614 1078 3618 1082
rect 3726 1078 3730 1082
rect 3814 1078 3818 1082
rect 3990 1078 3994 1082
rect 4046 1078 4050 1082
rect 4062 1078 4066 1082
rect 4086 1078 4090 1082
rect 4142 1078 4146 1082
rect 4158 1078 4162 1082
rect 4294 1078 4298 1082
rect 4406 1078 4410 1082
rect 4422 1078 4426 1082
rect 4478 1078 4482 1082
rect 2022 1068 2026 1072
rect 2086 1068 2090 1072
rect 2110 1068 2114 1072
rect 2126 1068 2130 1072
rect 2158 1068 2162 1072
rect 2190 1068 2194 1072
rect 2214 1068 2218 1072
rect 2222 1068 2226 1072
rect 2238 1068 2242 1072
rect 2254 1068 2258 1072
rect 2286 1068 2290 1072
rect 2350 1068 2354 1072
rect 2414 1068 2418 1072
rect 2486 1068 2490 1072
rect 2534 1068 2538 1072
rect 2566 1068 2570 1072
rect 2590 1068 2594 1072
rect 2654 1068 2658 1072
rect 2678 1068 2682 1072
rect 2718 1068 2722 1072
rect 2774 1068 2778 1072
rect 2782 1068 2786 1072
rect 2886 1068 2890 1072
rect 2902 1068 2906 1072
rect 2926 1068 2930 1072
rect 2998 1068 3002 1072
rect 3014 1068 3018 1072
rect 3030 1068 3034 1072
rect 3054 1068 3058 1072
rect 3118 1068 3122 1072
rect 3150 1068 3154 1072
rect 3166 1068 3170 1072
rect 3182 1068 3186 1072
rect 3190 1068 3194 1072
rect 3246 1068 3250 1072
rect 3254 1068 3258 1072
rect 3310 1068 3314 1072
rect 3350 1068 3354 1072
rect 1998 1058 2002 1062
rect 2014 1058 2018 1062
rect 2078 1058 2082 1062
rect 2142 1058 2146 1062
rect 2150 1058 2154 1062
rect 2182 1058 2186 1062
rect 2214 1058 2218 1062
rect 2246 1058 2250 1062
rect 2262 1058 2266 1062
rect 2294 1058 2298 1062
rect 2318 1058 2322 1062
rect 2350 1058 2354 1062
rect 2382 1058 2386 1062
rect 2390 1058 2394 1062
rect 2422 1058 2426 1062
rect 2478 1058 2482 1062
rect 2614 1058 2618 1062
rect 2646 1058 2650 1062
rect 2726 1058 2730 1062
rect 2766 1058 2770 1062
rect 2798 1058 2802 1062
rect 2822 1058 2826 1062
rect 2870 1058 2874 1062
rect 2918 1058 2922 1062
rect 2934 1058 2938 1062
rect 2974 1058 2978 1062
rect 2990 1058 2994 1062
rect 3022 1058 3026 1062
rect 3062 1058 3066 1062
rect 3094 1058 3098 1062
rect 3118 1058 3122 1062
rect 3158 1058 3162 1062
rect 3174 1058 3178 1062
rect 3198 1058 3202 1062
rect 3222 1058 3226 1062
rect 3238 1058 3242 1062
rect 3358 1066 3362 1070
rect 3382 1068 3386 1072
rect 3398 1068 3402 1072
rect 3438 1068 3442 1072
rect 3542 1068 3546 1072
rect 3574 1068 3578 1072
rect 3606 1068 3610 1072
rect 3638 1068 3642 1072
rect 3670 1068 3674 1072
rect 3694 1068 3698 1072
rect 3718 1068 3722 1072
rect 3782 1068 3786 1072
rect 3830 1068 3834 1072
rect 3862 1068 3866 1072
rect 3902 1068 3906 1072
rect 3910 1068 3914 1072
rect 3950 1068 3954 1072
rect 3334 1058 3338 1062
rect 3390 1058 3394 1062
rect 3438 1058 3442 1062
rect 3486 1058 3490 1062
rect 3510 1058 3514 1062
rect 3534 1058 3538 1062
rect 3646 1058 3650 1062
rect 3662 1058 3666 1062
rect 3702 1058 3706 1062
rect 3742 1058 3746 1062
rect 3750 1058 3754 1062
rect 3790 1058 3794 1062
rect 3838 1058 3842 1062
rect 3878 1058 3882 1062
rect 3894 1058 3898 1062
rect 3918 1058 3922 1062
rect 3926 1058 3930 1062
rect 4046 1068 4050 1072
rect 4062 1068 4066 1072
rect 4102 1068 4106 1072
rect 4134 1068 4138 1072
rect 4166 1068 4170 1072
rect 4222 1068 4226 1072
rect 4262 1068 4266 1072
rect 4278 1068 4282 1072
rect 4302 1068 4306 1072
rect 4334 1068 4338 1072
rect 4342 1068 4346 1072
rect 4454 1068 4458 1072
rect 4486 1068 4490 1072
rect 4518 1068 4522 1072
rect 4542 1068 4546 1072
rect 4550 1068 4554 1072
rect 3966 1058 3970 1062
rect 3982 1058 3986 1062
rect 4006 1058 4010 1062
rect 4014 1058 4018 1062
rect 4046 1058 4050 1062
rect 4590 1066 4594 1070
rect 4598 1068 4602 1072
rect 4118 1058 4122 1062
rect 4182 1058 4186 1062
rect 4206 1058 4210 1062
rect 4270 1058 4274 1062
rect 4310 1058 4314 1062
rect 4326 1058 4330 1062
rect 4350 1058 4354 1062
rect 4366 1058 4370 1062
rect 4382 1058 4386 1062
rect 4406 1058 4410 1062
rect 4422 1058 4426 1062
rect 4454 1058 4458 1062
rect 4462 1058 4466 1062
rect 4494 1058 4498 1062
rect 4510 1058 4514 1062
rect 4542 1058 4546 1062
rect 278 1048 282 1052
rect 294 1048 298 1052
rect 334 1048 338 1052
rect 398 1048 402 1052
rect 406 1048 410 1052
rect 926 1048 930 1052
rect 934 1048 938 1052
rect 1046 1048 1050 1052
rect 1174 1048 1178 1052
rect 1214 1048 1218 1052
rect 1294 1048 1298 1052
rect 1302 1048 1306 1052
rect 1430 1048 1434 1052
rect 1726 1048 1730 1052
rect 1766 1048 1770 1052
rect 1862 1048 1866 1052
rect 1958 1048 1962 1052
rect 2038 1048 2042 1052
rect 2054 1048 2058 1052
rect 2094 1048 2098 1052
rect 2102 1048 2106 1052
rect 2262 1048 2266 1052
rect 2278 1048 2282 1052
rect 2310 1048 2314 1052
rect 2342 1048 2346 1052
rect 2406 1048 2410 1052
rect 2446 1048 2450 1052
rect 2510 1048 2514 1052
rect 2550 1048 2554 1052
rect 2590 1048 2594 1052
rect 2598 1048 2602 1052
rect 2694 1048 2698 1052
rect 2702 1048 2706 1052
rect 2750 1048 2754 1052
rect 2878 1048 2882 1052
rect 2902 1048 2906 1052
rect 2974 1048 2978 1052
rect 3086 1048 3090 1052
rect 3126 1048 3130 1052
rect 3142 1048 3146 1052
rect 3214 1048 3218 1052
rect 3222 1048 3226 1052
rect 3270 1048 3274 1052
rect 3342 1048 3346 1052
rect 3406 1048 3410 1052
rect 3454 1048 3458 1052
rect 3582 1048 3586 1052
rect 3678 1048 3682 1052
rect 3702 1048 3706 1052
rect 3774 1048 3778 1052
rect 3790 1048 3794 1052
rect 3846 1048 3850 1052
rect 3934 1048 3938 1052
rect 3982 1048 3986 1052
rect 4038 1048 4042 1052
rect 4118 1048 4122 1052
rect 4238 1048 4242 1052
rect 4246 1048 4250 1052
rect 4398 1048 4402 1052
rect 4430 1048 4434 1052
rect 4526 1048 4530 1052
rect 6 1038 10 1042
rect 382 1038 386 1042
rect 694 1038 698 1042
rect 702 1038 706 1042
rect 790 1038 794 1042
rect 1390 1038 1394 1042
rect 1454 1038 1458 1042
rect 1846 1038 1850 1042
rect 1878 1038 1882 1042
rect 2862 1038 2866 1042
rect 2950 1038 2954 1042
rect 2966 1038 2970 1042
rect 3102 1038 3106 1042
rect 3334 1038 3338 1042
rect 3422 1038 3426 1042
rect 3518 1038 3522 1042
rect 3758 1038 3762 1042
rect 4214 1038 4218 1042
rect 4382 1038 4386 1042
rect 4462 1038 4466 1042
rect 358 1028 362 1032
rect 2870 1028 2874 1032
rect 4190 1028 4194 1032
rect 4294 1028 4298 1032
rect 374 1018 378 1022
rect 446 1018 450 1022
rect 918 1018 922 1022
rect 974 1018 978 1022
rect 1094 1018 1098 1022
rect 1182 1018 1186 1022
rect 1198 1018 1202 1022
rect 1230 1018 1234 1022
rect 1414 1018 1418 1022
rect 1670 1018 1674 1022
rect 1694 1018 1698 1022
rect 1782 1018 1786 1022
rect 1838 1018 1842 1022
rect 2078 1018 2082 1022
rect 2174 1018 2178 1022
rect 2422 1018 2426 1022
rect 2454 1018 2458 1022
rect 2838 1018 2842 1022
rect 2974 1018 2978 1022
rect 3014 1018 3018 1022
rect 3038 1018 3042 1022
rect 3198 1018 3202 1022
rect 3318 1018 3322 1022
rect 3470 1018 3474 1022
rect 3494 1018 3498 1022
rect 3646 1018 3650 1022
rect 3942 1018 3946 1022
rect 4150 1018 4154 1022
rect 4254 1018 4258 1022
rect 4318 1018 4322 1022
rect 4374 1018 4378 1022
rect 4494 1018 4498 1022
rect 498 1003 502 1007
rect 505 1003 509 1007
rect 1522 1003 1526 1007
rect 1529 1003 1533 1007
rect 2546 1003 2550 1007
rect 2553 1003 2557 1007
rect 3570 1003 3574 1007
rect 3577 1003 3581 1007
rect 158 988 162 992
rect 326 988 330 992
rect 422 988 426 992
rect 870 988 874 992
rect 910 988 914 992
rect 958 988 962 992
rect 1062 988 1066 992
rect 1422 988 1426 992
rect 1774 988 1778 992
rect 1886 988 1890 992
rect 1942 988 1946 992
rect 1998 988 2002 992
rect 2062 988 2066 992
rect 2102 988 2106 992
rect 2166 988 2170 992
rect 2206 988 2210 992
rect 2574 988 2578 992
rect 2638 988 2642 992
rect 2670 988 2674 992
rect 2790 988 2794 992
rect 2950 988 2954 992
rect 3262 988 3266 992
rect 3342 988 3346 992
rect 3662 988 3666 992
rect 3750 988 3754 992
rect 4006 988 4010 992
rect 4390 988 4394 992
rect 4454 988 4458 992
rect 4566 988 4570 992
rect 246 978 250 982
rect 1814 978 1818 982
rect 454 968 458 972
rect 486 968 490 972
rect 598 968 602 972
rect 654 968 658 972
rect 662 968 666 972
rect 854 968 858 972
rect 1878 968 1882 972
rect 1934 968 1938 972
rect 2054 968 2058 972
rect 2094 968 2098 972
rect 2238 968 2242 972
rect 2254 968 2258 972
rect 2374 968 2378 972
rect 2518 968 2522 972
rect 3014 968 3018 972
rect 3158 968 3162 972
rect 3398 968 3402 972
rect 3718 968 3722 972
rect 3862 968 3866 972
rect 4398 968 4402 972
rect 4462 968 4466 972
rect 4534 968 4538 972
rect 4574 968 4578 972
rect 142 958 146 962
rect 206 958 210 962
rect 310 958 314 962
rect 358 958 362 962
rect 390 958 394 962
rect 470 958 474 962
rect 502 958 506 962
rect 646 958 650 962
rect 702 958 706 962
rect 894 958 898 962
rect 926 958 930 962
rect 1014 958 1018 962
rect 1070 958 1074 962
rect 1134 958 1138 962
rect 1278 958 1282 962
rect 1318 957 1322 961
rect 1430 958 1434 962
rect 1510 958 1514 962
rect 1566 958 1570 962
rect 94 947 98 951
rect 206 948 210 952
rect 222 948 226 952
rect 294 948 298 952
rect 382 948 386 952
rect 406 948 410 952
rect 438 948 442 952
rect 446 948 450 952
rect 494 948 498 952
rect 6 938 10 942
rect 110 938 114 942
rect 126 938 130 942
rect 214 938 218 942
rect 230 938 234 942
rect 286 938 290 942
rect 310 938 314 942
rect 318 938 322 942
rect 382 938 386 942
rect 550 947 554 951
rect 638 948 642 952
rect 670 948 674 952
rect 742 948 746 952
rect 806 947 810 951
rect 918 948 922 952
rect 934 948 938 952
rect 950 948 954 952
rect 974 948 978 952
rect 1166 948 1170 952
rect 1222 948 1226 952
rect 1238 948 1242 952
rect 1358 948 1362 952
rect 1366 948 1370 952
rect 1438 948 1442 952
rect 1470 948 1474 952
rect 1486 948 1490 952
rect 1502 948 1506 952
rect 1694 958 1698 962
rect 1846 958 1850 962
rect 1894 958 1898 962
rect 1902 958 1906 962
rect 1950 958 1954 962
rect 2006 958 2010 962
rect 2070 958 2074 962
rect 2078 958 2082 962
rect 2134 958 2138 962
rect 2222 958 2226 962
rect 2294 958 2298 962
rect 2406 958 2410 962
rect 2526 958 2530 962
rect 2622 958 2626 962
rect 2822 958 2826 962
rect 2910 958 2914 962
rect 2966 958 2970 962
rect 2998 958 3002 962
rect 3142 958 3146 962
rect 3174 958 3178 962
rect 3278 958 3282 962
rect 3318 958 3322 962
rect 3326 958 3330 962
rect 3414 958 3418 962
rect 3454 958 3458 962
rect 3590 958 3594 962
rect 3630 958 3634 962
rect 3646 958 3650 962
rect 3678 958 3682 962
rect 3702 958 3706 962
rect 3734 958 3738 962
rect 3766 958 3770 962
rect 3798 958 3802 962
rect 3870 958 3874 962
rect 3910 958 3914 962
rect 1590 948 1594 952
rect 1622 948 1626 952
rect 1670 948 1674 952
rect 1686 948 1690 952
rect 1710 948 1714 952
rect 1726 948 1730 952
rect 1774 948 1778 952
rect 1790 948 1794 952
rect 1822 948 1826 952
rect 1830 948 1834 952
rect 1854 948 1858 952
rect 1886 948 1890 952
rect 1942 948 1946 952
rect 1982 948 1986 952
rect 2062 948 2066 952
rect 2094 948 2098 952
rect 2110 948 2114 952
rect 2126 948 2130 952
rect 2150 948 2154 952
rect 2190 948 2194 952
rect 2198 948 2202 952
rect 2238 948 2242 952
rect 2278 948 2282 952
rect 2294 948 2298 952
rect 2318 948 2322 952
rect 2334 948 2338 952
rect 2350 948 2354 952
rect 2382 948 2386 952
rect 2414 948 2418 952
rect 2462 948 2466 952
rect 2518 948 2522 952
rect 2566 948 2570 952
rect 2598 948 2602 952
rect 2614 948 2618 952
rect 2646 948 2650 952
rect 2670 948 2674 952
rect 2678 948 2682 952
rect 2710 948 2714 952
rect 2742 948 2746 952
rect 2774 948 2778 952
rect 446 938 450 942
rect 622 938 626 942
rect 790 938 794 942
rect 878 938 882 942
rect 950 938 954 942
rect 998 938 1002 942
rect 1078 938 1082 942
rect 1126 938 1130 942
rect 1158 938 1162 942
rect 1166 938 1170 942
rect 1214 938 1218 942
rect 1342 938 1346 942
rect 1374 938 1378 942
rect 1406 938 1410 942
rect 1446 938 1450 942
rect 1478 938 1482 942
rect 1494 938 1498 942
rect 1550 938 1554 942
rect 1654 938 1658 942
rect 1686 938 1690 942
rect 1726 938 1730 942
rect 1734 938 1738 942
rect 1782 938 1786 942
rect 1798 938 1802 942
rect 1918 938 1922 942
rect 2022 938 2026 942
rect 2830 948 2834 952
rect 2878 948 2882 952
rect 2902 948 2906 952
rect 2950 948 2954 952
rect 2990 948 2994 952
rect 3054 948 3058 952
rect 3094 948 3098 952
rect 3102 948 3106 952
rect 3166 948 3170 952
rect 3174 948 3178 952
rect 3190 948 3194 952
rect 3222 948 3226 952
rect 3254 948 3258 952
rect 3350 948 3354 952
rect 3382 948 3386 952
rect 3398 948 3402 952
rect 3430 948 3434 952
rect 3454 948 3458 952
rect 3470 948 3474 952
rect 3518 948 3522 952
rect 3542 948 3546 952
rect 3558 948 3562 952
rect 3630 948 3634 952
rect 3662 948 3666 952
rect 3718 948 3722 952
rect 3750 948 3754 952
rect 3782 948 3786 952
rect 3798 948 3802 952
rect 3830 948 3834 952
rect 3838 948 3842 952
rect 3886 948 3890 952
rect 3910 948 3914 952
rect 3934 958 3938 962
rect 3990 958 3994 962
rect 4070 958 4074 962
rect 4094 958 4098 962
rect 4142 958 4146 962
rect 4262 958 4266 962
rect 4286 958 4290 962
rect 4294 958 4298 962
rect 4374 958 4378 962
rect 4382 958 4386 962
rect 4414 958 4418 962
rect 4446 958 4450 962
rect 4478 958 4482 962
rect 4558 958 4562 962
rect 3982 948 3986 952
rect 4006 948 4010 952
rect 4014 948 4018 952
rect 4054 948 4058 952
rect 4070 948 4074 952
rect 4126 948 4130 952
rect 4174 948 4178 952
rect 4182 948 4186 952
rect 4246 948 4250 952
rect 4286 948 4290 952
rect 4342 948 4346 952
rect 4358 948 4362 952
rect 4390 948 4394 952
rect 4438 948 4442 952
rect 4454 948 4458 952
rect 4478 948 4482 952
rect 4494 948 4498 952
rect 4510 948 4514 952
rect 4566 948 4570 952
rect 2166 938 2170 942
rect 2182 938 2186 942
rect 2230 938 2234 942
rect 2246 938 2250 942
rect 2270 938 2274 942
rect 2302 938 2306 942
rect 2310 938 2314 942
rect 2342 938 2346 942
rect 2358 938 2362 942
rect 2382 938 2386 942
rect 2422 938 2426 942
rect 2454 938 2458 942
rect 2478 938 2482 942
rect 2502 938 2506 942
rect 2534 938 2538 942
rect 2550 938 2554 942
rect 2582 938 2586 942
rect 2606 938 2610 942
rect 2646 938 2650 942
rect 2750 938 2754 942
rect 2766 938 2770 942
rect 2798 938 2802 942
rect 2806 938 2810 942
rect 2822 938 2826 942
rect 2870 938 2874 942
rect 2886 938 2890 942
rect 2926 938 2930 942
rect 2958 938 2962 942
rect 2982 938 2986 942
rect 3030 938 3034 942
rect 3046 938 3050 942
rect 3110 938 3114 942
rect 3126 938 3130 942
rect 3166 938 3170 942
rect 3198 938 3202 942
rect 3222 938 3226 942
rect 3270 938 3274 942
rect 3302 938 3306 942
rect 3350 938 3354 942
rect 3358 938 3362 942
rect 3390 938 3394 942
rect 3422 938 3426 942
rect 3478 938 3482 942
rect 3494 938 3498 942
rect 3534 938 3538 942
rect 3550 938 3554 942
rect 3622 938 3626 942
rect 3654 938 3658 942
rect 3686 938 3690 942
rect 3710 938 3714 942
rect 3742 938 3746 942
rect 3774 938 3778 942
rect 3830 938 3834 942
rect 3846 938 3850 942
rect 3894 938 3898 942
rect 3902 938 3906 942
rect 3950 938 3954 942
rect 4022 938 4026 942
rect 4086 938 4090 942
rect 4118 938 4122 942
rect 4150 938 4154 942
rect 4190 938 4194 942
rect 4230 938 4234 942
rect 4238 938 4242 942
rect 4302 938 4306 942
rect 4318 938 4322 942
rect 4430 938 4434 942
rect 4502 938 4506 942
rect 94 928 98 932
rect 166 928 170 932
rect 190 928 194 932
rect 278 928 282 932
rect 494 928 498 932
rect 550 928 554 932
rect 974 928 978 932
rect 990 928 994 932
rect 1038 928 1042 932
rect 1222 928 1226 932
rect 1246 928 1250 932
rect 1286 928 1290 932
rect 1310 928 1314 932
rect 1334 928 1338 932
rect 1406 928 1410 932
rect 1462 928 1466 932
rect 1614 928 1618 932
rect 1750 928 1754 932
rect 1814 928 1818 932
rect 1990 928 1994 932
rect 2166 928 2170 932
rect 2214 928 2218 932
rect 2262 928 2266 932
rect 2406 928 2410 932
rect 2430 928 2434 932
rect 2438 928 2442 932
rect 2446 928 2450 932
rect 2486 928 2490 932
rect 2502 928 2506 932
rect 2590 928 2594 932
rect 2654 928 2658 932
rect 2670 928 2674 932
rect 2694 928 2698 932
rect 2782 928 2786 932
rect 2846 928 2850 932
rect 2854 928 2858 932
rect 2862 928 2866 932
rect 2886 928 2890 932
rect 2966 928 2970 932
rect 3030 928 3034 932
rect 3110 928 3114 932
rect 3206 928 3210 932
rect 3230 928 3234 932
rect 3286 928 3290 932
rect 3454 928 3458 932
rect 3486 928 3490 932
rect 3590 928 3594 932
rect 3614 928 3618 932
rect 3694 928 3698 932
rect 3806 928 3810 932
rect 4038 928 4042 932
rect 4206 928 4210 932
rect 4326 928 4330 932
rect 4414 928 4418 932
rect 4526 928 4530 932
rect 4550 928 4554 932
rect 182 918 186 922
rect 358 918 362 922
rect 390 918 394 922
rect 614 918 618 922
rect 886 918 890 922
rect 982 918 986 922
rect 1030 918 1034 922
rect 1102 918 1106 922
rect 1134 918 1138 922
rect 1190 918 1194 922
rect 1270 918 1274 922
rect 1382 918 1386 922
rect 1454 918 1458 922
rect 1518 918 1522 922
rect 1574 918 1578 922
rect 1638 918 1642 922
rect 1694 918 1698 922
rect 1910 918 1914 922
rect 1966 918 1970 922
rect 2006 918 2010 922
rect 2118 918 2122 922
rect 2318 918 2322 922
rect 2758 918 2762 922
rect 2838 918 2842 922
rect 3078 918 3082 922
rect 3238 918 3242 922
rect 3318 918 3322 922
rect 3814 918 3818 922
rect 3966 918 3970 922
rect 4142 918 4146 922
rect 4198 918 4202 922
rect 4222 918 4226 922
rect 4374 918 4378 922
rect 1002 903 1006 907
rect 1009 903 1013 907
rect 2026 903 2030 907
rect 2033 903 2037 907
rect 3050 903 3054 907
rect 3057 903 3061 907
rect 4082 903 4086 907
rect 4089 903 4093 907
rect 230 888 234 892
rect 262 888 266 892
rect 446 888 450 892
rect 678 888 682 892
rect 878 888 882 892
rect 1046 888 1050 892
rect 1118 888 1122 892
rect 1182 888 1186 892
rect 1214 888 1218 892
rect 1246 888 1250 892
rect 1262 888 1266 892
rect 1566 888 1570 892
rect 1590 888 1594 892
rect 1766 888 1770 892
rect 1870 888 1874 892
rect 1966 888 1970 892
rect 1998 888 2002 892
rect 2014 888 2018 892
rect 2078 888 2082 892
rect 2094 888 2098 892
rect 2150 888 2154 892
rect 2446 888 2450 892
rect 2534 888 2538 892
rect 2662 888 2666 892
rect 2694 888 2698 892
rect 2718 888 2722 892
rect 2966 888 2970 892
rect 3070 888 3074 892
rect 3118 888 3122 892
rect 3190 888 3194 892
rect 3262 888 3266 892
rect 3294 888 3298 892
rect 3334 888 3338 892
rect 3406 888 3410 892
rect 3526 888 3530 892
rect 3614 888 3618 892
rect 3622 888 3626 892
rect 3694 888 3698 892
rect 3742 888 3746 892
rect 3782 888 3786 892
rect 3806 888 3810 892
rect 3990 888 3994 892
rect 4038 888 4042 892
rect 4174 888 4178 892
rect 4446 888 4450 892
rect 4478 888 4482 892
rect 4550 888 4554 892
rect 270 878 274 882
rect 1142 878 1146 882
rect 1206 878 1210 882
rect 1470 878 1474 882
rect 1558 878 1562 882
rect 1598 878 1602 882
rect 1678 878 1682 882
rect 1758 878 1762 882
rect 1798 878 1802 882
rect 1854 878 1858 882
rect 1902 878 1906 882
rect 1934 878 1938 882
rect 1958 878 1962 882
rect 2006 878 2010 882
rect 2142 878 2146 882
rect 2174 878 2178 882
rect 2230 878 2234 882
rect 2246 878 2250 882
rect 2278 878 2282 882
rect 2470 878 2474 882
rect 2686 878 2690 882
rect 2766 878 2770 882
rect 2830 878 2834 882
rect 2942 878 2946 882
rect 3038 878 3042 882
rect 3462 878 3466 882
rect 3518 878 3522 882
rect 3670 878 3674 882
rect 3734 878 3738 882
rect 3750 878 3754 882
rect 3774 878 3778 882
rect 3958 878 3962 882
rect 4150 878 4154 882
rect 4182 878 4186 882
rect 4238 878 4242 882
rect 4246 878 4250 882
rect 4278 878 4282 882
rect 4302 878 4306 882
rect 4486 878 4490 882
rect 4518 878 4522 882
rect 4558 878 4562 882
rect 6 868 10 872
rect 30 868 34 872
rect 94 868 98 872
rect 134 868 138 872
rect 150 868 154 872
rect 214 868 218 872
rect 222 868 226 872
rect 238 868 242 872
rect 254 868 258 872
rect 286 868 290 872
rect 438 868 442 872
rect 550 868 554 872
rect 598 868 602 872
rect 750 868 754 872
rect 798 868 802 872
rect 886 868 890 872
rect 934 868 938 872
rect 950 868 954 872
rect 1054 868 1058 872
rect 1110 868 1114 872
rect 1150 868 1154 872
rect 1166 868 1170 872
rect 1198 868 1202 872
rect 1222 868 1226 872
rect 1238 868 1242 872
rect 1278 868 1282 872
rect 1286 868 1290 872
rect 1302 868 1306 872
rect 1318 868 1322 872
rect 1350 868 1354 872
rect 1398 868 1402 872
rect 1430 868 1434 872
rect 1462 868 1466 872
rect 1478 868 1482 872
rect 1534 868 1538 872
rect 1574 868 1578 872
rect 1614 868 1618 872
rect 1630 868 1634 872
rect 1646 868 1650 872
rect 1734 868 1738 872
rect 1750 868 1754 872
rect 1894 868 1898 872
rect 1910 868 1914 872
rect 1934 868 1938 872
rect 1974 868 1978 872
rect 2030 868 2034 872
rect 2046 868 2050 872
rect 22 858 26 862
rect 118 859 122 863
rect 246 858 250 862
rect 302 859 306 863
rect 382 858 386 862
rect 478 858 482 862
rect 510 859 514 863
rect 566 858 570 862
rect 622 858 626 862
rect 694 858 698 862
rect 718 858 722 862
rect 726 858 730 862
rect 814 859 818 863
rect 966 859 970 863
rect 1174 858 1178 862
rect 1230 858 1234 862
rect 1294 858 1298 862
rect 1326 858 1330 862
rect 1350 858 1354 862
rect 1422 858 1426 862
rect 1454 858 1458 862
rect 1478 858 1482 862
rect 1582 858 1586 862
rect 1606 858 1610 862
rect 1622 858 1626 862
rect 1638 858 1642 862
rect 1670 858 1674 862
rect 1702 858 1706 862
rect 1742 858 1746 862
rect 1782 858 1786 862
rect 1814 858 1818 862
rect 1838 858 1842 862
rect 1846 858 1850 862
rect 1886 858 1890 862
rect 1950 858 1954 862
rect 2062 866 2066 870
rect 2086 868 2090 872
rect 2110 868 2114 872
rect 2174 868 2178 872
rect 2190 868 2194 872
rect 2214 868 2218 872
rect 2230 868 2234 872
rect 2254 868 2258 872
rect 2278 868 2282 872
rect 2318 868 2322 872
rect 2350 868 2354 872
rect 2382 868 2386 872
rect 2398 868 2402 872
rect 2430 868 2434 872
rect 2454 868 2458 872
rect 2486 868 2490 872
rect 2502 868 2506 872
rect 2518 868 2522 872
rect 2550 868 2554 872
rect 2582 868 2586 872
rect 2598 868 2602 872
rect 2630 868 2634 872
rect 2678 868 2682 872
rect 2742 868 2746 872
rect 2774 868 2778 872
rect 2806 868 2810 872
rect 2846 868 2850 872
rect 2878 868 2882 872
rect 2926 868 2930 872
rect 3030 868 3034 872
rect 3046 868 3050 872
rect 3078 868 3082 872
rect 3142 868 3146 872
rect 3166 868 3170 872
rect 3230 868 3234 872
rect 3238 868 3242 872
rect 3270 868 3274 872
rect 3302 868 3306 872
rect 3358 868 3362 872
rect 3390 868 3394 872
rect 3414 868 3418 872
rect 3446 868 3450 872
rect 3534 868 3538 872
rect 3566 868 3570 872
rect 3590 868 3594 872
rect 3646 868 3650 872
rect 3678 868 3682 872
rect 3702 868 3706 872
rect 3798 868 3802 872
rect 3822 868 3826 872
rect 3862 868 3866 872
rect 3870 868 3874 872
rect 3942 868 3946 872
rect 3982 868 3986 872
rect 1990 858 1994 862
rect 2102 858 2106 862
rect 2166 858 2170 862
rect 2182 858 2186 862
rect 2198 858 2202 862
rect 2206 858 2210 862
rect 2254 858 2258 862
rect 2302 858 2306 862
rect 2310 858 2314 862
rect 2358 858 2362 862
rect 2374 858 2378 862
rect 2462 858 2466 862
rect 2494 858 2498 862
rect 2510 858 2514 862
rect 2606 858 2610 862
rect 2702 858 2706 862
rect 2726 858 2730 862
rect 2750 858 2754 862
rect 2782 858 2786 862
rect 2838 858 2842 862
rect 2854 858 2858 862
rect 2910 858 2914 862
rect 2918 858 2922 862
rect 2950 858 2954 862
rect 2958 858 2962 862
rect 2982 858 2986 862
rect 3006 858 3010 862
rect 3094 858 3098 862
rect 3110 858 3114 862
rect 3134 858 3138 862
rect 3174 858 3178 862
rect 3222 858 3226 862
rect 3246 858 3250 862
rect 3278 858 3282 862
rect 3310 858 3314 862
rect 3350 858 3354 862
rect 3382 858 3386 862
rect 3438 858 3442 862
rect 3478 858 3482 862
rect 3510 858 3514 862
rect 3542 858 3546 862
rect 3566 858 3570 862
rect 3638 858 3642 862
rect 3654 858 3658 862
rect 3726 858 3730 862
rect 3758 858 3762 862
rect 3830 858 3834 862
rect 3838 858 3842 862
rect 3862 858 3866 862
rect 3886 858 3890 862
rect 3934 858 3938 862
rect 3982 858 3986 862
rect 4014 868 4018 872
rect 4046 868 4050 872
rect 4102 868 4106 872
rect 4126 868 4130 872
rect 4134 868 4138 872
rect 4166 868 4170 872
rect 4190 868 4194 872
rect 4206 868 4210 872
rect 4270 868 4274 872
rect 4326 868 4330 872
rect 4334 868 4338 872
rect 4374 868 4378 872
rect 4414 868 4418 872
rect 4422 868 4426 872
rect 4438 868 4442 872
rect 4454 868 4458 872
rect 4502 868 4506 872
rect 4558 868 4562 872
rect 4582 868 4586 872
rect 4022 858 4026 862
rect 4054 858 4058 862
rect 4086 858 4090 862
rect 4110 858 4114 862
rect 4126 858 4130 862
rect 4158 858 4162 862
rect 4198 858 4202 862
rect 4214 858 4218 862
rect 4262 858 4266 862
rect 4294 858 4298 862
rect 4318 858 4322 862
rect 4326 858 4330 862
rect 4406 858 4410 862
rect 4438 858 4442 862
rect 4462 858 4466 862
rect 4510 858 4514 862
rect 4534 858 4538 862
rect 4574 858 4578 862
rect 238 848 242 852
rect 542 848 546 852
rect 558 848 562 852
rect 366 838 370 842
rect 550 838 554 842
rect 574 838 578 842
rect 1182 848 1186 852
rect 1262 848 1266 852
rect 1310 848 1314 852
rect 1342 848 1346 852
rect 1406 848 1410 852
rect 1438 848 1442 852
rect 1718 848 1722 852
rect 1726 848 1730 852
rect 2014 848 2018 852
rect 2102 848 2106 852
rect 2134 848 2138 852
rect 2230 848 2234 852
rect 2286 848 2290 852
rect 2342 848 2346 852
rect 2374 848 2378 852
rect 2382 848 2386 852
rect 2422 848 2426 852
rect 2526 848 2530 852
rect 2534 848 2538 852
rect 2614 848 2618 852
rect 2630 848 2634 852
rect 2638 848 2642 852
rect 2662 848 2666 852
rect 2734 848 2738 852
rect 2766 848 2770 852
rect 2822 848 2826 852
rect 2862 848 2866 852
rect 2998 848 3002 852
rect 3062 848 3066 852
rect 3110 848 3114 852
rect 3118 848 3122 852
rect 3150 848 3154 852
rect 3166 848 3170 852
rect 3206 848 3210 852
rect 3262 848 3266 852
rect 3294 848 3298 852
rect 3326 848 3330 852
rect 3366 848 3370 852
rect 3382 848 3386 852
rect 3398 848 3402 852
rect 3422 848 3426 852
rect 3494 848 3498 852
rect 3550 848 3554 852
rect 3574 848 3578 852
rect 3614 848 3618 852
rect 3622 848 3626 852
rect 3662 848 3666 852
rect 3694 848 3698 852
rect 3726 848 3730 852
rect 3782 848 3786 852
rect 3806 848 3810 852
rect 3886 848 3890 852
rect 3910 848 3914 852
rect 3966 848 3970 852
rect 3990 848 3994 852
rect 4038 848 4042 852
rect 4070 848 4074 852
rect 4078 848 4082 852
rect 4150 848 4154 852
rect 4214 848 4218 852
rect 4246 848 4250 852
rect 4390 848 4394 852
rect 4590 848 4594 852
rect 702 838 706 842
rect 726 838 730 842
rect 734 838 738 842
rect 1950 838 1954 842
rect 2470 838 2474 842
rect 2718 838 2722 842
rect 3014 838 3018 842
rect 3222 838 3226 842
rect 3758 838 3762 842
rect 3958 838 3962 842
rect 4222 838 4226 842
rect 694 828 698 832
rect 2278 828 2282 832
rect 3438 828 3442 832
rect 758 818 762 822
rect 910 818 914 822
rect 1078 818 1082 822
rect 1366 818 1370 822
rect 1422 818 1426 822
rect 1454 818 1458 822
rect 1502 818 1506 822
rect 1702 818 1706 822
rect 1822 818 1826 822
rect 2118 818 2122 822
rect 2326 818 2330 822
rect 2582 818 2586 822
rect 2646 818 2650 822
rect 2782 818 2786 822
rect 2870 818 2874 822
rect 2894 818 2898 822
rect 2942 818 2946 822
rect 3006 818 3010 822
rect 3134 818 3138 822
rect 4286 818 4290 822
rect 4350 818 4354 822
rect 498 803 502 807
rect 505 803 509 807
rect 1522 803 1526 807
rect 1529 803 1533 807
rect 2546 803 2550 807
rect 2553 803 2557 807
rect 3570 803 3574 807
rect 3577 803 3581 807
rect 318 788 322 792
rect 1238 788 1242 792
rect 1694 788 1698 792
rect 1814 788 1818 792
rect 1894 788 1898 792
rect 2086 788 2090 792
rect 2102 788 2106 792
rect 2134 788 2138 792
rect 2198 788 2202 792
rect 2246 788 2250 792
rect 2310 788 2314 792
rect 2830 788 2834 792
rect 3086 788 3090 792
rect 3238 788 3242 792
rect 3254 788 3258 792
rect 3414 788 3418 792
rect 3550 788 3554 792
rect 3654 788 3658 792
rect 3718 788 3722 792
rect 3838 788 3842 792
rect 3870 788 3874 792
rect 3902 788 3906 792
rect 3982 788 3986 792
rect 4238 788 4242 792
rect 4326 788 4330 792
rect 4430 788 4434 792
rect 4518 788 4522 792
rect 566 778 570 782
rect 2382 778 2386 782
rect 2582 778 2586 782
rect 302 768 306 772
rect 326 768 330 772
rect 1350 768 1354 772
rect 1886 768 1890 772
rect 2006 768 2010 772
rect 2590 768 2594 772
rect 2934 768 2938 772
rect 3846 768 3850 772
rect 3998 768 4002 772
rect 4110 768 4114 772
rect 4198 768 4202 772
rect 4222 768 4226 772
rect 4230 768 4234 772
rect 4262 768 4266 772
rect 4350 768 4354 772
rect 4382 768 4386 772
rect 134 758 138 762
rect 150 758 154 762
rect 222 758 226 762
rect 278 758 282 762
rect 70 747 74 751
rect 134 748 138 752
rect 166 748 170 752
rect 182 748 186 752
rect 222 748 226 752
rect 254 748 258 752
rect 262 748 266 752
rect 342 758 346 762
rect 302 748 306 752
rect 334 748 338 752
rect 358 748 362 752
rect 382 758 386 762
rect 558 758 562 762
rect 574 758 578 762
rect 638 758 642 762
rect 678 758 682 762
rect 750 758 754 762
rect 774 758 778 762
rect 414 748 418 752
rect 446 748 450 752
rect 470 748 474 752
rect 478 748 482 752
rect 534 748 538 752
rect 622 748 626 752
rect 630 748 634 752
rect 646 748 650 752
rect 678 748 682 752
rect 702 748 706 752
rect 734 748 738 752
rect 142 738 146 742
rect 174 738 178 742
rect 198 738 202 742
rect 310 738 314 742
rect 350 738 354 742
rect 406 738 410 742
rect 494 738 498 742
rect 558 738 562 742
rect 574 738 578 742
rect 694 738 698 742
rect 870 747 874 751
rect 950 748 954 752
rect 1174 748 1178 752
rect 1222 758 1226 762
rect 1342 758 1346 762
rect 1366 758 1370 762
rect 1430 758 1434 762
rect 1454 758 1458 762
rect 1470 758 1474 762
rect 1654 758 1658 762
rect 1710 758 1714 762
rect 1750 758 1754 762
rect 1798 758 1802 762
rect 1870 758 1874 762
rect 1902 758 1906 762
rect 1990 758 1994 762
rect 2014 758 2018 762
rect 2070 758 2074 762
rect 2118 758 2122 762
rect 2214 758 2218 762
rect 2318 758 2322 762
rect 2446 758 2450 762
rect 2534 758 2538 762
rect 2566 758 2570 762
rect 2694 758 2698 762
rect 2798 758 2802 762
rect 2814 758 2818 762
rect 2846 758 2850 762
rect 2910 758 2914 762
rect 2966 758 2970 762
rect 2990 758 2994 762
rect 3102 758 3106 762
rect 3142 758 3146 762
rect 3166 758 3170 762
rect 3174 758 3178 762
rect 3198 758 3202 762
rect 3230 758 3234 762
rect 3294 758 3298 762
rect 3382 758 3386 762
rect 1206 748 1210 752
rect 1230 748 1234 752
rect 1246 748 1250 752
rect 1470 748 1474 752
rect 1566 748 1570 752
rect 1606 748 1610 752
rect 1694 748 1698 752
rect 1718 748 1722 752
rect 1758 748 1762 752
rect 1774 748 1778 752
rect 1790 748 1794 752
rect 1814 748 1818 752
rect 1830 748 1834 752
rect 1846 748 1850 752
rect 1878 748 1882 752
rect 1918 748 1922 752
rect 1958 748 1962 752
rect 1966 748 1970 752
rect 2102 748 2106 752
rect 2134 748 2138 752
rect 2182 748 2186 752
rect 2190 748 2194 752
rect 2222 748 2226 752
rect 2254 748 2258 752
rect 2262 748 2266 752
rect 2286 748 2290 752
rect 2390 748 2394 752
rect 2406 748 2410 752
rect 2430 748 2434 752
rect 2478 748 2482 752
rect 2486 748 2490 752
rect 2494 748 2498 752
rect 2518 748 2522 752
rect 2582 748 2586 752
rect 2654 748 2658 752
rect 2670 748 2674 752
rect 2694 748 2698 752
rect 2734 748 2738 752
rect 2790 748 2794 752
rect 2830 748 2834 752
rect 2854 748 2858 752
rect 2894 748 2898 752
rect 2934 748 2938 752
rect 758 738 762 742
rect 1062 738 1066 742
rect 3022 748 3026 752
rect 3054 748 3058 752
rect 3102 748 3106 752
rect 3190 748 3194 752
rect 3222 748 3226 752
rect 3278 748 3282 752
rect 3302 748 3306 752
rect 3310 748 3314 752
rect 3334 748 3338 752
rect 3342 748 3346 752
rect 3422 748 3426 752
rect 3430 748 3434 752
rect 3438 748 3442 752
rect 3462 748 3466 752
rect 3486 748 3490 752
rect 3494 748 3498 752
rect 3510 758 3514 762
rect 3534 758 3538 762
rect 3598 758 3602 762
rect 3758 758 3762 762
rect 3614 748 3618 752
rect 3686 748 3690 752
rect 3702 748 3706 752
rect 3726 748 3730 752
rect 3734 748 3738 752
rect 3830 758 3834 762
rect 4006 758 4010 762
rect 4214 758 4218 762
rect 4246 758 4250 762
rect 4294 758 4298 762
rect 4350 758 4354 762
rect 4414 758 4418 762
rect 4470 758 4474 762
rect 3782 748 3786 752
rect 3822 748 3826 752
rect 3846 748 3850 752
rect 3942 748 3946 752
rect 3950 748 3954 752
rect 3998 748 4002 752
rect 4014 748 4018 752
rect 4030 748 4034 752
rect 4046 748 4050 752
rect 4110 748 4114 752
rect 4158 748 4162 752
rect 4190 748 4194 752
rect 4222 748 4226 752
rect 4262 748 4266 752
rect 4286 748 4290 752
rect 4310 748 4314 752
rect 4342 748 4346 752
rect 4358 748 4362 752
rect 4406 748 4410 752
rect 4430 748 4434 752
rect 4454 748 4458 752
rect 4470 748 4474 752
rect 4478 748 4482 752
rect 4542 748 4546 752
rect 1086 738 1090 742
rect 1094 738 1098 742
rect 1142 738 1146 742
rect 1150 738 1154 742
rect 1166 738 1170 742
rect 1182 738 1186 742
rect 1198 738 1202 742
rect 1254 738 1258 742
rect 1270 738 1274 742
rect 1326 738 1330 742
rect 1342 738 1346 742
rect 1374 738 1378 742
rect 1422 738 1426 742
rect 1446 738 1450 742
rect 1478 738 1482 742
rect 1574 738 1578 742
rect 1614 738 1618 742
rect 1638 738 1642 742
rect 1686 738 1690 742
rect 1782 738 1786 742
rect 1822 738 1826 742
rect 1854 738 1858 742
rect 1926 738 1930 742
rect 1934 738 1938 742
rect 2006 738 2010 742
rect 2030 738 2034 742
rect 2054 738 2058 742
rect 2094 738 2098 742
rect 2126 738 2130 742
rect 2174 738 2178 742
rect 2190 738 2194 742
rect 2230 738 2234 742
rect 2286 738 2290 742
rect 2294 738 2298 742
rect 2334 738 2338 742
rect 2358 738 2362 742
rect 2366 738 2370 742
rect 2398 738 2402 742
rect 2470 738 2474 742
rect 2550 738 2554 742
rect 2614 738 2618 742
rect 2646 738 2650 742
rect 2662 738 2666 742
rect 2678 738 2682 742
rect 2702 738 2706 742
rect 2718 738 2722 742
rect 2726 738 2730 742
rect 2742 738 2746 742
rect 2782 738 2786 742
rect 2798 738 2802 742
rect 2822 738 2826 742
rect 2862 738 2866 742
rect 2886 738 2890 742
rect 2942 738 2946 742
rect 2950 738 2954 742
rect 2974 738 2978 742
rect 2990 738 2994 742
rect 3014 738 3018 742
rect 3022 738 3026 742
rect 3062 738 3066 742
rect 3094 738 3098 742
rect 3126 738 3130 742
rect 3150 738 3154 742
rect 3190 738 3194 742
rect 3222 738 3226 742
rect 3246 738 3250 742
rect 3270 738 3274 742
rect 3286 738 3290 742
rect 3342 738 3346 742
rect 3398 738 3402 742
rect 3470 738 3474 742
rect 3478 738 3482 742
rect 3526 738 3530 742
rect 3558 738 3562 742
rect 3606 738 3610 742
rect 3622 738 3626 742
rect 3638 740 3642 744
rect 3742 738 3746 742
rect 3774 738 3778 742
rect 3790 738 3794 742
rect 3918 738 3922 742
rect 4022 738 4026 742
rect 4070 738 4074 742
rect 4102 738 4106 742
rect 4150 738 4154 742
rect 4318 738 4322 742
rect 4374 738 4378 742
rect 4398 738 4402 742
rect 4438 738 4442 742
rect 4446 738 4450 742
rect 4486 738 4490 742
rect 4510 738 4514 742
rect 4534 738 4538 742
rect 4542 738 4546 742
rect 4598 738 4602 742
rect 70 728 74 732
rect 102 728 106 732
rect 182 728 186 732
rect 230 728 234 732
rect 422 728 426 732
rect 582 728 586 732
rect 926 728 930 732
rect 1230 728 1234 732
rect 1334 728 1338 732
rect 1486 728 1490 732
rect 1542 728 1546 732
rect 1582 728 1586 732
rect 1622 728 1626 732
rect 1662 728 1666 732
rect 1678 728 1682 732
rect 1734 728 1738 732
rect 1742 728 1746 732
rect 1766 728 1770 732
rect 1830 728 1834 732
rect 1846 728 1850 732
rect 1982 728 1986 732
rect 2078 728 2082 732
rect 2158 728 2162 732
rect 2246 728 2250 732
rect 2326 728 2330 732
rect 2382 728 2386 732
rect 2414 728 2418 732
rect 2606 728 2610 732
rect 2766 728 2770 732
rect 2878 728 2882 732
rect 2998 728 3002 732
rect 3030 728 3034 732
rect 3062 728 3066 732
rect 3262 728 3266 732
rect 3406 728 3410 732
rect 3590 728 3594 732
rect 3670 728 3674 732
rect 3862 728 3866 732
rect 3926 728 3930 732
rect 4054 728 4058 732
rect 4134 728 4138 732
rect 4166 728 4170 732
rect 4374 728 4378 732
rect 4382 728 4386 732
rect 4502 728 4506 732
rect 6 718 10 722
rect 150 718 154 722
rect 374 718 378 722
rect 454 718 458 722
rect 550 718 554 722
rect 662 718 666 722
rect 742 718 746 722
rect 766 718 770 722
rect 782 718 786 722
rect 990 718 994 722
rect 1038 718 1042 722
rect 1126 718 1130 722
rect 1158 718 1162 722
rect 1262 718 1266 722
rect 1294 718 1298 722
rect 1398 718 1402 722
rect 1510 718 1514 722
rect 1654 718 1658 722
rect 1726 718 1730 722
rect 1750 718 1754 722
rect 2014 718 2018 722
rect 2062 718 2066 722
rect 2462 718 2466 722
rect 2510 718 2514 722
rect 2542 718 2546 722
rect 2686 718 2690 722
rect 2750 718 2754 722
rect 2870 718 2874 722
rect 2910 718 2914 722
rect 2966 718 2970 722
rect 2990 718 2994 722
rect 3158 718 3162 722
rect 3182 718 3186 722
rect 3366 718 3370 722
rect 3390 718 3394 722
rect 3806 718 3810 722
rect 3902 718 3906 722
rect 3966 718 3970 722
rect 4174 718 4178 722
rect 4566 718 4570 722
rect 1002 703 1006 707
rect 1009 703 1013 707
rect 2026 703 2030 707
rect 2033 703 2037 707
rect 3050 703 3054 707
rect 3057 703 3061 707
rect 4082 703 4086 707
rect 4089 703 4093 707
rect 142 688 146 692
rect 662 688 666 692
rect 958 688 962 692
rect 1222 688 1226 692
rect 1294 688 1298 692
rect 1398 688 1402 692
rect 1558 688 1562 692
rect 1622 688 1626 692
rect 1662 688 1666 692
rect 1774 688 1778 692
rect 1870 688 1874 692
rect 1934 688 1938 692
rect 1982 688 1986 692
rect 1998 688 2002 692
rect 2030 688 2034 692
rect 2118 688 2122 692
rect 2134 688 2138 692
rect 2214 688 2218 692
rect 2254 688 2258 692
rect 2374 688 2378 692
rect 2414 688 2418 692
rect 2446 688 2450 692
rect 2502 688 2506 692
rect 2598 688 2602 692
rect 2622 688 2626 692
rect 2678 688 2682 692
rect 2710 688 2714 692
rect 2742 688 2746 692
rect 2902 688 2906 692
rect 2982 688 2986 692
rect 3038 688 3042 692
rect 3094 688 3098 692
rect 3174 688 3178 692
rect 3198 688 3202 692
rect 3238 688 3242 692
rect 3270 688 3274 692
rect 3342 688 3346 692
rect 3374 688 3378 692
rect 3462 688 3466 692
rect 3502 688 3506 692
rect 3518 688 3522 692
rect 3558 688 3562 692
rect 3606 688 3610 692
rect 3614 688 3618 692
rect 3806 688 3810 692
rect 3830 688 3834 692
rect 3878 688 3882 692
rect 3998 688 4002 692
rect 4206 688 4210 692
rect 4246 688 4250 692
rect 4286 688 4290 692
rect 4414 688 4418 692
rect 4478 688 4482 692
rect 4526 688 4530 692
rect 4542 688 4546 692
rect 654 678 658 682
rect 806 678 810 682
rect 1062 678 1066 682
rect 126 668 130 672
rect 142 668 146 672
rect 206 668 210 672
rect 214 668 218 672
rect 406 668 410 672
rect 478 668 482 672
rect 582 668 586 672
rect 702 668 706 672
rect 926 668 930 672
rect 966 668 970 672
rect 1022 668 1026 672
rect 1046 668 1050 672
rect 1054 668 1058 672
rect 1070 668 1074 672
rect 1118 668 1122 672
rect 22 658 26 662
rect 70 658 74 662
rect 94 659 98 663
rect 166 658 170 662
rect 190 658 194 662
rect 198 658 202 662
rect 222 658 226 662
rect 230 658 234 662
rect 246 658 250 662
rect 270 658 274 662
rect 302 658 306 662
rect 334 658 338 662
rect 358 658 362 662
rect 390 658 394 662
rect 518 658 522 662
rect 526 658 530 662
rect 542 658 546 662
rect 590 658 594 662
rect 670 658 674 662
rect 678 658 682 662
rect 710 658 714 662
rect 758 658 762 662
rect 830 658 834 662
rect 894 659 898 663
rect 1174 668 1178 672
rect 1198 678 1202 682
rect 1214 668 1218 672
rect 1334 678 1338 682
rect 1342 678 1346 682
rect 1358 678 1362 682
rect 1374 678 1378 682
rect 1430 678 1434 682
rect 1550 678 1554 682
rect 1646 678 1650 682
rect 1678 678 1682 682
rect 1974 678 1978 682
rect 2006 678 2010 682
rect 2126 678 2130 682
rect 2158 678 2162 682
rect 2302 678 2306 682
rect 2342 678 2346 682
rect 2398 678 2402 682
rect 2518 678 2522 682
rect 2654 678 2658 682
rect 2686 678 2690 682
rect 2718 678 2722 682
rect 2750 678 2754 682
rect 2974 678 2978 682
rect 3030 678 3034 682
rect 3142 678 3146 682
rect 3654 678 3658 682
rect 3798 678 3802 682
rect 3886 678 3890 682
rect 3950 678 3954 682
rect 4198 678 4202 682
rect 4254 678 4258 682
rect 4302 678 4306 682
rect 4318 678 4322 682
rect 4366 678 4370 682
rect 4574 678 4578 682
rect 1262 668 1266 672
rect 1310 668 1314 672
rect 1366 668 1370 672
rect 1438 668 1442 672
rect 1486 668 1490 672
rect 1494 668 1498 672
rect 1558 668 1562 672
rect 1614 668 1618 672
rect 1630 668 1634 672
rect 1670 668 1674 672
rect 1726 668 1730 672
rect 1734 668 1738 672
rect 1798 668 1802 672
rect 1822 668 1826 672
rect 1854 668 1858 672
rect 1894 668 1898 672
rect 2086 668 2090 672
rect 918 658 922 662
rect 1038 658 1042 662
rect 1126 658 1130 662
rect 1158 658 1162 662
rect 1198 658 1202 662
rect 2142 668 2146 672
rect 2182 668 2186 672
rect 2198 668 2202 672
rect 2238 668 2242 672
rect 2246 668 2250 672
rect 2278 668 2282 672
rect 2430 668 2434 672
rect 2438 668 2442 672
rect 2510 668 2514 672
rect 2582 668 2586 672
rect 2614 668 2618 672
rect 2654 668 2658 672
rect 2702 668 2706 672
rect 2734 668 2738 672
rect 2766 668 2770 672
rect 2782 668 2786 672
rect 2806 668 2810 672
rect 2846 668 2850 672
rect 2878 668 2882 672
rect 2910 668 2914 672
rect 2926 668 2930 672
rect 2942 668 2946 672
rect 2990 668 2994 672
rect 3006 668 3010 672
rect 3054 668 3058 672
rect 3078 668 3082 672
rect 3102 668 3106 672
rect 3166 668 3170 672
rect 3190 668 3194 672
rect 3214 668 3218 672
rect 3246 668 3250 672
rect 3278 668 3282 672
rect 3294 668 3298 672
rect 3326 668 3330 672
rect 3350 668 3354 672
rect 3358 668 3362 672
rect 3382 668 3386 672
rect 3414 668 3418 672
rect 3430 668 3434 672
rect 3438 668 3442 672
rect 3486 668 3490 672
rect 3510 668 3514 672
rect 3542 668 3546 672
rect 3590 668 3594 672
rect 3638 668 3642 672
rect 3662 668 3666 672
rect 3694 668 3698 672
rect 3710 668 3714 672
rect 3838 668 3842 672
rect 3862 668 3866 672
rect 3894 668 3898 672
rect 3950 668 3954 672
rect 3982 668 3986 672
rect 4014 668 4018 672
rect 4030 668 4034 672
rect 4070 668 4074 672
rect 4094 668 4098 672
rect 4110 668 4114 672
rect 4118 668 4122 672
rect 4150 668 4154 672
rect 4158 668 4162 672
rect 4190 668 4194 672
rect 4214 668 4218 672
rect 4238 668 4242 672
rect 4262 668 4266 672
rect 4294 668 4298 672
rect 4358 668 4362 672
rect 4406 668 4410 672
rect 1238 658 1242 662
rect 1318 658 1322 662
rect 1334 658 1338 662
rect 1406 658 1410 662
rect 1414 658 1418 662
rect 1422 658 1426 662
rect 1430 658 1434 662
rect 1502 658 1506 662
rect 1566 658 1570 662
rect 1606 658 1610 662
rect 1638 658 1642 662
rect 1694 658 1698 662
rect 1718 658 1722 662
rect 1742 658 1746 662
rect 1750 658 1754 662
rect 1782 658 1786 662
rect 1806 658 1810 662
rect 1846 658 1850 662
rect 1878 658 1882 662
rect 1950 658 1954 662
rect 1990 658 1994 662
rect 2014 658 2018 662
rect 2078 658 2082 662
rect 2094 658 2098 662
rect 2102 658 2106 662
rect 2150 658 2154 662
rect 2174 658 2178 662
rect 2214 658 2218 662
rect 2230 658 2234 662
rect 2270 658 2274 662
rect 2318 658 2322 662
rect 2342 658 2346 662
rect 2358 658 2362 662
rect 2382 658 2386 662
rect 2398 658 2402 662
rect 2486 658 2490 662
rect 2558 658 2562 662
rect 2574 658 2578 662
rect 2606 658 2610 662
rect 2630 658 2634 662
rect 2662 658 2666 662
rect 2694 658 2698 662
rect 2726 658 2730 662
rect 2774 658 2778 662
rect 2830 658 2834 662
rect 2870 658 2874 662
rect 2886 658 2890 662
rect 2918 658 2922 662
rect 2950 658 2954 662
rect 2998 658 3002 662
rect 3014 658 3018 662
rect 3110 658 3114 662
rect 3134 658 3138 662
rect 3158 658 3162 662
rect 3222 658 3226 662
rect 3254 658 3258 662
rect 3286 658 3290 662
rect 3422 658 3426 662
rect 3478 658 3482 662
rect 3630 658 3634 662
rect 3702 658 3706 662
rect 3726 658 3730 662
rect 3750 658 3754 662
rect 3758 658 3762 662
rect 3766 658 3770 662
rect 3798 658 3802 662
rect 3814 658 3818 662
rect 3870 658 3874 662
rect 3934 658 3938 662
rect 3950 658 3954 662
rect 4006 658 4010 662
rect 4038 658 4042 662
rect 4062 658 4066 662
rect 4126 658 4130 662
rect 4150 658 4154 662
rect 4166 658 4170 662
rect 4182 658 4186 662
rect 4222 658 4226 662
rect 4230 658 4234 662
rect 4270 658 4274 662
rect 4286 658 4290 662
rect 4318 658 4322 662
rect 4342 658 4346 662
rect 4374 658 4378 662
rect 4398 658 4402 662
rect 4430 658 4434 662
rect 4446 668 4450 672
rect 4486 658 4490 662
rect 4534 668 4538 672
rect 4558 668 4562 672
rect 4510 658 4514 662
rect 4550 658 4554 662
rect 142 648 146 652
rect 174 648 178 652
rect 182 648 186 652
rect 238 648 242 652
rect 318 648 322 652
rect 366 648 370 652
rect 398 648 402 652
rect 550 648 554 652
rect 726 648 730 652
rect 6 638 10 642
rect 158 638 162 642
rect 286 638 290 642
rect 350 638 354 642
rect 382 638 386 642
rect 534 638 538 642
rect 742 638 746 642
rect 750 638 754 642
rect 1382 648 1386 652
rect 1518 648 1522 652
rect 1758 648 1762 652
rect 1790 648 1794 652
rect 1830 648 1834 652
rect 1894 648 1898 652
rect 1910 648 1914 652
rect 1934 648 1938 652
rect 1942 648 1946 652
rect 2062 648 2066 652
rect 2118 648 2122 652
rect 2182 648 2186 652
rect 2294 648 2298 652
rect 2454 648 2458 652
rect 2494 648 2498 652
rect 2542 648 2546 652
rect 2758 648 2762 652
rect 2790 648 2794 652
rect 2814 648 2818 652
rect 2830 648 2834 652
rect 2902 648 2906 652
rect 2934 648 2938 652
rect 2966 648 2970 652
rect 3030 648 3034 652
rect 3038 648 3042 652
rect 3094 648 3098 652
rect 3126 648 3130 652
rect 3182 648 3186 652
rect 3206 648 3210 652
rect 3238 648 3242 652
rect 3270 648 3274 652
rect 3310 648 3314 652
rect 3334 648 3338 652
rect 3374 648 3378 652
rect 3398 648 3402 652
rect 3454 648 3458 652
rect 3494 648 3498 652
rect 3510 648 3514 652
rect 3550 648 3554 652
rect 3606 648 3610 652
rect 3614 648 3618 652
rect 3678 648 3682 652
rect 3822 648 3826 652
rect 3846 648 3850 652
rect 3974 648 3978 652
rect 3998 648 4002 652
rect 4046 648 4050 652
rect 4110 648 4114 652
rect 4182 648 4186 652
rect 4350 648 4354 652
rect 4414 648 4418 652
rect 4446 648 4450 652
rect 4462 648 4466 652
rect 4494 648 4498 652
rect 4526 648 4530 652
rect 1718 638 1722 642
rect 1774 638 1778 642
rect 1870 638 1874 642
rect 1918 638 1922 642
rect 1950 638 1954 642
rect 1958 638 1962 642
rect 3654 638 3658 642
rect 3902 638 3906 642
rect 3926 638 3930 642
rect 4334 638 4338 642
rect 4478 638 4482 642
rect 358 628 362 632
rect 646 628 650 632
rect 30 618 34 622
rect 390 618 394 622
rect 462 618 466 622
rect 990 618 994 622
rect 1094 618 1098 622
rect 1350 618 1354 622
rect 1502 618 1506 622
rect 1654 618 1658 622
rect 1982 618 1986 622
rect 2174 618 2178 622
rect 2470 618 2474 622
rect 2526 618 2530 622
rect 2574 618 2578 622
rect 2798 618 2802 622
rect 2854 618 2858 622
rect 2950 618 2954 622
rect 3742 618 3746 622
rect 3854 618 3858 622
rect 4014 618 4018 622
rect 4062 618 4066 622
rect 4126 618 4130 622
rect 4326 618 4330 622
rect 4582 618 4586 622
rect 498 603 502 607
rect 505 603 509 607
rect 1522 603 1526 607
rect 1529 603 1533 607
rect 2546 603 2550 607
rect 2553 603 2557 607
rect 3570 603 3574 607
rect 3577 603 3581 607
rect 254 588 258 592
rect 390 588 394 592
rect 526 588 530 592
rect 654 588 658 592
rect 1134 588 1138 592
rect 1150 588 1154 592
rect 1326 588 1330 592
rect 1390 588 1394 592
rect 1550 588 1554 592
rect 1630 588 1634 592
rect 1862 588 1866 592
rect 1886 588 1890 592
rect 1974 588 1978 592
rect 2054 588 2058 592
rect 2110 588 2114 592
rect 2126 588 2130 592
rect 2254 588 2258 592
rect 2294 588 2298 592
rect 2438 588 2442 592
rect 2614 588 2618 592
rect 2670 588 2674 592
rect 2710 588 2714 592
rect 2846 588 2850 592
rect 2870 588 2874 592
rect 2942 588 2946 592
rect 2990 588 2994 592
rect 3142 588 3146 592
rect 3222 588 3226 592
rect 3278 588 3282 592
rect 3286 588 3290 592
rect 3318 588 3322 592
rect 3398 588 3402 592
rect 3454 588 3458 592
rect 3478 588 3482 592
rect 3542 588 3546 592
rect 3686 588 3690 592
rect 4014 588 4018 592
rect 4246 588 4250 592
rect 4302 588 4306 592
rect 4350 588 4354 592
rect 4478 588 4482 592
rect 4542 588 4546 592
rect 4574 588 4578 592
rect 1470 578 1474 582
rect 3934 578 3938 582
rect 30 568 34 572
rect 70 568 74 572
rect 254 568 258 572
rect 262 568 266 572
rect 798 568 802 572
rect 854 568 858 572
rect 862 568 866 572
rect 902 568 906 572
rect 998 568 1002 572
rect 1446 568 1450 572
rect 1478 568 1482 572
rect 1486 568 1490 572
rect 2134 568 2138 572
rect 2342 568 2346 572
rect 2422 568 2426 572
rect 2982 568 2986 572
rect 3694 568 3698 572
rect 4326 568 4330 572
rect 4390 568 4394 572
rect 278 558 282 562
rect 662 558 666 562
rect 742 558 746 562
rect 22 548 26 552
rect 830 558 834 562
rect 870 558 874 562
rect 902 558 906 562
rect 1158 558 1162 562
rect 1382 558 1386 562
rect 1494 558 1498 562
rect 1502 558 1506 562
rect 118 547 122 551
rect 174 547 178 551
rect 206 548 210 552
rect 254 548 258 552
rect 326 547 330 551
rect 358 548 362 552
rect 422 547 426 551
rect 454 548 458 552
rect 590 547 594 551
rect 694 548 698 552
rect 718 548 722 552
rect 734 548 738 552
rect 750 548 754 552
rect 774 548 778 552
rect 782 548 786 552
rect 798 548 802 552
rect 814 548 818 552
rect 862 548 866 552
rect 894 548 898 552
rect 942 548 946 552
rect 966 548 970 552
rect 1014 548 1018 552
rect 6 538 10 542
rect 294 538 298 542
rect 310 538 314 542
rect 510 538 514 542
rect 574 538 578 542
rect 678 540 682 544
rect 686 538 690 542
rect 1070 547 1074 551
rect 1102 548 1106 552
rect 1262 547 1266 551
rect 1350 548 1354 552
rect 1366 548 1370 552
rect 1390 548 1394 552
rect 1486 548 1490 552
rect 1582 558 1586 562
rect 1662 558 1666 562
rect 1598 548 1602 552
rect 1702 558 1706 562
rect 1686 548 1690 552
rect 1726 548 1730 552
rect 1734 548 1738 552
rect 1758 548 1762 552
rect 1790 558 1794 562
rect 1822 558 1826 562
rect 1878 558 1882 562
rect 1910 558 1914 562
rect 1790 548 1794 552
rect 1814 548 1818 552
rect 1830 548 1834 552
rect 1862 548 1866 552
rect 1902 548 1906 552
rect 1990 558 1994 562
rect 1998 558 2002 562
rect 2078 558 2082 562
rect 2150 558 2154 562
rect 2238 558 2242 562
rect 2278 558 2282 562
rect 2326 558 2330 562
rect 2366 558 2370 562
rect 2454 558 2458 562
rect 2494 558 2498 562
rect 2510 558 2514 562
rect 2630 558 2634 562
rect 2654 558 2658 562
rect 2662 558 2666 562
rect 2742 558 2746 562
rect 2758 558 2762 562
rect 2790 558 2794 562
rect 2822 558 2826 562
rect 2910 558 2914 562
rect 2918 558 2922 562
rect 3006 558 3010 562
rect 3038 558 3042 562
rect 3094 558 3098 562
rect 3126 558 3130 562
rect 3166 558 3170 562
rect 3182 558 3186 562
rect 3262 558 3266 562
rect 3302 558 3306 562
rect 1974 548 1978 552
rect 1998 548 2002 552
rect 2014 548 2018 552
rect 2062 548 2066 552
rect 2118 548 2122 552
rect 2134 548 2138 552
rect 2158 548 2162 552
rect 2190 548 2194 552
rect 2198 548 2202 552
rect 2206 548 2210 552
rect 2262 548 2266 552
rect 2270 548 2274 552
rect 2318 548 2322 552
rect 2358 548 2362 552
rect 2366 548 2370 552
rect 2382 548 2386 552
rect 2390 548 2394 552
rect 2406 548 2410 552
rect 2438 548 2442 552
rect 2470 548 2474 552
rect 2486 548 2490 552
rect 2510 548 2514 552
rect 2574 548 2578 552
rect 2598 548 2602 552
rect 2614 548 2618 552
rect 2654 548 2658 552
rect 2686 548 2690 552
rect 2702 548 2706 552
rect 2734 548 2738 552
rect 2774 548 2778 552
rect 2806 548 2810 552
rect 2830 548 2834 552
rect 2870 548 2874 552
rect 2966 548 2970 552
rect 2982 548 2986 552
rect 3038 548 3042 552
rect 3110 548 3114 552
rect 3166 548 3170 552
rect 3182 548 3186 552
rect 3198 548 3202 552
rect 3206 548 3210 552
rect 3230 548 3234 552
rect 3262 548 3266 552
rect 3318 548 3322 552
rect 3358 548 3362 552
rect 3366 548 3370 552
rect 3382 558 3386 562
rect 3430 558 3434 562
rect 3382 548 3386 552
rect 3406 548 3410 552
rect 3486 558 3490 562
rect 3518 558 3522 562
rect 3454 548 3458 552
rect 3510 548 3514 552
rect 3542 548 3546 552
rect 3582 558 3586 562
rect 3622 558 3626 562
rect 3662 558 3666 562
rect 3670 558 3674 562
rect 3710 558 3714 562
rect 3758 558 3762 562
rect 3838 558 3842 562
rect 3854 558 3858 562
rect 3862 558 3866 562
rect 4062 558 4066 562
rect 4134 558 4138 562
rect 4230 558 4234 562
rect 4406 558 4410 562
rect 4438 558 4442 562
rect 4558 558 4562 562
rect 3646 548 3650 552
rect 3702 548 3706 552
rect 3718 548 3722 552
rect 3766 548 3770 552
rect 3782 548 3786 552
rect 3798 548 3802 552
rect 3806 548 3810 552
rect 3862 548 3866 552
rect 3878 548 3882 552
rect 3910 548 3914 552
rect 3934 548 3938 552
rect 3950 548 3954 552
rect 3990 548 3994 552
rect 3998 548 4002 552
rect 4006 548 4010 552
rect 4038 548 4042 552
rect 4054 548 4058 552
rect 4078 548 4082 552
rect 4110 548 4114 552
rect 4150 548 4154 552
rect 806 538 810 542
rect 918 538 922 542
rect 1142 538 1146 542
rect 1166 538 1170 542
rect 1246 538 1250 542
rect 1414 538 1418 542
rect 1462 538 1466 542
rect 1518 538 1522 542
rect 1558 538 1562 542
rect 1622 538 1626 542
rect 1646 538 1650 542
rect 1718 538 1722 542
rect 1798 538 1802 542
rect 1854 538 1858 542
rect 1918 538 1922 542
rect 1966 538 1970 542
rect 2022 538 2026 542
rect 2094 538 2098 542
rect 2110 538 2114 542
rect 2214 538 2218 542
rect 2262 538 2266 542
rect 2310 538 2314 542
rect 2350 538 2354 542
rect 2358 538 2362 542
rect 2398 538 2402 542
rect 2494 538 2498 542
rect 2534 538 2538 542
rect 2574 538 2578 542
rect 2606 538 2610 542
rect 2638 538 2642 542
rect 2678 538 2682 542
rect 2726 538 2730 542
rect 2766 538 2770 542
rect 2798 538 2802 542
rect 2854 538 2858 542
rect 2862 538 2866 542
rect 2894 538 2898 542
rect 2934 538 2938 542
rect 2958 538 2962 542
rect 3022 538 3026 542
rect 3030 538 3034 542
rect 3070 538 3074 542
rect 3102 538 3106 542
rect 3118 538 3122 542
rect 3190 538 3194 542
rect 3246 538 3250 542
rect 3350 538 3354 542
rect 3406 538 3410 542
rect 3414 538 3418 542
rect 3470 538 3474 542
rect 3494 538 3498 542
rect 3598 538 3602 542
rect 3606 538 3610 542
rect 3654 538 3658 542
rect 3678 538 3682 542
rect 3734 538 3738 542
rect 3790 538 3794 542
rect 3814 538 3818 542
rect 3830 538 3834 542
rect 3854 538 3858 542
rect 3918 538 3922 542
rect 3942 538 3946 542
rect 3974 538 3978 542
rect 4046 538 4050 542
rect 4070 538 4074 542
rect 4142 538 4146 542
rect 4166 538 4170 542
rect 4182 538 4186 542
rect 4198 548 4202 552
rect 4246 548 4250 552
rect 4262 548 4266 552
rect 4294 548 4298 552
rect 4318 548 4322 552
rect 4326 548 4330 552
rect 4374 548 4378 552
rect 4382 548 4386 552
rect 4430 548 4434 552
rect 4454 548 4458 552
rect 4462 548 4466 552
rect 4502 548 4506 552
rect 4510 548 4514 552
rect 4526 548 4530 552
rect 4574 548 4578 552
rect 4198 538 4202 542
rect 4206 538 4210 542
rect 4254 538 4258 542
rect 4286 538 4290 542
rect 4318 538 4322 542
rect 4366 538 4370 542
rect 4374 538 4378 542
rect 4414 538 4418 542
rect 4462 538 4466 542
rect 4470 538 4474 542
rect 4494 538 4498 542
rect 4510 538 4514 542
rect 4582 538 4586 542
rect 710 528 714 532
rect 1334 528 1338 532
rect 1406 528 1410 532
rect 1542 528 1546 532
rect 1566 528 1570 532
rect 1638 528 1642 532
rect 1846 528 1850 532
rect 1942 528 1946 532
rect 2046 528 2050 532
rect 2054 528 2058 532
rect 2078 528 2082 532
rect 2230 528 2234 532
rect 2286 528 2290 532
rect 2294 528 2298 532
rect 2382 528 2386 532
rect 2542 528 2546 532
rect 2582 528 2586 532
rect 2686 528 2690 532
rect 2790 528 2794 532
rect 2942 528 2946 532
rect 3270 528 3274 532
rect 3294 528 3298 532
rect 3342 528 3346 532
rect 3518 528 3522 532
rect 3830 528 3834 532
rect 3894 528 3898 532
rect 3918 528 3922 532
rect 3982 528 3986 532
rect 4022 528 4026 532
rect 4030 528 4034 532
rect 4110 528 4114 532
rect 4126 528 4130 532
rect 4166 528 4170 532
rect 4222 528 4226 532
rect 4278 528 4282 532
rect 4342 528 4346 532
rect 4534 528 4538 532
rect 4550 528 4554 532
rect 286 518 290 522
rect 486 518 490 522
rect 846 518 850 522
rect 1038 518 1042 522
rect 1222 518 1226 522
rect 1342 518 1346 522
rect 1382 518 1386 522
rect 1510 518 1514 522
rect 1614 518 1618 522
rect 1670 518 1674 522
rect 1710 518 1714 522
rect 1750 518 1754 522
rect 1838 518 1842 522
rect 2174 518 2178 522
rect 2222 518 2226 522
rect 2510 518 2514 522
rect 2822 518 2826 522
rect 2926 518 2930 522
rect 3630 518 3634 522
rect 3726 518 3730 522
rect 3822 518 3826 522
rect 3950 518 3954 522
rect 4174 518 4178 522
rect 4214 518 4218 522
rect 4270 518 4274 522
rect 4438 518 4442 522
rect 4542 518 4546 522
rect 1002 503 1006 507
rect 1009 503 1013 507
rect 2026 503 2030 507
rect 2033 503 2037 507
rect 3050 503 3054 507
rect 3057 503 3061 507
rect 4082 503 4086 507
rect 4089 503 4093 507
rect 126 488 130 492
rect 542 488 546 492
rect 718 488 722 492
rect 782 488 786 492
rect 1174 488 1178 492
rect 1270 488 1274 492
rect 1430 488 1434 492
rect 1502 488 1506 492
rect 1622 488 1626 492
rect 1654 488 1658 492
rect 1790 488 1794 492
rect 1854 488 1858 492
rect 1910 488 1914 492
rect 1966 488 1970 492
rect 2062 488 2066 492
rect 2078 488 2082 492
rect 2110 488 2114 492
rect 2206 488 2210 492
rect 2230 488 2234 492
rect 2286 488 2290 492
rect 2302 488 2306 492
rect 2366 488 2370 492
rect 2470 488 2474 492
rect 2518 488 2522 492
rect 2710 488 2714 492
rect 2790 488 2794 492
rect 2806 488 2810 492
rect 2838 488 2842 492
rect 2862 488 2866 492
rect 2902 488 2906 492
rect 2990 488 2994 492
rect 3014 488 3018 492
rect 3078 488 3082 492
rect 3150 488 3154 492
rect 3182 488 3186 492
rect 3222 488 3226 492
rect 3246 488 3250 492
rect 3278 488 3282 492
rect 3382 488 3386 492
rect 3398 488 3402 492
rect 3582 488 3586 492
rect 3806 488 3810 492
rect 3902 488 3906 492
rect 4006 488 4010 492
rect 4062 488 4066 492
rect 4310 488 4314 492
rect 4358 488 4362 492
rect 4374 488 4378 492
rect 4390 488 4394 492
rect 4398 488 4402 492
rect 4430 488 4434 492
rect 4446 488 4450 492
rect 4550 488 4554 492
rect 478 478 482 482
rect 622 478 626 482
rect 734 478 738 482
rect 1526 478 1530 482
rect 1718 478 1722 482
rect 1782 478 1786 482
rect 1846 478 1850 482
rect 1918 478 1922 482
rect 1998 478 2002 482
rect 2094 478 2098 482
rect 2118 478 2122 482
rect 2182 478 2186 482
rect 2294 478 2298 482
rect 2374 478 2378 482
rect 2398 478 2402 482
rect 2406 478 2410 482
rect 2478 478 2482 482
rect 2486 478 2490 482
rect 2670 478 2674 482
rect 2702 478 2706 482
rect 2782 478 2786 482
rect 2894 478 2898 482
rect 3038 478 3042 482
rect 3062 478 3066 482
rect 278 468 282 472
rect 390 468 394 472
rect 534 468 538 472
rect 558 468 562 472
rect 638 468 642 472
rect 670 468 674 472
rect 734 468 738 472
rect 750 468 754 472
rect 902 468 906 472
rect 1030 468 1034 472
rect 1094 468 1098 472
rect 1222 468 1226 472
rect 1278 468 1282 472
rect 1326 468 1330 472
rect 1334 468 1338 472
rect 1382 468 1386 472
rect 1390 468 1394 472
rect 1422 468 1426 472
rect 1438 468 1442 472
rect 1470 468 1474 472
rect 1478 468 1482 472
rect 1550 468 1554 472
rect 1598 468 1602 472
rect 1614 468 1618 472
rect 1630 468 1634 472
rect 1654 468 1658 472
rect 1670 468 1674 472
rect 1686 468 1690 472
rect 1822 468 1826 472
rect 1878 468 1882 472
rect 1886 468 1890 472
rect 1942 468 1946 472
rect 1990 468 1994 472
rect 2022 468 2026 472
rect 2046 468 2050 472
rect 2070 468 2074 472
rect 2094 468 2098 472
rect 2126 468 2130 472
rect 2158 468 2162 472
rect 2174 468 2178 472
rect 2214 468 2218 472
rect 2222 468 2226 472
rect 2254 468 2258 472
rect 2262 468 2266 472
rect 2398 468 2402 472
rect 2422 468 2426 472
rect 2438 468 2442 472
rect 2454 468 2458 472
rect 2502 468 2506 472
rect 2542 468 2546 472
rect 2590 468 2594 472
rect 2598 468 2602 472
rect 2630 468 2634 472
rect 2670 468 2674 472
rect 2686 468 2690 472
rect 2718 468 2722 472
rect 2758 468 2762 472
rect 2774 468 2778 472
rect 2822 468 2826 472
rect 2846 468 2850 472
rect 2886 468 2890 472
rect 2910 468 2914 472
rect 2950 468 2954 472
rect 2982 468 2986 472
rect 3006 468 3010 472
rect 3030 468 3034 472
rect 3238 478 3242 482
rect 3294 478 3298 482
rect 3622 478 3626 482
rect 3742 478 3746 482
rect 3814 478 3818 482
rect 3854 478 3858 482
rect 3870 478 3874 482
rect 3878 478 3882 482
rect 3982 478 3986 482
rect 4054 478 4058 482
rect 4102 478 4106 482
rect 4118 478 4122 482
rect 3094 468 3098 472
rect 3110 468 3114 472
rect 3126 468 3130 472
rect 3174 468 3178 472
rect 3206 468 3210 472
rect 3230 468 3234 472
rect 3254 468 3258 472
rect 3286 468 3290 472
rect 3318 468 3322 472
rect 3390 468 3394 472
rect 3422 468 3426 472
rect 3438 468 3442 472
rect 3462 468 3466 472
rect 3478 468 3482 472
rect 3542 468 3546 472
rect 3558 468 3562 472
rect 3678 468 3682 472
rect 3838 468 3842 472
rect 3886 468 3890 472
rect 3910 468 3914 472
rect 3918 468 3922 472
rect 4014 468 4018 472
rect 4046 468 4050 472
rect 4070 468 4074 472
rect 4150 468 4154 472
rect 4190 468 4194 472
rect 4246 468 4250 472
rect 4254 468 4258 472
rect 4270 468 4274 472
rect 4342 478 4346 482
rect 4382 478 4386 482
rect 4462 478 4466 482
rect 4502 478 4506 482
rect 4510 478 4514 482
rect 4302 468 4306 472
rect 4350 468 4354 472
rect 4406 468 4410 472
rect 4414 468 4418 472
rect 4518 468 4522 472
rect 4534 468 4538 472
rect 4574 468 4578 472
rect 22 458 26 462
rect 54 459 58 463
rect 86 458 90 462
rect 158 458 162 462
rect 190 459 194 463
rect 238 458 242 462
rect 270 458 274 462
rect 294 458 298 462
rect 318 458 322 462
rect 342 458 346 462
rect 366 458 370 462
rect 406 459 410 463
rect 518 458 522 462
rect 566 458 570 462
rect 606 458 610 462
rect 646 458 650 462
rect 662 458 666 462
rect 694 458 698 462
rect 766 458 770 462
rect 814 458 818 462
rect 846 459 850 463
rect 878 458 882 462
rect 894 458 898 462
rect 926 458 930 462
rect 958 458 962 462
rect 1014 459 1018 463
rect 1110 459 1114 463
rect 1206 459 1210 463
rect 1398 458 1402 462
rect 222 448 226 452
rect 286 448 290 452
rect 374 448 378 452
rect 614 448 618 452
rect 622 448 626 452
rect 702 448 706 452
rect 710 448 714 452
rect 774 448 778 452
rect 934 448 938 452
rect 982 448 986 452
rect 1414 448 1418 452
rect 1446 458 1450 462
rect 1462 458 1466 462
rect 1486 458 1490 462
rect 1510 458 1514 462
rect 1518 458 1522 462
rect 1526 458 1530 462
rect 1606 458 1610 462
rect 1646 458 1650 462
rect 1678 458 1682 462
rect 1694 458 1698 462
rect 1742 458 1746 462
rect 1766 458 1770 462
rect 1774 458 1778 462
rect 1814 458 1818 462
rect 1822 458 1826 462
rect 1870 458 1874 462
rect 1894 458 1898 462
rect 1934 458 1938 462
rect 1950 458 1954 462
rect 2014 458 2018 462
rect 2126 458 2130 462
rect 2230 458 2234 462
rect 2254 458 2258 462
rect 2270 458 2274 462
rect 2318 458 2322 462
rect 2342 458 2346 462
rect 2358 458 2362 462
rect 2382 458 2386 462
rect 2414 458 2418 462
rect 2462 458 2466 462
rect 2494 458 2498 462
rect 2510 458 2514 462
rect 2534 458 2538 462
rect 2582 458 2586 462
rect 2606 458 2610 462
rect 2638 458 2642 462
rect 2654 458 2658 462
rect 2662 458 2666 462
rect 2694 458 2698 462
rect 2718 458 2722 462
rect 2766 458 2770 462
rect 2806 458 2810 462
rect 2830 458 2834 462
rect 2862 458 2866 462
rect 2878 458 2882 462
rect 2918 458 2922 462
rect 2934 458 2938 462
rect 2942 458 2946 462
rect 2974 458 2978 462
rect 3070 458 3074 462
rect 3102 458 3106 462
rect 3134 458 3138 462
rect 3198 458 3202 462
rect 3262 458 3266 462
rect 3310 458 3314 462
rect 3326 458 3330 462
rect 3334 458 3338 462
rect 3350 458 3354 462
rect 3358 458 3362 462
rect 3430 458 3434 462
rect 3454 458 3458 462
rect 3470 458 3474 462
rect 3494 458 3498 462
rect 3502 458 3506 462
rect 3526 458 3530 462
rect 3566 458 3570 462
rect 3598 458 3602 462
rect 3622 458 3626 462
rect 3630 458 3634 462
rect 3662 458 3666 462
rect 3670 458 3674 462
rect 3718 458 3722 462
rect 3750 458 3754 462
rect 3758 458 3762 462
rect 3782 458 3786 462
rect 3798 458 3802 462
rect 3830 458 3834 462
rect 3854 458 3858 462
rect 3950 458 3954 462
rect 3998 458 4002 462
rect 4038 458 4042 462
rect 4118 458 4122 462
rect 4142 458 4146 462
rect 4174 458 4178 462
rect 4198 458 4202 462
rect 4214 458 4218 462
rect 4238 458 4242 462
rect 4278 458 4282 462
rect 4294 458 4298 462
rect 4326 458 4330 462
rect 4366 458 4370 462
rect 4478 458 4482 462
rect 4486 458 4490 462
rect 1446 448 1450 452
rect 1502 448 1506 452
rect 1710 448 1714 452
rect 1798 448 1802 452
rect 1814 448 1818 452
rect 1974 448 1978 452
rect 1998 448 2002 452
rect 2070 448 2074 452
rect 2158 448 2162 452
rect 2286 448 2290 452
rect 2326 448 2330 452
rect 2438 448 2442 452
rect 2518 448 2522 452
rect 2566 448 2570 452
rect 2622 448 2626 452
rect 2742 448 2746 452
rect 2750 448 2754 452
rect 2806 448 2810 452
rect 2830 448 2834 452
rect 2926 448 2930 452
rect 2958 448 2962 452
rect 2974 448 2978 452
rect 2990 448 2994 452
rect 3014 448 3018 452
rect 3118 448 3122 452
rect 3158 448 3162 452
rect 3182 448 3186 452
rect 3214 448 3218 452
rect 3270 448 3274 452
rect 3294 448 3298 452
rect 3374 448 3378 452
rect 3398 448 3402 452
rect 3486 448 3490 452
rect 3694 448 3698 452
rect 3822 448 3826 452
rect 3894 448 3898 452
rect 3934 448 3938 452
rect 3942 448 3946 452
rect 3974 448 3978 452
rect 3990 448 3994 452
rect 4022 448 4026 452
rect 4126 448 4130 452
rect 4158 448 4162 452
rect 4198 448 4202 452
rect 4214 448 4218 452
rect 4254 448 4258 452
rect 4318 448 4322 452
rect 4390 448 4394 452
rect 4430 448 4434 452
rect 4438 448 4442 452
rect 4518 448 4522 452
rect 4542 448 4546 452
rect 4558 448 4562 452
rect 6 438 10 442
rect 118 438 122 442
rect 238 438 242 442
rect 254 438 258 442
rect 302 438 306 442
rect 358 438 362 442
rect 478 438 482 442
rect 582 438 586 442
rect 598 438 602 442
rect 686 438 690 442
rect 694 438 698 442
rect 894 438 898 442
rect 918 438 922 442
rect 926 438 930 442
rect 950 438 954 442
rect 1078 438 1082 442
rect 1158 438 1162 442
rect 2726 438 2730 442
rect 3838 438 3842 442
rect 3958 438 3962 442
rect 230 428 234 432
rect 270 428 274 432
rect 294 428 298 432
rect 4326 428 4330 432
rect 326 418 330 422
rect 366 418 370 422
rect 590 418 594 422
rect 926 418 930 422
rect 1302 418 1306 422
rect 1358 418 1362 422
rect 1398 418 1402 422
rect 1694 418 1698 422
rect 1726 418 1730 422
rect 1758 418 1762 422
rect 2446 418 2450 422
rect 2606 418 2610 422
rect 2654 418 2658 422
rect 3518 418 3522 422
rect 3718 418 3722 422
rect 3774 418 3778 422
rect 3926 418 3930 422
rect 3950 418 3954 422
rect 4038 418 4042 422
rect 4174 418 4178 422
rect 4238 418 4242 422
rect 498 403 502 407
rect 505 403 509 407
rect 1522 403 1526 407
rect 1529 403 1533 407
rect 2546 403 2550 407
rect 2553 403 2557 407
rect 3570 403 3574 407
rect 3577 403 3581 407
rect 286 388 290 392
rect 350 388 354 392
rect 606 388 610 392
rect 726 388 730 392
rect 806 388 810 392
rect 1166 388 1170 392
rect 1486 388 1490 392
rect 1534 388 1538 392
rect 1790 388 1794 392
rect 1822 388 1826 392
rect 1846 388 1850 392
rect 1870 388 1874 392
rect 2030 388 2034 392
rect 2078 388 2082 392
rect 2094 388 2098 392
rect 2134 388 2138 392
rect 2158 388 2162 392
rect 2190 388 2194 392
rect 2350 388 2354 392
rect 2422 388 2426 392
rect 2622 388 2626 392
rect 2646 388 2650 392
rect 2766 388 2770 392
rect 2806 388 2810 392
rect 2886 388 2890 392
rect 2942 388 2946 392
rect 2990 388 2994 392
rect 3030 388 3034 392
rect 3078 388 3082 392
rect 3110 388 3114 392
rect 3198 388 3202 392
rect 3262 388 3266 392
rect 3302 388 3306 392
rect 3366 388 3370 392
rect 3414 388 3418 392
rect 3454 388 3458 392
rect 3606 388 3610 392
rect 3670 388 3674 392
rect 3830 388 3834 392
rect 3934 388 3938 392
rect 4038 388 4042 392
rect 4118 388 4122 392
rect 4206 388 4210 392
rect 4262 388 4266 392
rect 4342 388 4346 392
rect 4470 388 4474 392
rect 4558 388 4562 392
rect 78 378 82 382
rect 1662 378 1666 382
rect 310 368 314 372
rect 326 368 330 372
rect 358 368 362 372
rect 582 368 586 372
rect 1774 368 1778 372
rect 2166 368 2170 372
rect 2262 368 2266 372
rect 3166 368 3170 372
rect 4126 368 4130 372
rect 4142 368 4146 372
rect 22 358 26 362
rect 118 358 122 362
rect 126 358 130 362
rect 222 358 226 362
rect 278 358 282 362
rect 302 358 306 362
rect 342 358 346 362
rect 374 358 378 362
rect 470 358 474 362
rect 518 358 522 362
rect 598 358 602 362
rect 742 358 746 362
rect 750 358 754 362
rect 790 358 794 362
rect 1478 358 1482 362
rect 1606 358 1610 362
rect 1710 358 1714 362
rect 1718 358 1722 362
rect 1750 358 1754 362
rect 1806 358 1810 362
rect 1862 358 1866 362
rect 1934 358 1938 362
rect 1966 358 1970 362
rect 1998 358 2002 362
rect 2014 358 2018 362
rect 2062 358 2066 362
rect 2118 358 2122 362
rect 2150 358 2154 362
rect 2302 358 2306 362
rect 2334 358 2338 362
rect 2390 358 2394 362
rect 2438 358 2442 362
rect 2446 358 2450 362
rect 30 348 34 352
rect 78 348 82 352
rect 126 348 130 352
rect 198 348 202 352
rect 222 348 226 352
rect 238 348 242 352
rect 262 348 266 352
rect 270 348 274 352
rect 294 348 298 352
rect 326 348 330 352
rect 366 348 370 352
rect 406 348 410 352
rect 462 348 466 352
rect 478 348 482 352
rect 486 348 490 352
rect 550 348 554 352
rect 590 348 594 352
rect 646 348 650 352
rect 726 348 730 352
rect 742 348 746 352
rect 902 348 906 352
rect 926 348 930 352
rect 6 338 10 342
rect 22 338 26 342
rect 94 338 98 342
rect 174 338 178 342
rect 246 338 250 342
rect 254 338 258 342
rect 318 338 322 342
rect 398 338 402 342
rect 1006 347 1010 351
rect 1030 348 1034 352
rect 1102 347 1106 351
rect 1134 348 1138 352
rect 1198 347 1202 351
rect 1230 348 1234 352
rect 1294 347 1298 351
rect 1422 348 1426 352
rect 1438 348 1442 352
rect 1446 348 1450 352
rect 1502 348 1506 352
rect 1582 348 1586 352
rect 1734 348 1738 352
rect 1790 348 1794 352
rect 1822 348 1826 352
rect 1846 348 1850 352
rect 1918 348 1922 352
rect 1942 348 1946 352
rect 1974 348 1978 352
rect 2006 348 2010 352
rect 2046 348 2050 352
rect 2078 348 2082 352
rect 2094 348 2098 352
rect 2134 348 2138 352
rect 2158 348 2162 352
rect 2182 348 2186 352
rect 2214 348 2218 352
rect 2238 348 2242 352
rect 2262 348 2266 352
rect 2278 348 2282 352
rect 2310 348 2314 352
rect 2350 348 2354 352
rect 2382 348 2386 352
rect 2446 348 2450 352
rect 2462 348 2466 352
rect 2486 348 2490 352
rect 2510 358 2514 362
rect 2590 358 2594 362
rect 2662 358 2666 362
rect 2710 358 2714 362
rect 2750 358 2754 362
rect 2846 358 2850 362
rect 2582 348 2586 352
rect 2614 348 2618 352
rect 2654 348 2658 352
rect 2694 348 2698 352
rect 2710 348 2714 352
rect 2742 348 2746 352
rect 2766 348 2770 352
rect 2782 348 2786 352
rect 2814 348 2818 352
rect 2830 348 2834 352
rect 2854 348 2858 352
rect 2862 348 2866 352
rect 2886 348 2890 352
rect 2910 358 2914 362
rect 2958 358 2962 362
rect 3006 358 3010 362
rect 3014 358 3018 362
rect 3062 358 3066 362
rect 3190 358 3194 362
rect 3318 358 3322 362
rect 2934 348 2938 352
rect 3030 348 3034 352
rect 3078 348 3082 352
rect 3086 348 3090 352
rect 3102 348 3106 352
rect 3134 348 3138 352
rect 3142 348 3146 352
rect 3150 348 3154 352
rect 3174 348 3178 352
rect 3238 348 3242 352
rect 3246 348 3250 352
rect 3254 348 3258 352
rect 3278 348 3282 352
rect 3302 348 3306 352
rect 3398 358 3402 362
rect 3430 358 3434 362
rect 3438 358 3442 362
rect 3518 358 3522 362
rect 3526 358 3530 362
rect 3622 358 3626 362
rect 3630 358 3634 362
rect 3654 358 3658 362
rect 3734 358 3738 362
rect 3806 358 3810 362
rect 3838 358 3842 362
rect 3366 348 3370 352
rect 3414 348 3418 352
rect 3462 348 3466 352
rect 3494 348 3498 352
rect 3550 348 3554 352
rect 3678 348 3682 352
rect 3702 348 3706 352
rect 3718 348 3722 352
rect 3742 348 3746 352
rect 3758 348 3762 352
rect 3814 348 3818 352
rect 3838 348 3842 352
rect 3854 348 3858 352
rect 3886 348 3890 352
rect 4006 358 4010 362
rect 4054 358 4058 362
rect 4110 358 4114 362
rect 4326 358 4330 362
rect 4438 358 4442 362
rect 4502 358 4506 362
rect 4574 358 4578 362
rect 542 338 546 342
rect 566 338 570 342
rect 686 338 690 342
rect 766 338 770 342
rect 862 338 866 342
rect 1310 338 1314 342
rect 1366 338 1370 342
rect 1414 338 1418 342
rect 1454 338 1458 342
rect 1494 338 1498 342
rect 1510 338 1514 342
rect 1550 338 1554 342
rect 1566 338 1570 342
rect 1590 338 1594 342
rect 1638 338 1642 342
rect 1646 338 1650 342
rect 1694 338 1698 342
rect 1702 338 1706 342
rect 1726 338 1730 342
rect 1798 338 1802 342
rect 1838 338 1842 342
rect 1886 338 1890 342
rect 1918 338 1922 342
rect 1950 338 1954 342
rect 1982 338 1986 342
rect 1998 338 2002 342
rect 2054 338 2058 342
rect 2086 338 2090 342
rect 2142 338 2146 342
rect 2190 338 2194 342
rect 2206 338 2210 342
rect 2278 338 2282 342
rect 2286 338 2290 342
rect 2310 338 2314 342
rect 2318 338 2322 342
rect 2358 338 2362 342
rect 2382 338 2386 342
rect 2406 338 2410 342
rect 2414 338 2418 342
rect 2470 338 2474 342
rect 2478 338 2482 342
rect 2526 338 2530 342
rect 2558 338 2562 342
rect 2574 338 2578 342
rect 2598 338 2602 342
rect 2630 338 2634 342
rect 2662 338 2666 342
rect 2678 338 2682 342
rect 2686 338 2690 342
rect 2734 338 2738 342
rect 2782 338 2786 342
rect 2790 338 2794 342
rect 2822 338 2826 342
rect 2870 338 2874 342
rect 2878 338 2882 342
rect 2934 338 2938 342
rect 2982 338 2986 342
rect 3038 338 3042 342
rect 3086 338 3090 342
rect 3206 338 3210 342
rect 3294 338 3298 342
rect 3342 338 3346 342
rect 3374 338 3378 342
rect 3382 338 3386 342
rect 3406 338 3410 342
rect 3462 338 3466 342
rect 3470 338 3474 342
rect 3502 338 3506 342
rect 3542 338 3546 342
rect 3558 338 3562 342
rect 3590 338 3594 342
rect 3646 338 3650 342
rect 3678 338 3682 342
rect 3694 338 3698 342
rect 3710 338 3714 342
rect 3766 338 3770 342
rect 3782 338 3786 342
rect 3862 338 3866 342
rect 3942 348 3946 352
rect 3950 348 3954 352
rect 3966 348 3970 352
rect 3998 348 4002 352
rect 4038 348 4042 352
rect 4062 348 4066 352
rect 4118 348 4122 352
rect 4142 348 4146 352
rect 4174 348 4178 352
rect 4190 348 4194 352
rect 4230 348 4234 352
rect 4238 348 4242 352
rect 4286 348 4290 352
rect 4302 348 4306 352
rect 4318 348 4322 352
rect 4342 348 4346 352
rect 4374 348 4378 352
rect 4390 348 4394 352
rect 4414 348 4418 352
rect 4422 348 4426 352
rect 4534 348 4538 352
rect 3942 338 3946 342
rect 3958 338 3962 342
rect 3974 338 3978 342
rect 3982 338 3986 342
rect 3990 338 3994 342
rect 4006 338 4010 342
rect 4022 338 4026 342
rect 4030 338 4034 342
rect 4070 338 4074 342
rect 4166 338 4170 342
rect 4198 338 4202 342
rect 4222 338 4226 342
rect 4246 338 4250 342
rect 4270 338 4274 342
rect 4310 338 4314 342
rect 4350 338 4354 342
rect 4374 338 4378 342
rect 4414 338 4418 342
rect 4478 338 4482 342
rect 4494 338 4498 342
rect 4542 338 4546 342
rect 4550 338 4554 342
rect 30 328 34 332
rect 46 328 50 332
rect 166 328 170 332
rect 198 328 202 332
rect 214 328 218 332
rect 390 328 394 332
rect 446 328 450 332
rect 566 328 570 332
rect 702 328 706 332
rect 782 328 786 332
rect 1470 328 1474 332
rect 1526 328 1530 332
rect 1574 328 1578 332
rect 1758 328 1762 332
rect 1870 328 1874 332
rect 1910 328 1914 332
rect 2110 328 2114 332
rect 2222 328 2226 332
rect 2326 328 2330 332
rect 2366 328 2370 332
rect 2638 328 2642 332
rect 2718 328 2722 332
rect 2726 328 2730 332
rect 2806 328 2810 332
rect 2838 328 2842 332
rect 2966 328 2970 332
rect 3398 328 3402 332
rect 3574 328 3578 332
rect 3686 328 3690 332
rect 3742 328 3746 332
rect 3774 328 3778 332
rect 3870 328 3874 332
rect 3910 328 3914 332
rect 4078 328 4082 332
rect 4086 328 4090 332
rect 4158 328 4162 332
rect 4190 328 4194 332
rect 4206 328 4210 332
rect 4262 328 4266 332
rect 4270 328 4274 332
rect 4294 328 4298 332
rect 4358 328 4362 332
rect 4446 328 4450 332
rect 4494 328 4498 332
rect 118 318 122 322
rect 150 318 154 322
rect 206 318 210 322
rect 398 318 402 322
rect 454 318 458 322
rect 558 318 562 322
rect 870 318 874 322
rect 1070 318 1074 322
rect 1262 318 1266 322
rect 1358 318 1362 322
rect 1390 318 1394 322
rect 1462 318 1466 322
rect 1750 318 1754 322
rect 2502 318 2506 322
rect 2574 318 2578 322
rect 3222 318 3226 322
rect 3510 318 3514 322
rect 3534 318 3538 322
rect 3566 318 3570 322
rect 3630 318 3634 322
rect 4518 318 4522 322
rect 1002 303 1006 307
rect 1009 303 1013 307
rect 2026 303 2030 307
rect 2033 303 2037 307
rect 3050 303 3054 307
rect 3057 303 3061 307
rect 4082 303 4086 307
rect 4089 303 4093 307
rect 326 288 330 292
rect 758 288 762 292
rect 1054 288 1058 292
rect 1326 288 1330 292
rect 1422 288 1426 292
rect 1662 288 1666 292
rect 1686 288 1690 292
rect 1734 288 1738 292
rect 1758 288 1762 292
rect 1878 288 1882 292
rect 1910 288 1914 292
rect 1950 288 1954 292
rect 1966 288 1970 292
rect 1998 288 2002 292
rect 2014 288 2018 292
rect 2102 288 2106 292
rect 2126 288 2130 292
rect 2166 288 2170 292
rect 2222 288 2226 292
rect 2286 288 2290 292
rect 2302 288 2306 292
rect 2382 288 2386 292
rect 2510 288 2514 292
rect 2534 288 2538 292
rect 2606 288 2610 292
rect 2726 288 2730 292
rect 2750 288 2754 292
rect 2766 288 2770 292
rect 2814 288 2818 292
rect 2846 288 2850 292
rect 2918 288 2922 292
rect 2950 288 2954 292
rect 3014 288 3018 292
rect 3070 288 3074 292
rect 3086 288 3090 292
rect 3110 288 3114 292
rect 3126 288 3130 292
rect 3150 288 3154 292
rect 3262 288 3266 292
rect 3294 288 3298 292
rect 3318 288 3322 292
rect 3366 288 3370 292
rect 3406 288 3410 292
rect 3430 288 3434 292
rect 3478 288 3482 292
rect 3518 288 3522 292
rect 3566 288 3570 292
rect 3622 288 3626 292
rect 3662 288 3666 292
rect 3694 288 3698 292
rect 3710 288 3714 292
rect 3750 288 3754 292
rect 3822 288 3826 292
rect 3846 288 3850 292
rect 3982 288 3986 292
rect 4022 288 4026 292
rect 4054 288 4058 292
rect 4142 288 4146 292
rect 4182 288 4186 292
rect 4198 288 4202 292
rect 4246 288 4250 292
rect 4286 288 4290 292
rect 4342 288 4346 292
rect 4382 288 4386 292
rect 4398 288 4402 292
rect 4566 288 4570 292
rect 126 278 130 282
rect 486 278 490 282
rect 502 278 506 282
rect 582 278 586 282
rect 1166 278 1170 282
rect 1262 278 1266 282
rect 1494 278 1498 282
rect 1742 278 1746 282
rect 1830 278 1834 282
rect 1958 278 1962 282
rect 1990 278 1994 282
rect 2054 278 2058 282
rect 2070 278 2074 282
rect 2134 278 2138 282
rect 2294 278 2298 282
rect 2334 278 2338 282
rect 2350 278 2354 282
rect 2414 278 2418 282
rect 2462 278 2466 282
rect 2542 278 2546 282
rect 2662 278 2666 282
rect 2758 278 2762 282
rect 3382 278 3386 282
rect 3526 278 3530 282
rect 3686 278 3690 282
rect 3854 278 3858 282
rect 3894 278 3898 282
rect 3934 278 3938 282
rect 4110 278 4114 282
rect 4150 278 4154 282
rect 4190 278 4194 282
rect 4454 278 4458 282
rect 4502 278 4506 282
rect 4518 278 4522 282
rect 38 268 42 272
rect 86 268 90 272
rect 142 268 146 272
rect 158 268 162 272
rect 214 268 218 272
rect 262 268 266 272
rect 286 268 290 272
rect 318 268 322 272
rect 374 268 378 272
rect 406 268 410 272
rect 430 268 434 272
rect 454 268 458 272
rect 478 268 482 272
rect 542 268 546 272
rect 590 268 594 272
rect 622 268 626 272
rect 638 268 642 272
rect 646 268 650 272
rect 662 268 666 272
rect 702 268 706 272
rect 726 268 730 272
rect 774 268 778 272
rect 806 268 810 272
rect 846 268 850 272
rect 902 268 906 272
rect 934 268 938 272
rect 974 268 978 272
rect 1070 268 1074 272
rect 1086 268 1090 272
rect 1478 268 1482 272
rect 1550 268 1554 272
rect 1582 268 1586 272
rect 1670 268 1674 272
rect 1718 268 1722 272
rect 1750 268 1754 272
rect 1822 268 1826 272
rect 1830 268 1834 272
rect 1846 268 1850 272
rect 1886 268 1890 272
rect 1910 268 1914 272
rect 1926 268 1930 272
rect 1990 268 1994 272
rect 2030 268 2034 272
rect 2070 268 2074 272
rect 2110 268 2114 272
rect 2142 268 2146 272
rect 2174 268 2178 272
rect 2214 268 2218 272
rect 2238 268 2242 272
rect 2254 268 2258 272
rect 2270 268 2274 272
rect 2326 268 2330 272
rect 2358 268 2362 272
rect 2390 268 2394 272
rect 2422 268 2426 272
rect 2446 268 2450 272
rect 2486 268 2490 272
rect 2526 268 2530 272
rect 2566 268 2570 272
rect 2582 268 2586 272
rect 2630 268 2634 272
rect 2646 268 2650 272
rect 2702 268 2706 272
rect 2734 268 2738 272
rect 2774 268 2778 272
rect 2854 268 2858 272
rect 2886 268 2890 272
rect 2942 268 2946 272
rect 2958 268 2962 272
rect 2982 268 2986 272
rect 2990 268 2994 272
rect 3030 268 3034 272
rect 3038 268 3042 272
rect 3094 268 3098 272
rect 3126 268 3130 272
rect 3142 268 3146 272
rect 3174 268 3178 272
rect 3182 268 3186 272
rect 3198 268 3202 272
rect 3238 268 3242 272
rect 3310 268 3314 272
rect 3334 268 3338 272
rect 3342 268 3346 272
rect 3382 268 3386 272
rect 3390 268 3394 272
rect 3414 268 3418 272
rect 3438 268 3442 272
rect 3462 268 3466 272
rect 3470 268 3474 272
rect 3494 268 3498 272
rect 3550 268 3554 272
rect 3558 268 3562 272
rect 3598 268 3602 272
rect 3654 268 3658 272
rect 3678 268 3682 272
rect 3734 268 3738 272
rect 3758 268 3762 272
rect 3798 268 3802 272
rect 3838 268 3842 272
rect 3854 268 3858 272
rect 3886 268 3890 272
rect 3942 268 3946 272
rect 3958 268 3962 272
rect 3990 268 3994 272
rect 3998 268 4002 272
rect 4030 268 4034 272
rect 4062 268 4066 272
rect 4086 268 4090 272
rect 4118 268 4122 272
rect 4134 268 4138 272
rect 4158 268 4162 272
rect 4206 268 4210 272
rect 4222 268 4226 272
rect 4254 268 4258 272
rect 4318 268 4322 272
rect 4350 268 4354 272
rect 4422 268 4426 272
rect 4446 268 4450 272
rect 4486 268 4490 272
rect 4510 268 4514 272
rect 4542 268 4546 272
rect 22 258 26 262
rect 54 259 58 263
rect 134 258 138 262
rect 150 258 154 262
rect 166 258 170 262
rect 206 258 210 262
rect 238 258 242 262
rect 262 258 266 262
rect 294 258 298 262
rect 310 258 314 262
rect 358 258 362 262
rect 382 258 386 262
rect 486 258 490 262
rect 502 258 506 262
rect 558 258 562 262
rect 606 258 610 262
rect 678 258 682 262
rect 694 258 698 262
rect 798 258 802 262
rect 830 258 834 262
rect 854 258 858 262
rect 894 258 898 262
rect 926 258 930 262
rect 182 248 186 252
rect 238 248 242 252
rect 246 248 250 252
rect 6 238 10 242
rect 118 238 122 242
rect 230 238 234 242
rect 334 248 338 252
rect 366 248 370 252
rect 406 248 410 252
rect 422 248 426 252
rect 462 248 466 252
rect 550 248 554 252
rect 614 248 618 252
rect 622 248 626 252
rect 646 248 650 252
rect 662 248 666 252
rect 718 248 722 252
rect 782 248 786 252
rect 838 248 842 252
rect 870 248 874 252
rect 926 248 930 252
rect 982 258 986 262
rect 1006 258 1010 262
rect 1038 258 1042 262
rect 1094 258 1098 262
rect 1102 258 1106 262
rect 1118 258 1122 262
rect 1134 258 1138 262
rect 1166 259 1170 263
rect 1270 258 1274 262
rect 1358 259 1362 263
rect 1390 258 1394 262
rect 1606 258 1610 262
rect 1822 258 1826 262
rect 1854 258 1858 262
rect 1862 258 1866 262
rect 1894 258 1898 262
rect 1934 258 1938 262
rect 1942 258 1946 262
rect 2006 258 2010 262
rect 2046 258 2050 262
rect 2118 258 2122 262
rect 2134 258 2138 262
rect 2190 258 2194 262
rect 2230 258 2234 262
rect 2270 258 2274 262
rect 2318 258 2322 262
rect 2350 258 2354 262
rect 2366 258 2370 262
rect 2398 258 2402 262
rect 2414 258 2418 262
rect 2438 258 2442 262
rect 2454 258 2458 262
rect 2478 258 2482 262
rect 2494 258 2498 262
rect 2510 258 2514 262
rect 2606 258 2610 262
rect 2622 258 2626 262
rect 2638 258 2642 262
rect 2686 258 2690 262
rect 2710 258 2714 262
rect 2782 258 2786 262
rect 2790 258 2794 262
rect 2798 258 2802 262
rect 2822 258 2826 262
rect 2878 258 2882 262
rect 2894 258 2898 262
rect 2902 258 2906 262
rect 2926 258 2930 262
rect 3190 258 3194 262
rect 3214 258 3218 262
rect 3230 258 3234 262
rect 3246 258 3250 262
rect 3254 258 3258 262
rect 3350 258 3354 262
rect 3430 258 3434 262
rect 3454 258 3458 262
rect 3542 258 3546 262
rect 3606 258 3610 262
rect 3622 258 3626 262
rect 3662 258 3666 262
rect 3702 258 3706 262
rect 3726 258 3730 262
rect 3734 258 3738 262
rect 3774 258 3778 262
rect 3830 258 3834 262
rect 3878 258 3882 262
rect 3910 258 3914 262
rect 3934 258 3938 262
rect 3950 258 3954 262
rect 4006 258 4010 262
rect 4038 258 4042 262
rect 4054 258 4058 262
rect 4070 258 4074 262
rect 4110 258 4114 262
rect 4126 258 4130 262
rect 4166 258 4170 262
rect 4214 258 4218 262
rect 4230 258 4234 262
rect 4326 258 4330 262
rect 4358 258 4362 262
rect 4398 258 4402 262
rect 4438 258 4442 262
rect 4454 258 4458 262
rect 4470 258 4474 262
rect 4478 258 4482 262
rect 4518 258 4522 262
rect 4534 258 4538 262
rect 4542 258 4546 262
rect 966 248 970 252
rect 1046 248 1050 252
rect 1054 248 1058 252
rect 1110 248 1114 252
rect 1782 248 1786 252
rect 1966 248 1970 252
rect 2086 248 2090 252
rect 2094 248 2098 252
rect 2158 248 2162 252
rect 2182 248 2186 252
rect 2230 248 2234 252
rect 2262 248 2266 252
rect 2382 248 2386 252
rect 2454 248 2458 252
rect 2510 248 2514 252
rect 2598 248 2602 252
rect 2606 248 2610 252
rect 2662 248 2666 252
rect 2686 248 2690 252
rect 2726 248 2730 252
rect 2750 248 2754 252
rect 2838 248 2842 252
rect 2862 248 2866 252
rect 2878 248 2882 252
rect 2958 248 2962 252
rect 2966 248 2970 252
rect 3006 248 3010 252
rect 3014 248 3018 252
rect 3054 248 3058 252
rect 3102 248 3106 252
rect 3126 248 3130 252
rect 3150 248 3154 252
rect 3206 248 3210 252
rect 3214 248 3218 252
rect 3294 248 3298 252
rect 3318 248 3322 252
rect 3366 248 3370 252
rect 3406 248 3410 252
rect 3430 248 3434 252
rect 3486 248 3490 252
rect 3518 248 3522 252
rect 3526 248 3530 252
rect 3590 248 3594 252
rect 3630 248 3634 252
rect 3646 248 3650 252
rect 3662 248 3666 252
rect 3710 248 3714 252
rect 3790 248 3794 252
rect 3822 248 3826 252
rect 3862 248 3866 252
rect 3966 248 3970 252
rect 3974 248 3978 252
rect 4022 248 4026 252
rect 4182 248 4186 252
rect 4246 248 4250 252
rect 4262 248 4266 252
rect 4278 248 4282 252
rect 4302 248 4306 252
rect 4382 248 4386 252
rect 4390 248 4394 252
rect 4422 248 4426 252
rect 270 238 274 242
rect 350 238 354 242
rect 798 238 802 242
rect 822 238 826 242
rect 894 238 898 242
rect 910 238 914 242
rect 950 238 954 242
rect 958 238 962 242
rect 998 238 1002 242
rect 1030 238 1034 242
rect 1086 238 1090 242
rect 1126 238 1130 242
rect 1230 238 1234 242
rect 2198 238 2202 242
rect 2678 238 2682 242
rect 3438 238 3442 242
rect 4406 238 4410 242
rect 206 228 210 232
rect 2574 228 2578 232
rect 2686 228 2690 232
rect 222 218 226 222
rect 294 218 298 222
rect 358 218 362 222
rect 382 218 386 222
rect 534 218 538 222
rect 814 218 818 222
rect 958 218 962 222
rect 1038 218 1042 222
rect 1454 218 1458 222
rect 2190 218 2194 222
rect 2742 218 2746 222
rect 2998 218 3002 222
rect 4470 218 4474 222
rect 4502 218 4506 222
rect 498 203 502 207
rect 505 203 509 207
rect 1522 203 1526 207
rect 1529 203 1533 207
rect 2546 203 2550 207
rect 2553 203 2557 207
rect 3570 203 3574 207
rect 3577 203 3581 207
rect 102 188 106 192
rect 654 188 658 192
rect 846 188 850 192
rect 950 188 954 192
rect 1078 188 1082 192
rect 1758 188 1762 192
rect 1854 188 1858 192
rect 1974 188 1978 192
rect 2350 188 2354 192
rect 2358 188 2362 192
rect 2438 188 2442 192
rect 2470 188 2474 192
rect 2510 188 2514 192
rect 2534 188 2538 192
rect 2598 188 2602 192
rect 2638 188 2642 192
rect 2678 188 2682 192
rect 2798 188 2802 192
rect 2838 188 2842 192
rect 2894 188 2898 192
rect 2934 188 2938 192
rect 2958 188 2962 192
rect 3022 188 3026 192
rect 3046 188 3050 192
rect 3086 188 3090 192
rect 3126 188 3130 192
rect 3150 188 3154 192
rect 3214 188 3218 192
rect 3294 188 3298 192
rect 3366 188 3370 192
rect 3398 188 3402 192
rect 3622 188 3626 192
rect 3678 188 3682 192
rect 3766 188 3770 192
rect 3862 188 3866 192
rect 3910 188 3914 192
rect 3958 188 3962 192
rect 4046 188 4050 192
rect 4102 188 4106 192
rect 4222 188 4226 192
rect 4238 188 4242 192
rect 4310 188 4314 192
rect 4342 188 4346 192
rect 4414 188 4418 192
rect 4454 188 4458 192
rect 4494 188 4498 192
rect 4518 188 4522 192
rect 4558 188 4562 192
rect 566 178 570 182
rect 3942 178 3946 182
rect 214 168 218 172
rect 238 168 242 172
rect 246 168 250 172
rect 342 168 346 172
rect 382 168 386 172
rect 854 168 858 172
rect 942 168 946 172
rect 1086 168 1090 172
rect 1334 168 1338 172
rect 2774 168 2778 172
rect 3166 168 3170 172
rect 3806 168 3810 172
rect 3870 168 3874 172
rect 4086 168 4090 172
rect 4366 168 4370 172
rect 198 158 202 162
rect 366 158 370 162
rect 390 158 394 162
rect 550 158 554 162
rect 582 158 586 162
rect 638 158 642 162
rect 38 148 42 152
rect 70 147 74 151
rect 134 148 138 152
rect 166 147 170 151
rect 206 148 210 152
rect 222 148 226 152
rect 230 148 234 152
rect 238 148 242 152
rect 350 148 354 152
rect 358 148 362 152
rect 374 148 378 152
rect 422 147 426 151
rect 510 148 514 152
rect 574 148 578 152
rect 622 148 626 152
rect 630 148 634 152
rect 654 148 658 152
rect 678 158 682 162
rect 926 158 930 162
rect 1102 158 1106 162
rect 702 148 706 152
rect 718 148 722 152
rect 774 148 778 152
rect 86 138 90 142
rect 262 138 266 142
rect 326 138 330 142
rect 342 138 346 142
rect 406 138 410 142
rect 534 138 538 142
rect 558 138 562 142
rect 598 138 602 142
rect 614 138 618 142
rect 646 138 650 142
rect 694 138 698 142
rect 806 147 810 151
rect 838 148 842 152
rect 846 148 850 152
rect 870 148 874 152
rect 902 148 906 152
rect 918 148 922 152
rect 950 148 954 152
rect 958 148 962 152
rect 1014 148 1018 152
rect 1030 148 1034 152
rect 1094 148 1098 152
rect 1174 148 1178 152
rect 1182 148 1186 152
rect 1198 158 1202 162
rect 1222 158 1226 162
rect 1238 158 1242 162
rect 1862 158 1866 162
rect 878 138 882 142
rect 1110 138 1114 142
rect 1158 138 1162 142
rect 1270 147 1274 151
rect 1294 148 1298 152
rect 1342 148 1346 152
rect 1366 148 1370 152
rect 1430 148 1434 152
rect 1526 147 1530 151
rect 1558 148 1562 152
rect 1694 147 1698 151
rect 1798 148 1802 152
rect 1910 147 1914 151
rect 2006 148 2010 152
rect 2046 158 2050 162
rect 2166 158 2170 162
rect 2206 158 2210 162
rect 2278 158 2282 162
rect 2382 158 2386 162
rect 2422 158 2426 162
rect 2454 158 2458 162
rect 2062 148 2066 152
rect 2078 148 2082 152
rect 2102 148 2106 152
rect 2126 148 2130 152
rect 2150 148 2154 152
rect 2158 148 2162 152
rect 2206 148 2210 152
rect 2238 148 2242 152
rect 2254 148 2258 152
rect 2318 148 2322 152
rect 2350 148 2354 152
rect 2358 148 2362 152
rect 2374 148 2378 152
rect 2438 148 2442 152
rect 2462 148 2466 152
rect 2494 148 2498 152
rect 2558 158 2562 162
rect 2574 158 2578 162
rect 2702 158 2706 162
rect 2750 158 2754 162
rect 2758 158 2762 162
rect 2806 158 2810 162
rect 2878 158 2882 162
rect 2926 158 2930 162
rect 2974 158 2978 162
rect 3006 158 3010 162
rect 3030 158 3034 162
rect 3102 158 3106 162
rect 3110 158 3114 162
rect 3142 158 3146 162
rect 3182 158 3186 162
rect 3246 158 3250 162
rect 3254 158 3258 162
rect 3270 158 3274 162
rect 2534 148 2538 152
rect 2550 148 2554 152
rect 2622 148 2626 152
rect 2630 148 2634 152
rect 2662 148 2666 152
rect 2686 148 2690 152
rect 2694 148 2698 152
rect 2718 148 2722 152
rect 2734 148 2738 152
rect 2750 148 2754 152
rect 2774 148 2778 152
rect 2838 148 2842 152
rect 2950 148 2954 152
rect 2958 148 2962 152
rect 2990 148 2994 152
rect 3054 148 3058 152
rect 3086 148 3090 152
rect 3126 148 3130 152
rect 3230 148 3234 152
rect 3238 148 3242 152
rect 3270 148 3274 152
rect 3286 148 3290 152
rect 3318 158 3322 162
rect 3350 158 3354 162
rect 3518 158 3522 162
rect 3638 158 3642 162
rect 3702 158 3706 162
rect 3790 158 3794 162
rect 3822 158 3826 162
rect 3854 158 3858 162
rect 3334 148 3338 152
rect 3366 148 3370 152
rect 3382 148 3386 152
rect 3414 148 3418 152
rect 3422 148 3426 152
rect 3430 148 3434 152
rect 3462 148 3466 152
rect 3486 148 3490 152
rect 3518 148 3522 152
rect 3550 148 3554 152
rect 3574 148 3578 152
rect 3590 148 3594 152
rect 3622 148 3626 152
rect 1214 138 1218 142
rect 1598 138 1602 142
rect 1662 138 1666 142
rect 1678 138 1682 142
rect 1710 138 1714 142
rect 1774 138 1778 142
rect 1878 138 1882 142
rect 1894 138 1898 142
rect 2014 138 2018 142
rect 2062 138 2066 142
rect 2182 138 2186 142
rect 2246 138 2250 142
rect 2262 138 2266 142
rect 2294 138 2298 142
rect 2310 138 2314 142
rect 2398 138 2402 142
rect 2406 138 2410 142
rect 2430 138 2434 142
rect 2470 138 2474 142
rect 2486 138 2490 142
rect 2518 138 2522 142
rect 2590 138 2594 142
rect 2614 138 2618 142
rect 2718 138 2722 142
rect 2782 138 2786 142
rect 2790 138 2794 142
rect 2862 138 2866 142
rect 2918 138 2922 142
rect 2942 138 2946 142
rect 2982 138 2986 142
rect 3062 138 3066 142
rect 3078 138 3082 142
rect 3134 138 3138 142
rect 3166 138 3170 142
rect 3198 138 3202 142
rect 3222 138 3226 142
rect 3278 138 3282 142
rect 3286 138 3290 142
rect 3342 138 3346 142
rect 3374 138 3378 142
rect 3438 138 3442 142
rect 3478 138 3482 142
rect 3510 138 3514 142
rect 3534 138 3538 142
rect 3662 148 3666 152
rect 3686 148 3690 152
rect 3694 148 3698 152
rect 3718 148 3722 152
rect 3734 148 3738 152
rect 3774 148 3778 152
rect 3798 148 3802 152
rect 3830 148 3834 152
rect 3838 148 3842 152
rect 3862 148 3866 152
rect 3886 148 3890 152
rect 3926 148 3930 152
rect 3942 148 3946 152
rect 3982 148 3986 152
rect 4054 158 4058 162
rect 4118 158 4122 162
rect 4134 158 4138 162
rect 4006 148 4010 152
rect 4022 148 4026 152
rect 4078 148 4082 152
rect 4118 148 4122 152
rect 4158 148 4162 152
rect 4326 158 4330 162
rect 4382 158 4386 162
rect 4510 158 4514 162
rect 4190 148 4194 152
rect 4198 148 4202 152
rect 4238 148 4242 152
rect 4254 148 4258 152
rect 4278 148 4282 152
rect 4294 148 4298 152
rect 4318 148 4322 152
rect 4342 148 4346 152
rect 4358 148 4362 152
rect 4422 148 4426 152
rect 4438 148 4442 152
rect 4454 148 4458 152
rect 4470 148 4474 152
rect 4518 148 4522 152
rect 4542 148 4546 152
rect 3710 138 3714 142
rect 3726 138 3730 142
rect 3750 138 3754 142
rect 3798 138 3802 142
rect 3894 138 3898 142
rect 3918 138 3922 142
rect 3950 138 3954 142
rect 3974 138 3978 142
rect 3998 138 4002 142
rect 4014 138 4018 142
rect 4030 138 4034 142
rect 4070 138 4074 142
rect 4094 138 4098 142
rect 4126 138 4130 142
rect 4150 138 4154 142
rect 4166 138 4170 142
rect 4190 138 4194 142
rect 4206 138 4210 142
rect 4230 138 4234 142
rect 4262 138 4266 142
rect 4286 138 4290 142
rect 4350 138 4354 142
rect 4358 138 4362 142
rect 4398 138 4402 142
rect 4446 138 4450 142
rect 4478 138 4482 142
rect 606 128 610 132
rect 702 128 706 132
rect 894 128 898 132
rect 1046 128 1050 132
rect 1454 128 1458 132
rect 1982 128 1986 132
rect 2230 128 2234 132
rect 2334 128 2338 132
rect 2374 128 2378 132
rect 2598 128 2602 132
rect 2646 128 2650 132
rect 2814 128 2818 132
rect 3190 128 3194 132
rect 3454 128 3458 132
rect 3566 128 3570 132
rect 3606 128 3610 132
rect 3630 128 3634 132
rect 3750 128 3754 132
rect 3782 128 3786 132
rect 3846 128 3850 132
rect 3910 128 3914 132
rect 3958 128 3962 132
rect 4046 128 4050 132
rect 4222 128 4226 132
rect 4270 128 4274 132
rect 4302 128 4306 132
rect 4414 128 4418 132
rect 4438 128 4442 132
rect 4534 128 4538 132
rect 6 118 10 122
rect 486 118 490 122
rect 526 118 530 122
rect 742 118 746 122
rect 974 118 978 122
rect 1358 118 1362 122
rect 1382 118 1386 122
rect 1390 118 1394 122
rect 1590 118 1594 122
rect 1862 118 1866 122
rect 2094 118 2098 122
rect 2142 118 2146 122
rect 2422 118 2426 122
rect 3518 118 3522 122
rect 1002 103 1006 107
rect 1009 103 1013 107
rect 2026 103 2030 107
rect 2033 103 2037 107
rect 3050 103 3054 107
rect 3057 103 3061 107
rect 4082 103 4086 107
rect 4089 103 4093 107
rect 38 88 42 92
rect 214 88 218 92
rect 454 88 458 92
rect 518 88 522 92
rect 734 88 738 92
rect 790 88 794 92
rect 926 88 930 92
rect 1110 88 1114 92
rect 1526 88 1530 92
rect 1878 88 1882 92
rect 1910 88 1914 92
rect 1926 88 1930 92
rect 1950 88 1954 92
rect 1998 88 2002 92
rect 2046 88 2050 92
rect 2110 88 2114 92
rect 2174 88 2178 92
rect 2206 88 2210 92
rect 2238 88 2242 92
rect 2270 88 2274 92
rect 2374 88 2378 92
rect 2574 88 2578 92
rect 2598 88 2602 92
rect 2614 88 2618 92
rect 2694 88 2698 92
rect 2718 88 2722 92
rect 2878 88 2882 92
rect 2918 88 2922 92
rect 2998 88 3002 92
rect 3134 88 3138 92
rect 3182 88 3186 92
rect 3222 88 3226 92
rect 3294 88 3298 92
rect 3358 88 3362 92
rect 3374 88 3378 92
rect 3446 88 3450 92
rect 3470 88 3474 92
rect 3494 88 3498 92
rect 3526 88 3530 92
rect 3542 88 3546 92
rect 3590 88 3594 92
rect 3614 88 3618 92
rect 3670 88 3674 92
rect 3734 88 3738 92
rect 4014 88 4018 92
rect 4102 88 4106 92
rect 4214 88 4218 92
rect 4542 88 4546 92
rect 182 78 186 82
rect 1046 78 1050 82
rect 1454 78 1458 82
rect 1646 78 1650 82
rect 1710 78 1714 82
rect 1830 78 1834 82
rect 1886 78 1890 82
rect 2006 78 2010 82
rect 2078 78 2082 82
rect 2158 78 2162 82
rect 94 68 98 72
rect 134 68 138 72
rect 406 68 410 72
rect 574 68 578 72
rect 654 68 658 72
rect 806 68 810 72
rect 846 68 850 72
rect 1294 68 1298 72
rect 1630 68 1634 72
rect 22 58 26 62
rect 118 58 122 62
rect 150 59 154 63
rect 278 58 282 62
rect 310 59 314 63
rect 358 58 362 62
rect 390 59 394 63
rect 462 58 466 62
rect 518 58 522 62
rect 574 58 578 62
rect 622 58 626 62
rect 670 59 674 63
rect 758 58 762 62
rect 782 58 786 62
rect 830 58 834 62
rect 862 59 866 63
rect 934 58 938 62
rect 958 58 962 62
rect 982 58 986 62
rect 1046 59 1050 63
rect 1134 58 1138 62
rect 1166 59 1170 63
rect 1198 58 1202 62
rect 1310 58 1314 62
rect 1382 58 1386 62
rect 1406 58 1410 62
rect 1462 58 1466 62
rect 1526 58 1530 62
rect 1566 58 1570 62
rect 1614 59 1618 63
rect 1918 68 1922 72
rect 1974 68 1978 72
rect 1982 68 1986 72
rect 2070 68 2074 72
rect 2102 68 2106 72
rect 2134 68 2138 72
rect 2358 78 2362 82
rect 2382 78 2386 82
rect 2414 78 2418 82
rect 2430 78 2434 82
rect 2470 78 2474 82
rect 2654 78 2658 82
rect 2686 78 2690 82
rect 2734 78 2738 82
rect 2910 78 2914 82
rect 2926 78 2930 82
rect 2974 78 2978 82
rect 3094 78 3098 82
rect 3190 78 3194 82
rect 3254 78 3258 82
rect 3270 78 3274 82
rect 3318 78 3322 82
rect 3350 78 3354 82
rect 3478 78 3482 82
rect 3550 78 3554 82
rect 3654 78 3658 82
rect 3758 78 3762 82
rect 3870 78 3874 82
rect 4070 78 4074 82
rect 4110 78 4114 82
rect 4286 78 4290 82
rect 4310 78 4314 82
rect 4326 78 4330 82
rect 4342 78 4346 82
rect 4366 78 4370 82
rect 4390 78 4394 82
rect 4478 78 4482 82
rect 4534 78 4538 82
rect 2182 68 2186 72
rect 2214 68 2218 72
rect 2222 68 2226 72
rect 2310 68 2314 72
rect 2398 68 2402 72
rect 2414 68 2418 72
rect 2502 68 2506 72
rect 2534 68 2538 72
rect 2582 68 2586 72
rect 2622 68 2626 72
rect 2630 68 2634 72
rect 2662 68 2666 72
rect 2766 68 2770 72
rect 2782 68 2786 72
rect 2846 68 2850 72
rect 2854 68 2858 72
rect 2886 68 2890 72
rect 2982 68 2986 72
rect 3038 68 3042 72
rect 3102 68 3106 72
rect 3142 68 3146 72
rect 3158 68 3162 72
rect 3166 68 3170 72
rect 3206 68 3210 72
rect 3230 68 3234 72
rect 3254 68 3258 72
rect 3278 68 3282 72
rect 3318 68 3322 72
rect 3390 68 3394 72
rect 3398 68 3402 72
rect 3422 68 3426 72
rect 3454 68 3458 72
rect 3510 68 3514 72
rect 3550 68 3554 72
rect 3598 68 3602 72
rect 3622 68 3626 72
rect 3678 68 3682 72
rect 3702 68 3706 72
rect 3766 68 3770 72
rect 3790 68 3794 72
rect 3846 68 3850 72
rect 3862 68 3866 72
rect 3878 68 3882 72
rect 3894 68 3898 72
rect 3910 68 3914 72
rect 3926 68 3930 72
rect 3958 68 3962 72
rect 3990 68 3994 72
rect 4030 68 4034 72
rect 4062 68 4066 72
rect 4118 68 4122 72
rect 4158 68 4162 72
rect 4174 68 4178 72
rect 4190 68 4194 72
rect 4254 68 4258 72
rect 4278 68 4282 72
rect 4326 68 4330 72
rect 4374 68 4378 72
rect 4398 68 4402 72
rect 4446 68 4450 72
rect 4454 68 4458 72
rect 4478 68 4482 72
rect 4558 68 4562 72
rect 1718 58 1722 62
rect 1790 58 1794 62
rect 1798 58 1802 62
rect 1814 58 1818 62
rect 1822 58 1826 62
rect 1854 58 1858 62
rect 1870 58 1874 62
rect 1942 58 1946 62
rect 2022 58 2026 62
rect 2062 58 2066 62
rect 2078 58 2082 62
rect 2094 58 2098 62
rect 2110 58 2114 62
rect 2126 58 2130 62
rect 2142 58 2146 62
rect 2158 58 2162 62
rect 2246 58 2250 62
rect 2254 58 2258 62
rect 2286 58 2290 62
rect 2334 58 2338 62
rect 2366 58 2370 62
rect 2390 58 2394 62
rect 2454 58 2458 62
rect 2526 58 2530 62
rect 2534 58 2538 62
rect 2558 58 2562 62
rect 2638 58 2642 62
rect 2702 58 2706 62
rect 2758 58 2762 62
rect 2798 58 2802 62
rect 2814 58 2818 62
rect 2838 58 2842 62
rect 2942 58 2946 62
rect 3006 58 3010 62
rect 3022 58 3026 62
rect 3070 58 3074 62
rect 3126 58 3130 62
rect 3302 58 3306 62
rect 3366 58 3370 62
rect 3422 58 3426 62
rect 3462 58 3466 62
rect 3502 58 3506 62
rect 3534 58 3538 62
rect 3638 58 3642 62
rect 3654 58 3658 62
rect 3710 58 3714 62
rect 3718 58 3722 62
rect 3742 58 3746 62
rect 3798 58 3802 62
rect 3846 58 3850 62
rect 3854 58 3858 62
rect 3886 58 3890 62
rect 3902 58 3906 62
rect 3918 58 3922 62
rect 3934 58 3938 62
rect 3950 58 3954 62
rect 3982 58 3986 62
rect 3998 58 4002 62
rect 4038 58 4042 62
rect 4054 58 4058 62
rect 4070 58 4074 62
rect 4126 58 4130 62
rect 4150 58 4154 62
rect 4182 58 4186 62
rect 4246 58 4250 62
rect 4294 58 4298 62
rect 4342 58 4346 62
rect 4366 58 4370 62
rect 4374 58 4378 62
rect 4406 58 4410 62
rect 4414 58 4418 62
rect 4494 58 4498 62
rect 4526 58 4530 62
rect 4550 58 4554 62
rect 4558 58 4562 62
rect 790 48 794 52
rect 1870 48 1874 52
rect 1910 48 1914 52
rect 1998 48 2002 52
rect 2198 48 2202 52
rect 2238 48 2242 52
rect 2486 48 2490 52
rect 2526 48 2530 52
rect 2574 48 2578 52
rect 2598 48 2602 52
rect 2678 48 2682 52
rect 2798 48 2802 52
rect 2902 48 2906 52
rect 2950 48 2954 52
rect 2966 48 2970 52
rect 3038 48 3042 52
rect 3046 48 3050 52
rect 3118 48 3122 52
rect 3182 48 3186 52
rect 3222 48 3226 52
rect 3246 48 3250 52
rect 3294 48 3298 52
rect 3342 48 3346 52
rect 3398 48 3402 52
rect 3414 48 3418 52
rect 3438 48 3442 52
rect 3526 48 3530 52
rect 3574 48 3578 52
rect 3614 48 3618 52
rect 3702 48 3706 52
rect 3782 48 3786 52
rect 3814 48 3818 52
rect 3822 48 3826 52
rect 3934 48 3938 52
rect 3966 48 3970 52
rect 4230 48 4234 52
rect 4430 48 4434 52
rect 4470 48 4474 52
rect 4582 48 4586 52
rect 6 38 10 42
rect 2030 38 2034 42
rect 2334 38 2338 42
rect 3014 38 3018 42
rect 3302 38 3306 42
rect 3798 38 3802 42
rect 4566 38 4570 42
rect 3110 28 3114 32
rect 3334 28 3338 32
rect 4142 28 4146 32
rect 4486 28 4490 32
rect 102 18 106 22
rect 222 18 226 22
rect 342 18 346 22
rect 478 18 482 22
rect 486 18 490 22
rect 638 18 642 22
rect 742 18 746 22
rect 766 18 770 22
rect 814 18 818 22
rect 950 18 954 22
rect 974 18 978 22
rect 998 18 1002 22
rect 1118 18 1122 22
rect 1254 18 1258 22
rect 1374 18 1378 22
rect 1398 18 1402 22
rect 1422 18 1426 22
rect 1558 18 1562 22
rect 1582 18 1586 22
rect 3086 18 3090 22
rect 4054 18 4058 22
rect 4158 18 4162 22
rect 4262 18 4266 22
rect 498 3 502 7
rect 505 3 509 7
rect 1522 3 1526 7
rect 1529 3 1533 7
rect 2546 3 2550 7
rect 2553 3 2557 7
rect 3570 3 3574 7
rect 3577 3 3581 7
<< metal2 >>
rect 150 4431 154 4432
rect 150 4428 161 4431
rect 34 4358 38 4361
rect 114 4348 118 4351
rect 6 4332 9 4348
rect 26 4338 30 4341
rect 58 4338 62 4341
rect 6 4252 9 4278
rect 26 4268 30 4271
rect 58 4268 62 4271
rect 46 4262 49 4268
rect 70 4262 73 4348
rect 106 4338 110 4341
rect 158 4332 161 4428
rect 1998 4428 2002 4432
rect 2262 4431 2266 4432
rect 2750 4431 2754 4432
rect 2774 4431 2778 4432
rect 3134 4431 3138 4432
rect 3158 4431 3162 4432
rect 2262 4428 2273 4431
rect 496 4403 498 4407
rect 502 4403 505 4407
rect 509 4403 512 4407
rect 1520 4403 1522 4407
rect 1526 4403 1529 4407
rect 1533 4403 1536 4407
rect 1998 4402 2001 4428
rect 2270 4392 2273 4428
rect 2742 4428 2754 4431
rect 2766 4428 2778 4431
rect 3126 4428 3138 4431
rect 3150 4428 3162 4431
rect 3182 4431 3186 4432
rect 3206 4431 3210 4432
rect 3286 4431 3290 4432
rect 3326 4431 3330 4432
rect 3382 4431 3386 4432
rect 3406 4431 3410 4432
rect 3462 4431 3466 4432
rect 3182 4428 3193 4431
rect 3206 4428 3217 4431
rect 3286 4428 3297 4431
rect 2544 4403 2546 4407
rect 2550 4403 2553 4407
rect 2557 4403 2560 4407
rect 2742 4392 2745 4428
rect 2766 4392 2769 4428
rect 3126 4392 3129 4428
rect 3150 4392 3153 4428
rect 3190 4392 3193 4428
rect 3214 4392 3217 4428
rect 3294 4392 3297 4428
rect 3318 4428 3330 4431
rect 3374 4428 3386 4431
rect 3398 4428 3410 4431
rect 3454 4428 3466 4431
rect 3518 4431 3522 4432
rect 3518 4428 3529 4431
rect 3318 4392 3321 4428
rect 3374 4392 3377 4428
rect 3398 4392 3401 4428
rect 3454 4392 3457 4428
rect 3526 4392 3529 4428
rect 3558 4428 3562 4432
rect 3686 4428 3690 4432
rect 3750 4428 3754 4432
rect 3766 4428 3770 4432
rect 3790 4428 3794 4432
rect 3830 4428 3834 4432
rect 3878 4428 3882 4432
rect 3902 4431 3906 4432
rect 3894 4428 3906 4431
rect 3918 4428 3922 4432
rect 3942 4428 3946 4432
rect 3966 4428 3970 4432
rect 3982 4428 3986 4432
rect 4006 4428 4010 4432
rect 4022 4428 4026 4432
rect 4046 4431 4050 4432
rect 4038 4428 4050 4431
rect 4062 4428 4066 4432
rect 4102 4428 4106 4432
rect 4126 4428 4130 4432
rect 4142 4428 4146 4432
rect 4214 4428 4218 4432
rect 4230 4428 4234 4432
rect 4342 4428 4346 4432
rect 4382 4428 4386 4432
rect 4430 4428 4434 4432
rect 2026 4378 2030 4381
rect 774 4362 777 4368
rect 1510 4362 1513 4368
rect 794 4358 798 4361
rect 930 4358 937 4361
rect 190 4351 193 4358
rect 546 4348 550 4351
rect 286 4342 289 4347
rect 406 4342 409 4348
rect 462 4342 465 4348
rect 614 4342 617 4348
rect 586 4338 590 4341
rect 270 4332 273 4338
rect 78 4282 81 4328
rect 126 4322 129 4328
rect 30 4192 33 4248
rect 54 4152 57 4258
rect 46 4148 54 4151
rect 6 4132 9 4148
rect 26 4138 30 4141
rect 6 3932 9 3968
rect 6 3852 9 3878
rect 30 3872 33 4068
rect 38 4022 41 4058
rect 46 3952 49 4148
rect 58 4138 62 4141
rect 78 4132 81 4278
rect 190 4272 193 4328
rect 110 4263 113 4268
rect 142 4262 145 4268
rect 190 4262 193 4268
rect 114 4158 118 4161
rect 86 4142 89 4148
rect 134 4142 137 4178
rect 70 3992 73 4018
rect 50 3948 54 3951
rect 70 3932 73 3938
rect 78 3932 81 4128
rect 142 4102 145 4258
rect 206 4252 209 4259
rect 174 4202 177 4218
rect 230 4202 233 4288
rect 254 4272 257 4318
rect 350 4312 353 4318
rect 358 4302 361 4338
rect 338 4288 361 4291
rect 358 4282 361 4288
rect 350 4272 353 4278
rect 298 4268 302 4271
rect 374 4262 377 4318
rect 406 4292 409 4298
rect 414 4292 417 4338
rect 438 4282 441 4298
rect 382 4272 385 4278
rect 430 4262 433 4268
rect 446 4261 449 4318
rect 458 4278 462 4281
rect 446 4258 454 4261
rect 302 4252 305 4258
rect 174 4152 177 4158
rect 214 4152 217 4158
rect 230 4152 233 4198
rect 254 4192 257 4238
rect 254 4162 257 4168
rect 250 4158 254 4161
rect 262 4152 265 4248
rect 374 4242 377 4248
rect 270 4212 273 4218
rect 366 4192 369 4238
rect 430 4232 433 4258
rect 510 4242 513 4258
rect 514 4238 521 4241
rect 466 4228 470 4231
rect 446 4192 449 4198
rect 318 4152 321 4158
rect 230 4142 233 4148
rect 246 4138 254 4141
rect 182 4132 185 4138
rect 194 4128 198 4131
rect 182 4102 185 4118
rect 206 4112 209 4138
rect 238 4132 241 4138
rect 218 4128 222 4131
rect 246 4121 249 4138
rect 262 4131 265 4148
rect 286 4142 289 4148
rect 258 4128 265 4131
rect 238 4118 249 4121
rect 110 4092 113 4098
rect 178 4078 182 4081
rect 178 4068 182 4071
rect 42 3928 46 3931
rect 94 3882 97 4018
rect 78 3862 81 3868
rect 14 3752 17 3818
rect 34 3758 38 3761
rect 6 3732 9 3748
rect 26 3738 30 3741
rect 38 3682 41 3688
rect 46 3682 49 3859
rect 58 3738 62 3741
rect 86 3682 89 3728
rect 6 3672 9 3678
rect 50 3658 54 3661
rect 70 3652 73 3678
rect 6 3532 9 3548
rect 22 3542 25 3548
rect 62 3542 65 3548
rect 74 3538 78 3541
rect 86 3532 89 3678
rect 94 3662 97 3748
rect 102 3732 105 3928
rect 110 3892 113 4018
rect 166 3982 169 4068
rect 190 4062 193 4068
rect 198 4062 201 4068
rect 206 4062 209 4108
rect 222 4072 225 4088
rect 230 4072 233 4078
rect 214 4062 217 4068
rect 238 4062 241 4118
rect 270 4072 273 4138
rect 294 4132 297 4138
rect 286 4122 289 4128
rect 302 4122 305 4138
rect 310 4132 313 4138
rect 126 3752 129 3948
rect 206 3942 209 3948
rect 214 3932 217 4018
rect 222 3931 225 3948
rect 230 3942 233 4058
rect 238 3992 241 4058
rect 246 4052 249 4058
rect 254 4022 257 4068
rect 270 4012 273 4058
rect 294 4031 297 4098
rect 302 4072 305 4118
rect 318 4112 321 4148
rect 326 4142 329 4168
rect 338 4138 342 4141
rect 350 4132 353 4148
rect 366 4142 369 4188
rect 382 4151 385 4158
rect 314 4078 318 4081
rect 310 4072 313 4078
rect 326 4062 329 4128
rect 334 4102 337 4118
rect 350 4092 353 4128
rect 382 4082 385 4108
rect 310 4032 313 4058
rect 326 4032 329 4058
rect 342 4052 345 4058
rect 294 4028 305 4031
rect 286 3992 289 4008
rect 254 3952 257 3988
rect 270 3952 273 3968
rect 294 3952 297 4018
rect 302 3952 305 4028
rect 262 3942 265 3948
rect 282 3938 286 3941
rect 298 3938 302 3941
rect 222 3928 233 3931
rect 206 3922 209 3928
rect 142 3863 145 3918
rect 230 3892 233 3928
rect 310 3922 313 3938
rect 214 3872 217 3878
rect 318 3872 321 4008
rect 330 3958 334 3961
rect 326 3932 329 3938
rect 334 3922 337 3948
rect 342 3932 345 4018
rect 350 3992 353 4068
rect 374 4062 377 4068
rect 362 4058 366 4061
rect 362 4048 366 4051
rect 374 4022 377 4038
rect 350 3972 353 3978
rect 358 3942 361 3948
rect 374 3942 377 3948
rect 382 3942 385 4078
rect 390 3972 393 4018
rect 398 3992 401 4128
rect 430 4122 433 4178
rect 430 4075 433 4118
rect 446 4092 449 4148
rect 454 4142 457 4228
rect 478 4192 481 4228
rect 496 4203 498 4207
rect 502 4203 505 4207
rect 509 4203 512 4207
rect 446 4072 449 4088
rect 426 4038 430 4041
rect 406 3942 409 4028
rect 454 3982 457 4138
rect 490 4128 494 4131
rect 518 4101 521 4238
rect 534 4151 537 4288
rect 542 4282 545 4338
rect 614 4332 617 4338
rect 586 4328 590 4331
rect 610 4318 614 4321
rect 622 4281 625 4318
rect 630 4292 633 4358
rect 638 4342 641 4348
rect 654 4342 657 4358
rect 726 4352 729 4358
rect 698 4348 702 4351
rect 638 4282 641 4338
rect 670 4322 673 4338
rect 682 4318 686 4321
rect 694 4311 697 4338
rect 686 4308 697 4311
rect 622 4278 633 4281
rect 578 4268 582 4271
rect 618 4268 622 4271
rect 542 4263 545 4268
rect 542 4192 545 4259
rect 582 4242 585 4268
rect 630 4262 633 4278
rect 646 4272 649 4288
rect 662 4272 665 4278
rect 590 4252 593 4258
rect 598 4232 601 4258
rect 670 4242 673 4268
rect 678 4252 681 4308
rect 686 4292 689 4308
rect 682 4248 686 4251
rect 702 4242 705 4328
rect 710 4312 713 4338
rect 622 4202 625 4218
rect 630 4192 633 4228
rect 694 4182 697 4188
rect 558 4162 561 4168
rect 570 4158 574 4161
rect 602 4158 606 4161
rect 534 4148 545 4151
rect 510 4098 521 4101
rect 470 4062 473 4098
rect 510 4072 513 4098
rect 526 4082 529 4118
rect 534 4112 537 4138
rect 534 4072 537 4108
rect 462 4042 465 4048
rect 414 3942 417 3948
rect 326 3892 329 3918
rect 358 3902 361 3938
rect 374 3892 377 3928
rect 382 3892 385 3918
rect 158 3862 161 3868
rect 118 3742 121 3748
rect 122 3728 126 3731
rect 130 3718 134 3721
rect 142 3721 145 3748
rect 158 3732 161 3858
rect 210 3838 214 3841
rect 270 3802 273 3868
rect 302 3852 305 3858
rect 238 3792 241 3798
rect 318 3792 321 3868
rect 338 3866 342 3869
rect 362 3868 366 3871
rect 398 3870 401 3938
rect 414 3872 417 3908
rect 430 3892 433 3958
rect 446 3952 449 3968
rect 462 3932 465 3948
rect 470 3942 473 4018
rect 478 3952 481 4058
rect 486 3992 489 4048
rect 526 4032 529 4059
rect 496 4003 498 4007
rect 502 4003 505 4007
rect 509 4003 512 4007
rect 506 3988 510 3991
rect 486 3942 489 3978
rect 450 3918 454 3921
rect 486 3912 489 3938
rect 510 3902 513 3948
rect 462 3872 465 3888
rect 518 3872 521 3938
rect 350 3862 353 3868
rect 374 3852 377 3858
rect 510 3842 513 3859
rect 330 3788 334 3791
rect 174 3751 177 3758
rect 142 3718 153 3721
rect 138 3678 142 3681
rect 106 3668 110 3671
rect 138 3668 142 3671
rect 130 3658 134 3661
rect 94 3552 97 3658
rect 114 3649 118 3651
rect 114 3648 121 3649
rect 126 3551 129 3558
rect 26 3528 30 3531
rect 86 3522 89 3528
rect 6 3452 9 3478
rect 26 3468 30 3471
rect 46 3462 49 3518
rect 74 3478 78 3481
rect 58 3468 62 3471
rect 30 3372 33 3418
rect 34 3358 38 3361
rect 58 3348 62 3351
rect 6 3332 9 3348
rect 26 3338 30 3341
rect 58 3338 62 3341
rect 70 3332 73 3478
rect 94 3472 97 3548
rect 126 3492 129 3528
rect 138 3478 142 3481
rect 150 3472 153 3718
rect 174 3672 177 3728
rect 254 3692 257 3738
rect 270 3722 273 3747
rect 366 3742 369 3747
rect 262 3672 265 3678
rect 286 3672 289 3738
rect 366 3672 369 3728
rect 158 3552 161 3668
rect 222 3662 225 3668
rect 326 3662 329 3668
rect 342 3662 345 3668
rect 190 3652 193 3659
rect 194 3568 198 3571
rect 222 3542 225 3658
rect 286 3562 289 3568
rect 318 3551 321 3558
rect 342 3552 345 3658
rect 374 3572 377 3658
rect 382 3592 385 3658
rect 230 3532 233 3548
rect 390 3532 393 3838
rect 496 3803 498 3807
rect 502 3803 505 3807
rect 509 3803 512 3807
rect 430 3792 433 3798
rect 502 3742 505 3768
rect 422 3692 425 3738
rect 446 3722 449 3728
rect 446 3701 449 3718
rect 446 3698 457 3701
rect 454 3682 457 3698
rect 502 3682 505 3738
rect 518 3732 521 3868
rect 534 3692 537 4028
rect 542 3932 545 4148
rect 638 4142 641 4148
rect 674 4138 678 4141
rect 558 4132 561 4138
rect 558 4032 561 4128
rect 574 4062 577 4118
rect 598 4112 601 4138
rect 606 4122 609 4138
rect 642 4128 646 4131
rect 590 4108 598 4111
rect 590 4092 593 4108
rect 598 4052 601 4058
rect 606 4042 609 4078
rect 614 4062 617 4118
rect 654 4072 657 4128
rect 670 4061 673 4118
rect 686 4112 689 4138
rect 686 4062 689 4078
rect 670 4058 681 4061
rect 630 4052 633 4058
rect 666 4048 670 4051
rect 566 3992 569 4018
rect 622 3992 625 4018
rect 630 3972 633 4048
rect 678 4042 681 4058
rect 694 3992 697 4168
rect 710 4151 713 4178
rect 718 4162 721 4259
rect 726 4152 729 4338
rect 734 4322 737 4348
rect 742 4342 745 4348
rect 758 4332 761 4358
rect 778 4348 782 4351
rect 794 4348 798 4351
rect 922 4348 926 4351
rect 766 4322 769 4338
rect 786 4328 793 4331
rect 802 4328 806 4331
rect 734 4272 737 4288
rect 750 4242 753 4318
rect 790 4292 793 4328
rect 806 4272 809 4278
rect 826 4258 830 4261
rect 810 4248 814 4251
rect 790 4232 793 4248
rect 810 4238 814 4241
rect 710 4148 721 4151
rect 702 4142 705 4148
rect 718 4142 721 4148
rect 738 4148 742 4151
rect 726 4142 729 4148
rect 774 4142 777 4148
rect 702 4092 705 4138
rect 710 4052 713 4118
rect 718 4102 721 4138
rect 718 4082 721 4088
rect 726 4072 729 4118
rect 734 4082 737 4138
rect 750 4082 753 4138
rect 750 4072 753 4078
rect 710 4042 713 4048
rect 702 4012 705 4018
rect 550 3942 553 3948
rect 598 3932 601 3938
rect 614 3932 617 3938
rect 542 3872 545 3928
rect 630 3922 633 3947
rect 702 3932 705 3988
rect 726 3932 729 4068
rect 758 4062 761 4098
rect 766 4092 769 4128
rect 782 4092 785 4218
rect 794 4158 798 4161
rect 806 4152 809 4168
rect 814 4152 817 4158
rect 802 4138 806 4141
rect 822 4132 825 4218
rect 838 4212 841 4318
rect 846 4312 849 4338
rect 846 4292 849 4308
rect 854 4281 857 4348
rect 866 4328 870 4331
rect 926 4322 929 4328
rect 934 4292 937 4358
rect 1538 4358 1542 4361
rect 942 4352 945 4358
rect 974 4342 977 4348
rect 982 4342 985 4348
rect 946 4338 950 4341
rect 958 4322 961 4328
rect 966 4292 969 4318
rect 990 4282 993 4318
rect 1000 4303 1002 4307
rect 1006 4303 1009 4307
rect 1013 4303 1016 4307
rect 846 4278 857 4281
rect 846 4272 849 4278
rect 862 4272 865 4278
rect 838 4142 841 4208
rect 818 4118 822 4121
rect 822 4082 825 4108
rect 830 4102 833 4138
rect 770 4078 774 4081
rect 798 4072 801 4078
rect 822 4072 825 4078
rect 830 4072 833 4088
rect 838 4072 841 4138
rect 846 4082 849 4268
rect 866 4258 870 4261
rect 878 4252 881 4258
rect 854 4222 857 4228
rect 886 4222 889 4268
rect 894 4262 897 4278
rect 918 4272 921 4278
rect 970 4268 974 4271
rect 906 4258 910 4261
rect 934 4252 937 4268
rect 954 4258 958 4261
rect 990 4261 993 4278
rect 986 4258 993 4261
rect 998 4252 1001 4278
rect 1038 4272 1041 4278
rect 1046 4272 1049 4278
rect 1062 4272 1065 4278
rect 1034 4258 1038 4261
rect 1046 4252 1049 4258
rect 1058 4248 1062 4251
rect 910 4222 913 4248
rect 890 4218 897 4221
rect 854 4162 857 4218
rect 870 4172 873 4188
rect 878 4172 881 4178
rect 894 4162 897 4218
rect 874 4148 878 4151
rect 854 4142 857 4148
rect 894 4142 897 4158
rect 926 4152 929 4158
rect 914 4138 918 4141
rect 830 4062 833 4068
rect 758 4052 761 4058
rect 782 4052 785 4058
rect 806 4052 809 4058
rect 846 4052 849 4068
rect 878 4061 881 4118
rect 898 4078 902 4081
rect 886 4072 889 4078
rect 906 4068 910 4071
rect 878 4058 886 4061
rect 926 4061 929 4148
rect 934 4072 937 4248
rect 942 4242 945 4248
rect 962 4238 966 4241
rect 946 4188 950 4191
rect 966 4172 969 4218
rect 1046 4182 1049 4248
rect 942 4122 945 4148
rect 958 4132 961 4168
rect 1010 4148 1014 4151
rect 958 4112 961 4128
rect 974 4122 977 4148
rect 1038 4132 1041 4178
rect 1070 4162 1073 4347
rect 1086 4332 1089 4338
rect 1134 4332 1137 4338
rect 1102 4282 1105 4318
rect 1158 4281 1161 4348
rect 1166 4311 1169 4328
rect 1166 4308 1177 4311
rect 1158 4278 1169 4281
rect 1094 4262 1097 4268
rect 1102 4262 1105 4278
rect 1114 4268 1118 4271
rect 1130 4268 1134 4271
rect 1106 4258 1118 4261
rect 1126 4252 1129 4268
rect 1138 4258 1142 4261
rect 1150 4252 1153 4278
rect 1118 4242 1121 4248
rect 1150 4242 1153 4248
rect 1082 4218 1086 4221
rect 1094 4192 1097 4198
rect 1062 4142 1065 4148
rect 1070 4142 1073 4158
rect 1078 4152 1081 4158
rect 1050 4138 1054 4141
rect 1086 4132 1089 4138
rect 1026 4128 1030 4131
rect 966 4092 969 4098
rect 982 4082 985 4088
rect 990 4082 993 4108
rect 1000 4103 1002 4107
rect 1006 4103 1009 4107
rect 1013 4103 1016 4107
rect 1022 4082 1025 4128
rect 994 4078 998 4081
rect 958 4072 961 4078
rect 974 4072 977 4078
rect 990 4062 993 4068
rect 922 4058 929 4061
rect 938 4058 942 4061
rect 862 4052 865 4058
rect 770 4048 774 4051
rect 794 4048 798 4051
rect 930 4048 934 4051
rect 846 4042 849 4048
rect 830 4031 833 4038
rect 854 4031 857 4038
rect 830 4028 857 4031
rect 734 4022 737 4028
rect 734 3941 737 3968
rect 746 3948 753 3951
rect 734 3938 745 3941
rect 558 3882 561 3898
rect 574 3892 577 3898
rect 558 3752 561 3878
rect 582 3872 585 3908
rect 630 3902 633 3918
rect 710 3892 713 3918
rect 742 3892 745 3938
rect 750 3922 753 3948
rect 766 3942 769 4028
rect 790 3952 793 3998
rect 886 3992 889 4038
rect 854 3962 857 3988
rect 894 3982 897 4048
rect 814 3952 817 3958
rect 830 3952 833 3958
rect 762 3938 766 3941
rect 610 3888 614 3891
rect 694 3882 697 3888
rect 722 3878 726 3881
rect 638 3872 641 3878
rect 686 3872 689 3878
rect 714 3868 718 3871
rect 766 3871 769 3888
rect 774 3882 777 3898
rect 790 3882 793 3948
rect 894 3942 897 3958
rect 810 3938 814 3941
rect 802 3928 806 3931
rect 802 3878 806 3881
rect 766 3868 777 3871
rect 558 3742 561 3748
rect 550 3722 553 3728
rect 542 3662 545 3668
rect 410 3548 414 3551
rect 438 3542 441 3548
rect 410 3538 414 3541
rect 446 3532 449 3558
rect 454 3552 457 3659
rect 574 3661 577 3868
rect 582 3671 585 3868
rect 630 3862 633 3868
rect 762 3858 766 3861
rect 614 3792 617 3798
rect 630 3782 633 3858
rect 710 3852 713 3858
rect 666 3848 670 3851
rect 650 3758 654 3761
rect 678 3742 681 3778
rect 774 3762 777 3868
rect 790 3862 793 3878
rect 830 3852 833 3918
rect 838 3902 841 3938
rect 850 3918 854 3921
rect 862 3901 865 3938
rect 858 3898 865 3901
rect 854 3882 857 3898
rect 870 3862 873 3918
rect 910 3882 913 4008
rect 950 3962 953 4058
rect 1006 3992 1009 4078
rect 1030 4072 1033 4118
rect 1038 4092 1041 4118
rect 1030 4002 1033 4068
rect 1062 4062 1065 4068
rect 1046 4052 1049 4058
rect 1070 4052 1073 4128
rect 1094 4072 1097 4178
rect 1110 4142 1113 4218
rect 1134 4152 1137 4188
rect 1142 4162 1145 4168
rect 1122 4148 1126 4151
rect 1086 4062 1089 4068
rect 1094 4042 1097 4068
rect 1110 4032 1113 4138
rect 1126 4122 1129 4138
rect 1134 4072 1137 4148
rect 1158 4122 1161 4268
rect 1166 4262 1169 4278
rect 1166 4192 1169 4258
rect 1038 3992 1041 4018
rect 954 3948 958 3951
rect 1050 3948 1054 3951
rect 926 3882 929 3947
rect 1038 3942 1041 3948
rect 1110 3942 1113 4018
rect 1000 3903 1002 3907
rect 1006 3903 1009 3907
rect 1013 3903 1016 3907
rect 938 3888 942 3891
rect 982 3872 985 3878
rect 914 3868 918 3871
rect 842 3858 846 3861
rect 902 3852 905 3858
rect 934 3852 937 3868
rect 950 3862 953 3868
rect 858 3848 862 3851
rect 930 3848 934 3851
rect 814 3842 817 3848
rect 874 3838 878 3841
rect 970 3818 974 3821
rect 750 3752 753 3758
rect 726 3742 729 3748
rect 758 3742 761 3748
rect 766 3742 769 3748
rect 774 3742 777 3758
rect 618 3738 622 3741
rect 590 3682 593 3688
rect 662 3682 665 3718
rect 670 3692 673 3738
rect 706 3718 710 3721
rect 726 3681 729 3738
rect 734 3722 737 3728
rect 726 3678 734 3681
rect 582 3668 593 3671
rect 574 3658 582 3661
rect 496 3603 498 3607
rect 502 3603 505 3607
rect 509 3603 512 3607
rect 486 3542 489 3568
rect 494 3542 497 3578
rect 530 3558 534 3561
rect 558 3542 561 3568
rect 566 3542 569 3548
rect 494 3532 497 3538
rect 190 3492 193 3518
rect 318 3492 321 3528
rect 378 3488 382 3491
rect 230 3482 233 3488
rect 314 3478 318 3481
rect 378 3478 382 3481
rect 78 3462 81 3468
rect 118 3462 121 3468
rect 126 3462 129 3468
rect 286 3462 289 3468
rect 218 3458 222 3461
rect 250 3458 254 3461
rect 306 3458 310 3461
rect 174 3452 177 3458
rect 318 3451 321 3468
rect 370 3458 374 3461
rect 310 3448 321 3451
rect 310 3392 313 3448
rect 110 3351 113 3358
rect 206 3351 209 3368
rect 366 3352 369 3358
rect 70 3302 73 3328
rect 110 3272 113 3328
rect 62 3262 65 3268
rect 38 3192 41 3258
rect 86 3192 89 3258
rect 98 3218 102 3221
rect 34 3168 38 3171
rect 82 3168 86 3171
rect 10 3148 14 3151
rect 34 3148 38 3151
rect 6 3132 9 3138
rect 46 3132 49 3158
rect 58 3148 62 3151
rect 82 3148 86 3151
rect 94 3132 97 3158
rect 102 3132 105 3158
rect 6 3072 9 3078
rect 38 3072 41 3078
rect 10 3058 14 3061
rect 34 3058 38 3061
rect 46 3052 49 3128
rect 54 3122 57 3128
rect 34 3038 38 3041
rect 6 2932 9 2948
rect 14 2942 17 2948
rect 46 2892 49 2947
rect 62 2942 65 3068
rect 78 3063 81 3068
rect 110 3062 113 3268
rect 126 3252 129 3259
rect 142 3152 145 3348
rect 298 3348 302 3351
rect 338 3338 342 3341
rect 370 3338 374 3341
rect 190 3332 193 3338
rect 382 3332 385 3478
rect 390 3472 393 3528
rect 178 3318 182 3321
rect 146 3148 150 3151
rect 122 3138 126 3141
rect 154 3138 158 3141
rect 174 3132 177 3298
rect 230 3292 233 3318
rect 230 3282 233 3288
rect 242 3278 246 3281
rect 254 3272 257 3328
rect 270 3322 273 3328
rect 294 3292 297 3308
rect 302 3292 305 3328
rect 318 3322 321 3328
rect 374 3322 377 3328
rect 398 3322 401 3328
rect 406 3322 409 3528
rect 414 3518 422 3521
rect 414 3482 417 3518
rect 446 3482 449 3528
rect 534 3492 537 3518
rect 474 3478 478 3481
rect 422 3472 425 3478
rect 442 3468 446 3471
rect 510 3462 513 3468
rect 518 3452 521 3458
rect 442 3448 446 3451
rect 466 3448 470 3451
rect 490 3448 494 3451
rect 502 3442 505 3448
rect 450 3438 454 3441
rect 430 3382 433 3418
rect 496 3403 498 3407
rect 502 3403 505 3407
rect 509 3403 512 3407
rect 430 3358 438 3361
rect 262 3282 265 3288
rect 338 3278 345 3281
rect 342 3272 345 3278
rect 234 3268 238 3271
rect 330 3268 334 3271
rect 286 3262 289 3268
rect 274 3258 278 3261
rect 190 3152 193 3218
rect 206 3192 209 3258
rect 214 3252 217 3258
rect 234 3248 238 3251
rect 198 3162 201 3168
rect 214 3162 217 3218
rect 242 3178 246 3181
rect 234 3168 238 3171
rect 278 3162 281 3258
rect 286 3252 289 3258
rect 294 3192 297 3248
rect 302 3192 305 3268
rect 310 3262 313 3268
rect 358 3262 361 3318
rect 382 3272 385 3288
rect 398 3272 401 3278
rect 414 3262 417 3338
rect 422 3312 425 3348
rect 430 3292 433 3358
rect 470 3332 473 3347
rect 526 3342 529 3468
rect 542 3372 545 3518
rect 558 3463 561 3478
rect 574 3472 577 3538
rect 582 3382 585 3658
rect 558 3362 561 3378
rect 566 3352 569 3358
rect 590 3351 593 3668
rect 630 3662 633 3668
rect 662 3663 665 3668
rect 662 3658 665 3659
rect 614 3632 617 3658
rect 626 3648 630 3651
rect 726 3642 729 3658
rect 774 3642 777 3659
rect 742 3572 745 3618
rect 738 3558 742 3561
rect 630 3542 633 3548
rect 646 3542 649 3548
rect 670 3532 673 3548
rect 758 3542 761 3548
rect 766 3542 769 3568
rect 774 3552 777 3628
rect 782 3552 785 3818
rect 902 3792 905 3798
rect 1022 3772 1025 3918
rect 1038 3881 1041 3938
rect 1030 3878 1041 3881
rect 790 3752 793 3758
rect 806 3692 809 3718
rect 790 3552 793 3558
rect 606 3362 609 3488
rect 662 3482 665 3528
rect 726 3512 729 3518
rect 662 3472 665 3478
rect 734 3472 737 3518
rect 750 3482 753 3488
rect 750 3463 753 3468
rect 658 3459 662 3461
rect 654 3458 662 3459
rect 750 3458 753 3459
rect 722 3438 726 3441
rect 590 3348 601 3351
rect 586 3338 590 3341
rect 438 3312 441 3318
rect 458 3278 462 3281
rect 470 3272 473 3278
rect 486 3272 489 3338
rect 598 3332 601 3348
rect 598 3322 601 3328
rect 534 3312 537 3318
rect 606 3302 609 3318
rect 622 3292 625 3418
rect 654 3362 657 3368
rect 638 3341 641 3348
rect 678 3342 681 3348
rect 634 3338 641 3341
rect 514 3278 518 3281
rect 446 3262 449 3268
rect 542 3262 545 3268
rect 370 3258 374 3261
rect 342 3242 345 3258
rect 558 3252 561 3259
rect 366 3248 374 3251
rect 366 3192 369 3248
rect 382 3192 385 3238
rect 290 3168 294 3171
rect 338 3168 342 3171
rect 354 3168 358 3171
rect 406 3162 409 3218
rect 250 3158 254 3161
rect 378 3158 382 3161
rect 194 3138 198 3141
rect 182 3132 185 3138
rect 146 3088 150 3091
rect 158 3062 161 3118
rect 174 3112 177 3128
rect 182 3092 185 3128
rect 214 3111 217 3158
rect 238 3152 241 3158
rect 246 3132 249 3158
rect 254 3132 257 3148
rect 262 3132 265 3138
rect 254 3118 262 3121
rect 214 3108 225 3111
rect 222 3082 225 3108
rect 242 3088 246 3091
rect 246 3072 249 3078
rect 174 3063 177 3068
rect 110 3052 113 3058
rect 190 3052 193 3068
rect 114 2988 118 2991
rect 150 2952 153 3028
rect 190 2992 193 3048
rect 254 2952 257 3118
rect 262 3072 265 3108
rect 270 3092 273 3158
rect 342 3152 345 3158
rect 422 3152 425 3248
rect 486 3218 494 3221
rect 486 3161 489 3218
rect 496 3203 498 3207
rect 502 3203 505 3207
rect 509 3203 512 3207
rect 486 3158 497 3161
rect 446 3152 449 3158
rect 298 3148 302 3151
rect 378 3148 382 3151
rect 278 3142 281 3148
rect 326 3132 329 3148
rect 366 3142 369 3148
rect 382 3142 385 3148
rect 314 3128 318 3131
rect 262 3052 265 3058
rect 270 3052 273 3088
rect 290 3058 294 3061
rect 282 3048 286 3051
rect 306 3038 310 3041
rect 270 2992 273 3028
rect 310 2962 313 3018
rect 142 2948 150 2951
rect 26 2878 30 2881
rect 74 2878 78 2881
rect 6 2852 9 2878
rect 62 2872 65 2878
rect 86 2872 89 2878
rect 106 2868 110 2871
rect 130 2868 134 2871
rect 142 2862 145 2948
rect 246 2942 249 2948
rect 154 2938 158 2941
rect 170 2928 174 2931
rect 162 2918 166 2921
rect 190 2882 193 2918
rect 254 2901 257 2948
rect 310 2922 313 2947
rect 318 2932 321 3108
rect 326 3082 329 3088
rect 334 3072 337 3128
rect 350 3092 353 3138
rect 398 3132 401 3148
rect 366 3092 369 3118
rect 398 3082 401 3128
rect 406 3122 409 3148
rect 422 3132 425 3138
rect 430 3132 433 3138
rect 454 3132 457 3138
rect 430 3082 433 3108
rect 438 3092 441 3108
rect 470 3082 473 3148
rect 486 3142 489 3148
rect 494 3142 497 3158
rect 526 3152 529 3218
rect 566 3152 569 3158
rect 506 3148 510 3151
rect 534 3142 537 3148
rect 582 3142 585 3258
rect 622 3242 625 3248
rect 638 3241 641 3338
rect 646 3332 649 3338
rect 694 3332 697 3378
rect 726 3351 729 3358
rect 710 3332 713 3338
rect 658 3318 665 3321
rect 654 3263 657 3298
rect 654 3258 657 3259
rect 630 3238 641 3241
rect 510 3092 513 3118
rect 390 3072 393 3078
rect 326 3052 329 3058
rect 246 2898 257 2901
rect 58 2858 62 2861
rect 138 2858 142 2861
rect 114 2849 118 2851
rect 114 2848 121 2849
rect 42 2748 46 2751
rect 6 2732 9 2738
rect 14 2731 17 2748
rect 22 2742 25 2748
rect 74 2738 78 2741
rect 14 2728 22 2731
rect 90 2728 94 2731
rect 74 2718 78 2721
rect 78 2692 81 2708
rect 14 2682 17 2688
rect 86 2682 89 2728
rect 6 2652 9 2678
rect 22 2672 25 2678
rect 42 2668 46 2671
rect 74 2668 78 2671
rect 102 2662 105 2748
rect 122 2668 126 2671
rect 134 2662 137 2748
rect 142 2742 145 2748
rect 158 2732 161 2878
rect 190 2852 193 2859
rect 142 2692 145 2718
rect 158 2682 161 2728
rect 190 2712 193 2747
rect 142 2672 145 2678
rect 74 2658 78 2661
rect 50 2558 54 2561
rect 6 2532 9 2558
rect 70 2552 73 2658
rect 134 2552 137 2658
rect 22 2542 25 2548
rect 74 2538 78 2541
rect 142 2532 145 2538
rect 158 2532 161 2678
rect 206 2672 209 2738
rect 222 2663 225 2668
rect 186 2658 190 2661
rect 246 2662 249 2898
rect 258 2888 262 2891
rect 270 2862 273 2918
rect 290 2858 294 2861
rect 274 2849 278 2851
rect 274 2848 281 2849
rect 254 2752 257 2768
rect 302 2752 305 2898
rect 318 2882 321 2928
rect 334 2892 337 3068
rect 346 3048 350 3051
rect 394 3048 398 3051
rect 430 3032 433 3058
rect 518 3052 521 3138
rect 526 3092 529 3138
rect 550 3132 553 3138
rect 582 3132 585 3138
rect 542 3122 545 3128
rect 598 3112 601 3147
rect 630 3092 633 3238
rect 662 3222 665 3318
rect 678 3262 681 3328
rect 694 3302 697 3328
rect 774 3321 777 3548
rect 806 3542 809 3658
rect 822 3642 825 3738
rect 838 3692 841 3747
rect 934 3742 937 3748
rect 870 3732 873 3738
rect 914 3728 918 3731
rect 870 3672 873 3678
rect 910 3672 913 3718
rect 966 3692 969 3748
rect 1018 3718 1022 3721
rect 1000 3703 1002 3707
rect 1006 3703 1009 3707
rect 1013 3703 1016 3707
rect 990 3682 993 3688
rect 922 3668 926 3671
rect 1030 3662 1033 3878
rect 1070 3872 1073 3878
rect 1038 3842 1041 3868
rect 1062 3751 1065 3758
rect 1070 3742 1073 3868
rect 1102 3792 1105 3858
rect 1110 3842 1113 3938
rect 1118 3782 1121 3918
rect 1126 3902 1129 4059
rect 1158 3952 1161 4058
rect 1174 4042 1177 4308
rect 1222 4272 1225 4347
rect 1318 4342 1321 4347
rect 1270 4282 1273 4328
rect 1286 4292 1289 4338
rect 1254 4272 1257 4278
rect 1318 4272 1321 4328
rect 1386 4318 1390 4321
rect 1414 4272 1417 4328
rect 1422 4282 1425 4348
rect 1498 4338 1502 4341
rect 1510 4322 1513 4338
rect 1478 4272 1481 4278
rect 1234 4268 1238 4271
rect 1498 4268 1502 4271
rect 1182 4252 1185 4268
rect 1202 4258 1206 4261
rect 1182 4132 1185 4248
rect 1206 4242 1209 4248
rect 1214 4202 1217 4268
rect 1222 4222 1225 4258
rect 1238 4212 1241 4258
rect 1246 4232 1249 4268
rect 1270 4262 1273 4268
rect 1254 4242 1257 4248
rect 1278 4232 1281 4258
rect 1286 4172 1289 4178
rect 1262 4162 1265 4168
rect 1334 4162 1337 4168
rect 1238 4152 1241 4158
rect 1318 4152 1321 4158
rect 1206 4142 1209 4147
rect 1194 4088 1198 4091
rect 1222 4082 1225 4138
rect 1246 4132 1249 4138
rect 1262 4102 1265 4138
rect 1270 4092 1273 4138
rect 1278 4092 1281 4148
rect 1302 4132 1305 4138
rect 1318 4132 1321 4138
rect 1286 4092 1289 4098
rect 1302 4082 1305 4128
rect 1326 4122 1329 4128
rect 1222 3991 1225 4059
rect 1218 3988 1225 3991
rect 1230 3972 1233 4068
rect 1306 4058 1310 4061
rect 1298 4038 1302 4041
rect 1306 4028 1310 4031
rect 1318 3992 1321 4048
rect 1154 3948 1158 3951
rect 1266 3948 1270 3951
rect 1182 3922 1185 3947
rect 1294 3942 1297 3948
rect 1310 3912 1313 3918
rect 1150 3882 1153 3888
rect 1190 3872 1193 3878
rect 1162 3868 1166 3871
rect 1214 3862 1217 3868
rect 1222 3862 1225 3908
rect 1270 3882 1273 3888
rect 1326 3881 1329 4088
rect 1334 3991 1337 4018
rect 1342 3991 1345 4268
rect 1510 4262 1513 4268
rect 1350 4252 1353 4259
rect 1406 4252 1409 4259
rect 1474 4238 1478 4241
rect 1518 4222 1521 4348
rect 1566 4332 1569 4338
rect 1582 4332 1585 4378
rect 1914 4368 1918 4371
rect 3138 4368 3145 4371
rect 1702 4352 1705 4358
rect 1726 4352 1729 4368
rect 3014 4362 3017 4368
rect 1738 4358 1742 4361
rect 1770 4358 1774 4361
rect 2154 4358 2158 4361
rect 2186 4358 2190 4361
rect 2242 4358 2246 4361
rect 2338 4358 2342 4361
rect 2418 4358 2422 4361
rect 2458 4358 2462 4361
rect 2674 4358 2678 4361
rect 2698 4358 2702 4361
rect 2970 4358 2974 4361
rect 1678 4348 1686 4351
rect 1738 4348 1742 4351
rect 1520 4203 1522 4207
rect 1526 4203 1529 4207
rect 1533 4203 1536 4207
rect 1494 4162 1497 4168
rect 1442 4158 1446 4161
rect 1398 4142 1401 4147
rect 1462 4138 1470 4141
rect 1414 4112 1417 4138
rect 1430 4132 1433 4138
rect 1438 4132 1441 4138
rect 1414 4072 1417 4088
rect 1390 4022 1393 4068
rect 1414 4062 1417 4068
rect 1398 4012 1401 4058
rect 1334 3988 1345 3991
rect 1342 3952 1345 3988
rect 1410 3958 1414 3961
rect 1374 3951 1377 3958
rect 1406 3932 1409 3948
rect 1322 3878 1329 3881
rect 1258 3868 1262 3871
rect 1170 3858 1177 3861
rect 1174 3792 1177 3858
rect 1182 3842 1185 3848
rect 1130 3788 1134 3791
rect 1134 3752 1137 3778
rect 1190 3752 1193 3858
rect 1206 3852 1209 3858
rect 1198 3792 1201 3848
rect 1214 3752 1217 3858
rect 1226 3848 1230 3851
rect 1270 3802 1273 3868
rect 1142 3742 1145 3748
rect 1166 3742 1169 3748
rect 1190 3742 1193 3748
rect 1214 3742 1217 3748
rect 1046 3682 1049 3738
rect 1110 3692 1113 3698
rect 1046 3672 1049 3678
rect 1142 3672 1145 3678
rect 914 3658 918 3661
rect 978 3658 982 3661
rect 842 3648 846 3651
rect 854 3641 857 3658
rect 846 3638 857 3641
rect 846 3552 849 3638
rect 862 3632 865 3658
rect 1054 3652 1057 3658
rect 1150 3652 1153 3718
rect 1158 3712 1161 3738
rect 1158 3682 1161 3698
rect 1182 3692 1185 3728
rect 1198 3722 1201 3738
rect 1262 3722 1265 3748
rect 1278 3742 1281 3858
rect 1286 3762 1289 3868
rect 1310 3862 1313 3878
rect 1330 3868 1334 3871
rect 1326 3862 1329 3868
rect 1382 3862 1385 3868
rect 1294 3772 1297 3858
rect 1374 3842 1377 3858
rect 1406 3852 1409 3858
rect 1422 3842 1425 4058
rect 1430 3992 1433 4108
rect 1462 4072 1465 4138
rect 1470 4132 1473 4138
rect 1518 4132 1521 4138
rect 1566 4132 1569 4328
rect 1614 4272 1617 4328
rect 1574 4262 1577 4268
rect 1590 4262 1593 4268
rect 1606 4242 1609 4259
rect 1622 4151 1625 4158
rect 1486 4102 1489 4128
rect 1550 4092 1553 4098
rect 1518 4072 1521 4078
rect 1498 4068 1502 4071
rect 1522 4068 1526 4071
rect 1542 4062 1545 4088
rect 1614 4082 1617 4138
rect 1638 4102 1641 4348
rect 1678 4262 1681 4348
rect 1758 4342 1761 4348
rect 1882 4347 1886 4350
rect 1694 4292 1697 4318
rect 1710 4271 1713 4338
rect 1766 4332 1769 4338
rect 1798 4332 1801 4338
rect 1726 4291 1729 4328
rect 1722 4288 1729 4291
rect 1846 4282 1849 4288
rect 1706 4268 1713 4271
rect 1662 4192 1665 4228
rect 1678 4222 1681 4258
rect 1702 4232 1705 4268
rect 1718 4261 1721 4278
rect 1714 4258 1721 4261
rect 1750 4262 1753 4268
rect 1782 4242 1785 4259
rect 1794 4188 1798 4191
rect 1702 4158 1710 4161
rect 1674 4148 1678 4151
rect 1642 4088 1646 4091
rect 1490 4058 1494 4061
rect 1462 4042 1465 4058
rect 1490 4048 1494 4051
rect 1502 4042 1505 4048
rect 1486 3942 1489 4018
rect 1494 3992 1497 4038
rect 1520 4003 1522 4007
rect 1526 4003 1529 4007
rect 1533 4003 1536 4007
rect 1542 3982 1545 3998
rect 1530 3958 1534 3961
rect 1582 3952 1585 4058
rect 1614 4052 1617 4059
rect 1606 3951 1609 4018
rect 1646 3982 1649 3988
rect 1430 3901 1433 3918
rect 1430 3898 1441 3901
rect 1438 3882 1441 3898
rect 1346 3838 1350 3841
rect 1326 3762 1329 3768
rect 1358 3762 1361 3818
rect 1390 3772 1393 3818
rect 1438 3802 1441 3859
rect 1466 3858 1470 3861
rect 1170 3688 1174 3691
rect 1214 3672 1217 3718
rect 1210 3668 1214 3671
rect 1230 3663 1233 3708
rect 1286 3682 1289 3758
rect 1294 3722 1297 3747
rect 1310 3692 1313 3728
rect 1302 3682 1305 3688
rect 1286 3672 1289 3678
rect 1350 3672 1353 3748
rect 1358 3742 1361 3758
rect 1398 3752 1401 3778
rect 1406 3742 1409 3748
rect 1430 3742 1433 3768
rect 1438 3752 1441 3768
rect 1446 3742 1449 3758
rect 1470 3742 1473 3758
rect 1478 3752 1481 3778
rect 1486 3762 1489 3938
rect 1502 3912 1505 3928
rect 1510 3922 1513 3928
rect 1542 3912 1545 3918
rect 1502 3892 1505 3898
rect 1526 3882 1529 3888
rect 1590 3863 1593 3878
rect 1606 3872 1609 3928
rect 1622 3872 1625 3888
rect 1562 3858 1566 3861
rect 1520 3803 1522 3807
rect 1526 3803 1529 3807
rect 1533 3803 1536 3807
rect 1506 3768 1510 3771
rect 1546 3748 1550 3751
rect 1378 3738 1382 3741
rect 1362 3728 1366 3731
rect 1354 3668 1358 3671
rect 1246 3662 1249 3668
rect 1122 3648 1126 3651
rect 886 3552 889 3568
rect 990 3542 993 3618
rect 1242 3588 1246 3591
rect 1142 3562 1145 3568
rect 1174 3551 1177 3558
rect 1262 3552 1265 3648
rect 1374 3642 1377 3659
rect 1406 3592 1409 3648
rect 1414 3592 1417 3738
rect 1422 3732 1425 3738
rect 1454 3692 1457 3698
rect 1446 3672 1449 3678
rect 1470 3672 1473 3738
rect 1498 3728 1502 3731
rect 1478 3722 1481 3728
rect 1434 3668 1438 3671
rect 1518 3663 1521 3698
rect 1386 3558 1390 3561
rect 1438 3552 1441 3618
rect 1520 3603 1522 3607
rect 1526 3603 1529 3607
rect 1533 3603 1536 3607
rect 1082 3547 1086 3550
rect 1250 3548 1254 3551
rect 1394 3548 1398 3551
rect 1350 3542 1353 3547
rect 1446 3542 1449 3548
rect 1514 3547 1518 3550
rect 1534 3542 1537 3548
rect 1558 3542 1561 3758
rect 1574 3742 1577 3747
rect 1606 3742 1609 3758
rect 1654 3692 1657 4098
rect 1662 4072 1665 4118
rect 1686 4112 1689 4138
rect 1694 4122 1697 4148
rect 1702 4102 1705 4158
rect 1722 4148 1726 4151
rect 1710 4142 1713 4148
rect 1742 4141 1745 4158
rect 1750 4152 1753 4158
rect 1774 4142 1777 4148
rect 1742 4138 1750 4141
rect 1718 4112 1721 4138
rect 1742 4122 1745 4128
rect 1742 4092 1745 4098
rect 1678 4062 1681 4078
rect 1710 4063 1713 4068
rect 1758 4062 1761 4128
rect 1782 4082 1785 4138
rect 1790 4112 1793 4178
rect 1806 4172 1809 4238
rect 1814 4222 1817 4268
rect 1822 4262 1825 4268
rect 1886 4262 1889 4328
rect 1882 4258 1886 4261
rect 1830 4248 1838 4251
rect 1814 4182 1817 4218
rect 1822 4212 1825 4218
rect 1830 4201 1833 4248
rect 1822 4198 1833 4201
rect 1822 4192 1825 4198
rect 1838 4172 1841 4198
rect 1806 4162 1809 4168
rect 1894 4152 1897 4228
rect 1902 4172 1905 4348
rect 1966 4332 1969 4338
rect 1910 4263 1913 4288
rect 1982 4282 1985 4347
rect 1950 4272 1953 4278
rect 1942 4192 1945 4248
rect 1966 4222 1969 4268
rect 2002 4258 2006 4261
rect 1974 4192 1977 4248
rect 1994 4238 1998 4241
rect 2014 4222 2017 4348
rect 2078 4332 2081 4338
rect 2024 4303 2026 4307
rect 2030 4303 2033 4307
rect 2037 4303 2040 4307
rect 2078 4302 2081 4328
rect 2094 4311 2097 4347
rect 2134 4332 2137 4338
rect 2094 4308 2105 4311
rect 2102 4292 2105 4308
rect 2126 4301 2129 4328
rect 2118 4298 2129 4301
rect 2118 4292 2121 4298
rect 2082 4288 2086 4291
rect 2022 4282 2025 4288
rect 2094 4282 2097 4288
rect 2034 4268 2038 4271
rect 2134 4262 2137 4298
rect 2010 4218 2014 4221
rect 1926 4172 1929 4178
rect 1850 4148 1854 4151
rect 1822 4142 1825 4148
rect 1862 4142 1865 4148
rect 1886 4142 1889 4148
rect 1766 4072 1769 4078
rect 1774 4072 1777 4078
rect 1790 4072 1793 4108
rect 1814 4082 1817 4138
rect 1810 4068 1814 4071
rect 1790 4062 1793 4068
rect 1838 4062 1841 4138
rect 1846 4072 1849 4078
rect 1870 4072 1873 4138
rect 1886 4072 1889 4138
rect 1854 4062 1857 4068
rect 1662 3952 1665 3968
rect 1678 3942 1681 4058
rect 1742 4052 1745 4058
rect 1822 4022 1825 4038
rect 1782 3992 1785 4008
rect 1762 3988 1766 3991
rect 1818 3988 1822 3991
rect 1694 3932 1697 3947
rect 1766 3912 1769 3958
rect 1782 3952 1785 3958
rect 1786 3938 1790 3941
rect 1798 3931 1801 3958
rect 1814 3952 1817 3958
rect 1862 3942 1865 4058
rect 1870 3992 1873 4068
rect 1878 4052 1881 4058
rect 1902 3962 1905 4168
rect 1942 4152 1945 4158
rect 1910 4142 1913 4148
rect 1910 3991 1913 4058
rect 1918 4002 1921 4058
rect 1926 4022 1929 4148
rect 1962 4138 1966 4141
rect 1970 4128 1974 4131
rect 1986 4128 1993 4131
rect 1950 4052 1953 4118
rect 1962 4058 1966 4061
rect 1934 4042 1937 4048
rect 1954 4038 1958 4041
rect 1910 3988 1921 3991
rect 1918 3952 1921 3988
rect 1926 3962 1929 4018
rect 1966 3962 1969 4018
rect 1974 3972 1977 4048
rect 1982 4012 1985 4118
rect 1990 4082 1993 4128
rect 1998 4082 2001 4208
rect 2010 4168 2014 4171
rect 2022 4152 2025 4248
rect 2078 4232 2081 4248
rect 2030 4192 2033 4208
rect 2038 4161 2041 4218
rect 2050 4168 2054 4171
rect 2038 4158 2049 4161
rect 2010 4148 2014 4151
rect 2024 4103 2026 4107
rect 2030 4103 2033 4107
rect 2037 4103 2040 4107
rect 1990 3992 1993 4078
rect 2010 4058 2014 4061
rect 2002 4038 2006 4041
rect 2014 3962 2017 4018
rect 1982 3952 1985 3958
rect 1790 3928 1801 3931
rect 1818 3938 1822 3941
rect 1842 3938 1846 3941
rect 1734 3892 1737 3908
rect 1790 3892 1793 3928
rect 1718 3872 1721 3878
rect 1726 3872 1729 3878
rect 1662 3792 1665 3858
rect 1686 3852 1689 3859
rect 1734 3791 1737 3838
rect 1726 3788 1737 3791
rect 1694 3782 1697 3788
rect 1682 3758 1686 3761
rect 1674 3748 1678 3751
rect 1678 3732 1681 3738
rect 1726 3702 1729 3788
rect 1750 3752 1753 3838
rect 1746 3748 1750 3751
rect 1742 3672 1745 3748
rect 1758 3742 1761 3868
rect 1774 3852 1777 3858
rect 1790 3852 1793 3858
rect 1806 3792 1809 3938
rect 1834 3928 1838 3931
rect 1830 3842 1833 3858
rect 1854 3852 1857 3938
rect 1862 3882 1865 3938
rect 1886 3932 1889 3948
rect 1894 3942 1897 3948
rect 1874 3928 1878 3931
rect 1862 3852 1865 3859
rect 1770 3747 1774 3750
rect 1806 3742 1809 3788
rect 1854 3772 1857 3848
rect 1878 3792 1881 3918
rect 1902 3872 1905 3938
rect 1910 3862 1913 3868
rect 1814 3732 1817 3748
rect 1830 3722 1833 3728
rect 1838 3712 1841 3758
rect 1854 3752 1857 3768
rect 1870 3742 1873 3788
rect 1878 3752 1881 3758
rect 1858 3738 1862 3741
rect 1754 3688 1758 3691
rect 1806 3672 1809 3698
rect 1838 3692 1841 3708
rect 1854 3692 1857 3728
rect 1878 3672 1881 3738
rect 1894 3732 1897 3848
rect 1918 3812 1921 3948
rect 1926 3792 1929 3868
rect 1934 3862 1937 3918
rect 1950 3862 1953 3928
rect 1958 3882 1961 3928
rect 1974 3882 1977 3928
rect 1950 3842 1953 3858
rect 1974 3832 1977 3878
rect 1982 3832 1985 3918
rect 1990 3852 1993 3958
rect 2046 3952 2049 4158
rect 2066 4148 2070 4151
rect 2086 4142 2089 4218
rect 2102 4202 2105 4218
rect 2094 4152 2097 4178
rect 2110 4152 2113 4158
rect 2082 4128 2086 4131
rect 2054 4072 2057 4078
rect 2062 4072 2065 4118
rect 2066 4058 2070 4061
rect 2082 4048 2086 4051
rect 2094 3972 2097 4148
rect 2118 4141 2121 4218
rect 2138 4188 2142 4191
rect 2110 4138 2121 4141
rect 2110 4062 2113 4138
rect 2122 4128 2126 4131
rect 2142 4122 2145 4128
rect 2118 4052 2121 4078
rect 2150 4052 2153 4358
rect 2162 4348 2166 4351
rect 2166 4342 2169 4348
rect 2174 4332 2177 4338
rect 2214 4332 2217 4338
rect 2202 4328 2206 4331
rect 2166 4252 2169 4259
rect 2182 4242 2185 4318
rect 2206 4261 2209 4318
rect 2230 4272 2233 4278
rect 2198 4258 2209 4261
rect 2166 4152 2169 4228
rect 2182 4172 2185 4198
rect 2178 4168 2182 4171
rect 2162 4148 2166 4151
rect 2198 4141 2201 4258
rect 2206 4242 2209 4248
rect 2214 4231 2217 4258
rect 2206 4228 2217 4231
rect 2206 4212 2209 4228
rect 2214 4212 2217 4218
rect 2206 4162 2209 4168
rect 2218 4158 2222 4161
rect 2222 4142 2225 4148
rect 2198 4138 2206 4141
rect 2186 4128 2190 4131
rect 2178 4118 2182 4121
rect 2222 4112 2225 4118
rect 2230 4082 2233 4248
rect 2238 4182 2241 4328
rect 2246 4242 2249 4318
rect 2254 4292 2257 4348
rect 2286 4322 2289 4348
rect 2302 4342 2305 4348
rect 2310 4332 2313 4348
rect 2406 4322 2409 4328
rect 2286 4271 2289 4318
rect 2326 4272 2329 4318
rect 2286 4268 2294 4271
rect 2350 4271 2353 4318
rect 2414 4291 2417 4358
rect 2526 4352 2529 4358
rect 2606 4352 2609 4358
rect 2990 4352 2993 4358
rect 3142 4352 3145 4368
rect 3174 4368 3182 4371
rect 3198 4368 3206 4371
rect 3498 4368 3502 4371
rect 3174 4352 3177 4368
rect 3198 4352 3201 4368
rect 3438 4362 3441 4368
rect 3478 4362 3481 4368
rect 3558 4362 3561 4428
rect 3568 4403 3570 4407
rect 3574 4403 3577 4407
rect 3581 4403 3584 4407
rect 3686 4402 3689 4428
rect 3750 4402 3753 4428
rect 3598 4362 3601 4368
rect 3622 4362 3625 4368
rect 3306 4358 3310 4361
rect 3338 4358 3342 4361
rect 3418 4358 3422 4361
rect 2826 4348 2830 4351
rect 2422 4342 2425 4348
rect 2650 4338 2654 4341
rect 2682 4338 2686 4341
rect 2722 4338 2726 4341
rect 2414 4288 2425 4291
rect 2350 4268 2361 4271
rect 2322 4258 2326 4261
rect 2254 4232 2257 4258
rect 2274 4248 2278 4251
rect 2250 4218 2254 4221
rect 2262 4202 2265 4238
rect 2286 4232 2289 4258
rect 2302 4252 2305 4258
rect 2350 4252 2353 4258
rect 2314 4238 2318 4241
rect 2294 4202 2297 4238
rect 2326 4202 2329 4218
rect 2334 4192 2337 4208
rect 2246 4182 2249 4188
rect 2278 4162 2281 4188
rect 2326 4172 2329 4178
rect 2310 4132 2313 4138
rect 2258 4128 2262 4131
rect 2246 4082 2249 4128
rect 2182 4052 2185 4078
rect 2190 4062 2193 4068
rect 2254 4052 2257 4078
rect 2262 4062 2265 4118
rect 2270 4112 2273 4118
rect 2114 4048 2118 4051
rect 2130 4048 2134 4051
rect 2210 4048 2214 4051
rect 2106 4038 2110 4041
rect 2138 4038 2142 4041
rect 2110 4012 2113 4018
rect 2126 3962 2129 4018
rect 2150 3972 2153 4048
rect 2202 4038 2206 4041
rect 2226 4038 2230 4041
rect 2278 4041 2281 4118
rect 2302 4092 2305 4098
rect 2274 4038 2281 4041
rect 2150 3962 2153 3968
rect 2094 3952 2097 3958
rect 2002 3948 2006 3951
rect 2134 3942 2137 3948
rect 1998 3882 2001 3908
rect 2014 3892 2017 3918
rect 2024 3903 2026 3907
rect 2030 3903 2033 3907
rect 2037 3903 2040 3907
rect 1998 3862 2001 3878
rect 2026 3868 2030 3871
rect 2002 3838 2006 3841
rect 1902 3752 1905 3758
rect 1918 3752 1921 3768
rect 1926 3752 1929 3788
rect 1886 3682 1889 3688
rect 1802 3668 1806 3671
rect 1726 3663 1729 3668
rect 1590 3652 1593 3659
rect 1918 3662 1921 3748
rect 1934 3742 1937 3818
rect 1958 3792 1961 3828
rect 1966 3772 1969 3818
rect 1978 3758 1982 3761
rect 1950 3742 1953 3748
rect 1990 3742 1993 3748
rect 1934 3712 1937 3728
rect 1934 3682 1937 3698
rect 1934 3672 1937 3678
rect 1982 3672 1985 3738
rect 1622 3592 1625 3658
rect 1822 3652 1825 3659
rect 1882 3658 1886 3661
rect 1982 3662 1985 3668
rect 1990 3662 1993 3698
rect 2006 3692 2009 3758
rect 2014 3752 2017 3868
rect 2046 3842 2049 3858
rect 2058 3848 2062 3851
rect 2054 3802 2057 3818
rect 2070 3762 2073 3938
rect 2078 3932 2081 3938
rect 2090 3928 2094 3931
rect 2086 3862 2089 3878
rect 2106 3868 2110 3871
rect 2118 3862 2121 3878
rect 2126 3862 2129 3918
rect 2150 3902 2153 3918
rect 2150 3862 2153 3868
rect 2082 3838 2086 3841
rect 2094 3801 2097 3848
rect 2114 3838 2118 3841
rect 2126 3812 2129 3848
rect 2142 3842 2145 3858
rect 2158 3852 2161 3938
rect 2174 3932 2177 4018
rect 2190 3962 2193 4018
rect 2206 3962 2209 4018
rect 2214 3952 2217 3978
rect 2278 3962 2281 4018
rect 2242 3958 2246 3961
rect 2186 3948 2190 3951
rect 2190 3932 2193 3938
rect 2174 3862 2177 3868
rect 2182 3862 2185 3878
rect 2170 3838 2174 3841
rect 2154 3818 2161 3821
rect 2094 3798 2105 3801
rect 2102 3782 2105 3798
rect 2150 3792 2153 3808
rect 2158 3792 2161 3818
rect 2190 3792 2193 3848
rect 2206 3842 2209 3918
rect 2230 3912 2233 3918
rect 2214 3862 2217 3868
rect 2246 3862 2249 3868
rect 2254 3861 2257 3918
rect 2254 3858 2265 3861
rect 2274 3858 2278 3861
rect 2218 3848 2222 3851
rect 2250 3848 2254 3851
rect 2262 3842 2265 3858
rect 2234 3838 2238 3841
rect 2286 3832 2289 4058
rect 2326 4052 2329 4168
rect 2334 4152 2337 4158
rect 2342 4082 2345 4248
rect 2358 4242 2361 4268
rect 2414 4262 2417 4278
rect 2374 4252 2377 4258
rect 2350 4152 2353 4218
rect 2382 4192 2385 4238
rect 2390 4232 2393 4258
rect 2394 4178 2398 4181
rect 2402 4158 2406 4161
rect 2366 4132 2369 4138
rect 2350 4102 2353 4128
rect 2358 4122 2361 4128
rect 2398 4112 2401 4138
rect 2334 4072 2337 4078
rect 2338 4058 2342 4061
rect 2350 4052 2353 4098
rect 2382 4082 2385 4098
rect 2358 4062 2361 4068
rect 2402 4058 2406 4061
rect 2414 4052 2417 4228
rect 2422 4162 2425 4288
rect 2438 4282 2441 4288
rect 2446 4262 2449 4338
rect 2598 4332 2601 4338
rect 2662 4332 2665 4338
rect 2758 4331 2761 4348
rect 2782 4331 2785 4348
rect 2946 4338 2950 4341
rect 2886 4332 2889 4338
rect 2974 4332 2977 4338
rect 2990 4332 2993 4348
rect 2674 4318 2678 4321
rect 2462 4302 2465 4318
rect 2454 4282 2457 4288
rect 2498 4278 2502 4281
rect 2478 4262 2481 4268
rect 2438 4252 2441 4258
rect 2446 4181 2449 4258
rect 2518 4252 2521 4318
rect 2526 4262 2529 4268
rect 2454 4242 2457 4248
rect 2542 4242 2545 4318
rect 2614 4271 2617 4318
rect 2702 4292 2705 4318
rect 2710 4312 2713 4328
rect 2754 4328 2761 4331
rect 2778 4328 2785 4331
rect 2814 4322 2817 4328
rect 2722 4278 2726 4281
rect 2614 4268 2625 4271
rect 2562 4258 2574 4261
rect 2594 4248 2598 4251
rect 2574 4242 2577 4248
rect 2530 4238 2534 4241
rect 2602 4238 2606 4241
rect 2486 4232 2489 4238
rect 2614 4232 2617 4258
rect 2622 4242 2625 4268
rect 2638 4262 2641 4268
rect 2686 4262 2689 4268
rect 2766 4262 2769 4268
rect 2666 4258 2670 4261
rect 2706 4258 2710 4261
rect 2670 4252 2673 4258
rect 2750 4252 2753 4258
rect 2658 4248 2662 4251
rect 2494 4222 2497 4228
rect 2544 4203 2546 4207
rect 2550 4203 2553 4207
rect 2557 4203 2560 4207
rect 2438 4178 2449 4181
rect 2430 4162 2433 4168
rect 2438 4152 2441 4178
rect 2450 4168 2454 4171
rect 2462 4162 2465 4188
rect 2502 4172 2505 4178
rect 2482 4168 2486 4171
rect 2530 4158 2534 4161
rect 2486 4152 2489 4158
rect 2466 4148 2470 4151
rect 2506 4148 2510 4151
rect 2422 4112 2425 4118
rect 2446 4072 2449 4078
rect 2454 4062 2457 4118
rect 2466 4078 2470 4081
rect 2442 4058 2446 4061
rect 2426 4048 2430 4051
rect 2326 4042 2329 4048
rect 2294 3862 2297 4028
rect 2334 3992 2337 4048
rect 2414 4042 2417 4048
rect 2370 4038 2374 4041
rect 2434 4038 2438 4041
rect 2478 4041 2481 4108
rect 2490 4058 2494 4061
rect 2502 4052 2505 4108
rect 2478 4038 2486 4041
rect 2346 3968 2350 3971
rect 2318 3962 2321 3968
rect 2358 3952 2361 4038
rect 2326 3932 2329 3938
rect 2342 3932 2345 3938
rect 2374 3932 2377 4018
rect 2470 3992 2473 4018
rect 2422 3952 2425 3978
rect 2454 3952 2457 3978
rect 2386 3948 2390 3951
rect 2494 3932 2497 4018
rect 2378 3918 2382 3921
rect 2122 3788 2126 3791
rect 2130 3778 2134 3781
rect 1858 3638 1862 3641
rect 1658 3618 1662 3621
rect 1886 3592 1889 3628
rect 1918 3582 1921 3588
rect 1942 3572 1945 3648
rect 1950 3642 1953 3659
rect 1746 3568 1750 3571
rect 1626 3548 1630 3551
rect 970 3538 974 3541
rect 1034 3538 1038 3541
rect 782 3422 785 3538
rect 806 3492 809 3538
rect 830 3482 833 3488
rect 894 3472 897 3538
rect 1062 3532 1065 3538
rect 1158 3532 1161 3538
rect 1000 3503 1002 3507
rect 1006 3503 1009 3507
rect 1013 3503 1016 3507
rect 1026 3488 1030 3491
rect 942 3472 945 3478
rect 1078 3472 1081 3528
rect 1138 3488 1142 3491
rect 1198 3472 1201 3538
rect 818 3428 822 3431
rect 790 3352 793 3368
rect 822 3351 825 3418
rect 774 3318 785 3321
rect 726 3282 729 3318
rect 678 3142 681 3258
rect 714 3238 718 3241
rect 726 3212 729 3278
rect 750 3262 753 3288
rect 774 3282 777 3308
rect 758 3232 761 3238
rect 694 3151 697 3178
rect 766 3172 769 3218
rect 678 3132 681 3138
rect 666 3118 670 3121
rect 762 3118 766 3121
rect 690 3078 694 3081
rect 578 3068 582 3071
rect 594 3058 598 3061
rect 490 3048 494 3051
rect 594 3048 598 3051
rect 622 3042 625 3058
rect 630 3052 633 3068
rect 610 3038 622 3041
rect 496 3003 498 3007
rect 502 3003 505 3007
rect 509 3003 512 3007
rect 374 2992 377 2998
rect 518 2991 521 2998
rect 510 2988 521 2991
rect 342 2952 345 2968
rect 406 2951 409 2958
rect 438 2952 441 2968
rect 494 2962 497 2978
rect 462 2892 465 2908
rect 334 2882 337 2888
rect 438 2872 441 2888
rect 366 2852 369 2859
rect 350 2762 353 2768
rect 390 2742 393 2858
rect 430 2842 433 2848
rect 438 2842 441 2868
rect 398 2752 401 2838
rect 446 2832 449 2838
rect 470 2792 473 2918
rect 478 2902 481 2938
rect 510 2892 513 2988
rect 526 2972 529 3018
rect 598 2981 601 3018
rect 590 2978 601 2981
rect 590 2972 593 2978
rect 602 2968 606 2971
rect 534 2962 537 2968
rect 546 2958 550 2961
rect 574 2948 582 2951
rect 534 2902 537 2948
rect 534 2882 537 2898
rect 542 2882 545 2938
rect 566 2932 569 2938
rect 566 2912 569 2928
rect 542 2872 545 2878
rect 550 2872 553 2898
rect 574 2892 577 2948
rect 622 2942 625 3038
rect 630 2952 633 3048
rect 646 3002 649 3068
rect 654 2982 657 3058
rect 662 3052 665 3078
rect 702 3072 705 3098
rect 774 3092 777 3278
rect 782 3262 785 3318
rect 790 3252 793 3258
rect 798 3252 801 3308
rect 830 3291 833 3438
rect 846 3352 849 3468
rect 894 3462 897 3468
rect 870 3432 873 3458
rect 926 3442 929 3448
rect 942 3352 945 3468
rect 1198 3462 1201 3468
rect 1206 3463 1209 3518
rect 1246 3492 1249 3538
rect 1270 3532 1273 3538
rect 1270 3472 1273 3528
rect 1334 3472 1337 3538
rect 1382 3532 1385 3538
rect 958 3452 961 3459
rect 1070 3392 1073 3459
rect 1238 3441 1241 3458
rect 1230 3438 1241 3441
rect 1146 3418 1150 3421
rect 1098 3388 1102 3391
rect 926 3342 929 3348
rect 942 3342 945 3348
rect 822 3288 833 3291
rect 822 3272 825 3288
rect 854 3282 857 3338
rect 886 3322 889 3338
rect 1014 3332 1017 3338
rect 1030 3322 1033 3347
rect 986 3318 990 3321
rect 1000 3303 1002 3307
rect 1006 3303 1009 3307
rect 1013 3303 1016 3307
rect 1038 3291 1041 3388
rect 1190 3352 1193 3368
rect 1198 3352 1201 3418
rect 1138 3348 1142 3351
rect 1206 3342 1209 3378
rect 1222 3362 1225 3368
rect 1230 3352 1233 3438
rect 1246 3392 1249 3468
rect 1254 3452 1257 3458
rect 1270 3382 1273 3468
rect 1310 3462 1313 3468
rect 1342 3463 1345 3478
rect 1398 3462 1401 3468
rect 1294 3352 1297 3438
rect 1330 3358 1334 3361
rect 1034 3288 1041 3291
rect 1062 3282 1065 3338
rect 1110 3332 1113 3338
rect 1222 3322 1225 3338
rect 1230 3332 1233 3348
rect 1266 3348 1270 3351
rect 1358 3342 1361 3458
rect 1378 3448 1382 3451
rect 1406 3391 1409 3538
rect 1422 3532 1425 3538
rect 1414 3482 1417 3488
rect 1438 3482 1441 3528
rect 1446 3472 1449 3528
rect 1398 3388 1409 3391
rect 1322 3318 1326 3321
rect 1126 3292 1129 3308
rect 810 3268 814 3271
rect 854 3263 857 3268
rect 854 3258 857 3259
rect 1190 3262 1193 3268
rect 786 3228 790 3231
rect 790 3151 793 3218
rect 798 3152 801 3248
rect 770 3078 774 3081
rect 702 3052 705 3058
rect 714 3048 718 3051
rect 674 3038 678 3041
rect 638 2952 641 2978
rect 670 2952 673 2958
rect 678 2952 681 2978
rect 602 2928 606 2931
rect 614 2922 617 2928
rect 582 2892 585 2908
rect 630 2902 633 2948
rect 594 2888 598 2891
rect 582 2872 585 2888
rect 614 2882 617 2898
rect 638 2892 641 2948
rect 662 2942 665 2948
rect 702 2942 705 2988
rect 726 2982 729 3068
rect 758 3062 761 3068
rect 774 3062 777 3068
rect 750 3052 753 3058
rect 782 3052 785 3108
rect 790 3062 793 3128
rect 814 3112 817 3258
rect 830 3072 833 3098
rect 770 3048 774 3051
rect 746 3018 750 3021
rect 710 2952 713 2958
rect 682 2938 686 2941
rect 646 2882 649 2938
rect 654 2892 657 2918
rect 662 2892 665 2928
rect 686 2912 689 2938
rect 718 2932 721 2948
rect 734 2942 737 2948
rect 670 2882 673 2908
rect 694 2902 697 2918
rect 478 2862 481 2868
rect 494 2852 497 2868
rect 550 2862 553 2868
rect 590 2862 593 2878
rect 522 2858 526 2861
rect 494 2842 497 2848
rect 542 2822 545 2828
rect 496 2803 498 2807
rect 502 2803 505 2807
rect 509 2803 512 2807
rect 466 2758 470 2761
rect 550 2752 553 2858
rect 558 2842 561 2858
rect 574 2832 577 2848
rect 598 2832 601 2878
rect 662 2862 665 2868
rect 634 2858 654 2861
rect 686 2852 689 2888
rect 702 2862 705 2918
rect 742 2882 745 2988
rect 750 2942 753 2958
rect 694 2842 697 2858
rect 710 2851 713 2868
rect 702 2848 713 2851
rect 590 2752 593 2818
rect 302 2672 305 2738
rect 398 2672 401 2738
rect 254 2662 257 2668
rect 302 2662 305 2668
rect 350 2662 353 2668
rect 398 2662 401 2668
rect 414 2663 417 2688
rect 190 2551 193 2558
rect 26 2528 30 2531
rect 42 2528 46 2531
rect 78 2482 81 2528
rect 74 2478 78 2481
rect 6 2452 9 2478
rect 26 2468 30 2471
rect 58 2468 62 2471
rect 58 2458 62 2461
rect 34 2449 38 2451
rect 34 2448 41 2449
rect 46 2382 49 2388
rect 110 2382 113 2468
rect 142 2462 145 2518
rect 158 2482 161 2528
rect 190 2472 193 2528
rect 246 2502 249 2658
rect 318 2652 321 2659
rect 486 2662 489 2718
rect 502 2682 505 2738
rect 558 2672 561 2728
rect 582 2682 585 2688
rect 366 2622 369 2648
rect 290 2618 294 2621
rect 286 2542 289 2548
rect 294 2522 297 2548
rect 258 2518 262 2521
rect 270 2482 273 2518
rect 118 2452 121 2458
rect 6 2332 9 2338
rect 14 2332 17 2338
rect 22 2332 25 2358
rect 30 2342 33 2348
rect 94 2282 97 2378
rect 174 2372 177 2418
rect 190 2382 193 2468
rect 206 2463 209 2468
rect 274 2428 278 2431
rect 142 2352 145 2358
rect 118 2312 121 2338
rect 150 2332 153 2338
rect 158 2321 161 2348
rect 154 2318 161 2321
rect 174 2282 177 2328
rect 126 2272 129 2278
rect 146 2268 150 2271
rect 178 2268 182 2271
rect 166 2262 169 2268
rect 190 2262 193 2358
rect 206 2352 209 2358
rect 262 2342 265 2378
rect 270 2342 273 2348
rect 210 2338 214 2341
rect 210 2328 214 2331
rect 218 2318 222 2321
rect 318 2312 321 2538
rect 366 2531 369 2618
rect 382 2572 385 2618
rect 398 2542 401 2658
rect 542 2652 545 2658
rect 482 2638 486 2641
rect 490 2618 494 2621
rect 542 2612 545 2648
rect 496 2603 498 2607
rect 502 2603 505 2607
rect 509 2603 512 2607
rect 558 2552 561 2668
rect 574 2661 577 2678
rect 570 2658 577 2661
rect 590 2662 593 2748
rect 598 2742 601 2828
rect 634 2818 638 2821
rect 614 2762 617 2768
rect 626 2758 630 2761
rect 686 2752 689 2818
rect 694 2762 697 2768
rect 634 2748 638 2751
rect 650 2748 654 2751
rect 614 2742 617 2748
rect 622 2742 625 2748
rect 598 2692 601 2738
rect 654 2732 657 2738
rect 670 2722 673 2738
rect 598 2672 601 2688
rect 626 2678 630 2681
rect 642 2678 646 2681
rect 654 2672 657 2688
rect 566 2642 569 2658
rect 606 2651 609 2658
rect 602 2648 609 2651
rect 614 2642 617 2668
rect 622 2652 625 2658
rect 646 2652 649 2658
rect 506 2548 510 2551
rect 422 2542 425 2548
rect 378 2538 382 2541
rect 398 2532 401 2538
rect 366 2528 377 2531
rect 338 2478 342 2481
rect 326 2462 329 2468
rect 342 2442 345 2458
rect 342 2392 345 2438
rect 326 2352 329 2368
rect 342 2362 345 2388
rect 358 2352 361 2498
rect 374 2482 377 2528
rect 406 2382 409 2468
rect 414 2452 417 2458
rect 358 2292 361 2348
rect 390 2342 393 2378
rect 462 2352 465 2548
rect 490 2528 494 2531
rect 470 2522 473 2528
rect 482 2518 486 2521
rect 470 2511 473 2518
rect 470 2508 481 2511
rect 478 2482 481 2508
rect 478 2462 481 2468
rect 478 2392 481 2448
rect 398 2322 401 2348
rect 454 2322 457 2328
rect 306 2288 310 2291
rect 330 2288 334 2291
rect 234 2278 238 2281
rect 6 2242 9 2248
rect 54 2192 57 2208
rect 78 2192 81 2228
rect 94 2192 97 2259
rect 34 2188 38 2191
rect 6 2172 9 2178
rect 22 2152 25 2178
rect 198 2172 201 2278
rect 230 2252 233 2259
rect 302 2252 305 2278
rect 350 2272 353 2278
rect 322 2268 326 2271
rect 342 2262 345 2268
rect 358 2262 361 2288
rect 454 2272 457 2308
rect 382 2262 385 2268
rect 298 2228 302 2231
rect 322 2178 326 2181
rect 114 2168 118 2171
rect 70 2152 73 2168
rect 118 2162 121 2168
rect 238 2151 241 2158
rect 30 2072 33 2078
rect 6 2042 9 2048
rect 22 2042 25 2058
rect 46 2002 49 2148
rect 94 1992 97 2148
rect 102 2132 105 2138
rect 110 2132 113 2148
rect 182 2142 185 2147
rect 182 2072 185 2128
rect 294 2111 297 2148
rect 310 2132 313 2158
rect 318 2142 321 2148
rect 306 2118 310 2121
rect 294 2108 305 2111
rect 302 2092 305 2108
rect 290 2078 294 2081
rect 118 2012 121 2059
rect 30 1972 33 1978
rect 54 1962 57 1968
rect 22 1952 25 1958
rect 118 1951 121 1958
rect 6 1942 9 1948
rect 46 1922 49 1948
rect 134 1942 137 2068
rect 214 2063 217 2068
rect 146 2038 150 2041
rect 150 1992 153 1998
rect 6 1872 9 1878
rect 22 1862 25 1888
rect 134 1872 137 1938
rect 30 1852 33 1868
rect 134 1862 137 1868
rect 150 1862 153 1868
rect 34 1788 38 1791
rect 6 1772 9 1778
rect 54 1762 57 1768
rect 50 1748 54 1751
rect 22 1692 25 1748
rect 70 1742 73 1748
rect 106 1747 110 1750
rect 30 1672 33 1678
rect 46 1662 49 1668
rect 54 1662 57 1688
rect 86 1662 89 1738
rect 118 1702 121 1859
rect 166 1792 169 2028
rect 214 1951 217 1968
rect 230 1942 233 2068
rect 246 2042 249 2078
rect 254 2042 257 2048
rect 254 1952 257 1978
rect 206 1792 209 1938
rect 214 1872 217 1878
rect 230 1872 233 1938
rect 246 1932 249 1938
rect 262 1912 265 2078
rect 310 2072 313 2078
rect 282 2068 286 2071
rect 270 2062 273 2068
rect 318 2062 321 2068
rect 326 2062 329 2118
rect 342 2092 345 2258
rect 334 2062 337 2088
rect 342 2062 345 2068
rect 290 2058 294 2061
rect 310 1992 313 2058
rect 358 2052 361 2068
rect 366 2062 369 2168
rect 382 2152 385 2158
rect 390 2142 393 2258
rect 430 2152 433 2168
rect 446 2152 449 2158
rect 462 2152 465 2348
rect 470 2272 473 2278
rect 470 2152 473 2228
rect 478 2172 481 2318
rect 486 2262 489 2508
rect 526 2492 529 2538
rect 550 2482 553 2528
rect 510 2442 513 2458
rect 518 2452 521 2478
rect 496 2403 498 2407
rect 502 2403 505 2407
rect 509 2403 512 2407
rect 558 2392 561 2518
rect 582 2502 585 2547
rect 598 2532 601 2538
rect 614 2532 617 2638
rect 654 2602 657 2668
rect 670 2662 673 2718
rect 686 2682 689 2748
rect 702 2732 705 2848
rect 742 2842 745 2859
rect 710 2752 713 2758
rect 758 2752 761 3018
rect 782 3002 785 3048
rect 790 2992 793 3058
rect 798 2982 801 3068
rect 782 2952 785 2978
rect 822 2952 825 2978
rect 794 2948 798 2951
rect 830 2942 833 3068
rect 838 3032 841 3248
rect 958 3242 961 3258
rect 958 3232 961 3238
rect 918 3202 921 3218
rect 982 3192 985 3258
rect 1014 3182 1017 3188
rect 1014 3152 1017 3178
rect 854 3112 857 3118
rect 862 3062 865 3068
rect 794 2938 798 2941
rect 766 2762 769 2918
rect 774 2912 777 2938
rect 806 2872 809 2918
rect 814 2912 817 2938
rect 810 2858 814 2861
rect 838 2852 841 2858
rect 846 2832 849 3058
rect 886 2892 889 3118
rect 894 3092 897 3148
rect 906 3138 913 3141
rect 910 3072 913 3138
rect 1026 3138 1030 3141
rect 950 3122 953 3128
rect 910 3062 913 3068
rect 934 3062 937 3108
rect 958 3102 961 3138
rect 1000 3103 1002 3107
rect 1006 3103 1009 3107
rect 1013 3103 1016 3107
rect 910 2952 913 3058
rect 926 2951 929 2968
rect 894 2942 897 2948
rect 910 2942 913 2948
rect 934 2922 937 3058
rect 990 3042 993 3048
rect 982 2892 985 2958
rect 990 2952 993 2968
rect 998 2942 1001 3088
rect 1022 3062 1025 3068
rect 1014 2972 1017 3028
rect 866 2878 870 2881
rect 886 2872 889 2888
rect 918 2872 921 2878
rect 810 2828 814 2831
rect 814 2812 817 2818
rect 854 2762 857 2868
rect 910 2862 913 2868
rect 950 2862 953 2878
rect 958 2872 961 2878
rect 882 2858 886 2861
rect 878 2852 881 2858
rect 894 2792 897 2858
rect 942 2842 945 2848
rect 950 2802 953 2858
rect 970 2848 974 2851
rect 990 2792 993 2938
rect 1000 2903 1002 2907
rect 1006 2903 1009 2907
rect 1013 2903 1016 2907
rect 1022 2882 1025 3058
rect 1038 2942 1041 3208
rect 1046 3042 1049 3058
rect 1062 2902 1065 3259
rect 1158 3212 1161 3259
rect 1118 3192 1121 3208
rect 1102 3182 1105 3188
rect 1206 3171 1209 3318
rect 1226 3288 1230 3291
rect 1198 3168 1209 3171
rect 1238 3262 1241 3268
rect 1262 3262 1265 3268
rect 1150 3152 1153 3158
rect 1102 3082 1105 3088
rect 1150 3072 1153 3148
rect 1082 2958 1086 2961
rect 1070 2952 1073 2958
rect 1070 2932 1073 2938
rect 1082 2928 1086 2931
rect 1034 2858 1038 2861
rect 818 2758 822 2761
rect 830 2752 833 2758
rect 842 2748 846 2751
rect 866 2748 870 2751
rect 1022 2751 1025 2758
rect 910 2742 913 2747
rect 866 2738 870 2741
rect 930 2738 934 2741
rect 718 2732 721 2738
rect 694 2712 697 2718
rect 718 2712 721 2728
rect 702 2672 705 2698
rect 722 2678 726 2681
rect 734 2672 737 2738
rect 818 2718 822 2721
rect 846 2712 849 2738
rect 878 2712 881 2738
rect 742 2672 745 2708
rect 770 2668 774 2671
rect 670 2652 673 2658
rect 662 2571 665 2618
rect 654 2568 665 2571
rect 686 2572 689 2668
rect 706 2658 710 2661
rect 730 2658 734 2661
rect 694 2642 697 2658
rect 702 2582 705 2658
rect 714 2648 718 2651
rect 654 2562 657 2568
rect 638 2552 641 2558
rect 654 2552 657 2558
rect 630 2542 633 2548
rect 570 2478 574 2481
rect 578 2468 582 2471
rect 614 2452 617 2478
rect 622 2472 625 2518
rect 638 2512 641 2548
rect 686 2532 689 2547
rect 650 2528 654 2531
rect 638 2492 641 2498
rect 694 2482 697 2538
rect 698 2459 702 2461
rect 694 2458 702 2459
rect 510 2322 513 2348
rect 510 2302 513 2318
rect 422 2142 425 2148
rect 390 2102 393 2138
rect 438 2072 441 2078
rect 394 2068 398 2071
rect 406 2068 414 2071
rect 346 2038 350 2041
rect 274 1958 278 1961
rect 294 1942 297 1978
rect 318 1972 321 2038
rect 330 1958 334 1961
rect 314 1948 318 1951
rect 274 1938 278 1941
rect 302 1932 305 1948
rect 302 1891 305 1928
rect 302 1888 310 1891
rect 326 1882 329 1888
rect 230 1862 233 1868
rect 250 1859 254 1862
rect 222 1742 225 1838
rect 334 1832 337 1918
rect 342 1882 345 1988
rect 366 1982 369 2058
rect 382 2052 385 2058
rect 398 1972 401 1978
rect 374 1962 377 1968
rect 382 1942 385 1958
rect 398 1952 401 1958
rect 342 1842 345 1878
rect 350 1862 353 1868
rect 358 1862 361 1938
rect 362 1858 366 1861
rect 374 1852 377 1918
rect 382 1872 385 1908
rect 382 1842 385 1858
rect 398 1852 401 1948
rect 406 1942 409 2068
rect 414 1992 417 1998
rect 422 1962 425 2058
rect 446 2052 449 2118
rect 454 1952 457 2098
rect 462 2052 465 2148
rect 470 2062 473 2088
rect 474 2058 478 2061
rect 466 2038 470 2041
rect 486 2022 489 2258
rect 534 2232 537 2338
rect 574 2332 577 2348
rect 582 2342 585 2368
rect 582 2282 585 2338
rect 542 2252 545 2258
rect 542 2242 545 2248
rect 496 2203 498 2207
rect 502 2203 505 2207
rect 509 2203 512 2207
rect 518 2182 521 2218
rect 542 2152 545 2238
rect 558 2142 561 2278
rect 598 2192 601 2418
rect 606 2332 609 2448
rect 630 2442 633 2458
rect 614 2352 617 2438
rect 654 2352 657 2448
rect 710 2352 713 2568
rect 718 2381 721 2548
rect 742 2522 745 2668
rect 814 2662 817 2678
rect 838 2662 841 2678
rect 754 2658 758 2661
rect 766 2652 769 2658
rect 750 2642 753 2648
rect 754 2588 758 2591
rect 758 2552 761 2558
rect 766 2552 769 2648
rect 790 2552 793 2578
rect 726 2462 729 2468
rect 718 2378 729 2381
rect 718 2352 721 2368
rect 726 2362 729 2378
rect 742 2352 745 2508
rect 758 2502 761 2548
rect 798 2542 801 2598
rect 818 2558 830 2561
rect 846 2552 849 2558
rect 842 2548 846 2551
rect 822 2542 825 2548
rect 854 2542 857 2708
rect 874 2688 878 2691
rect 886 2672 889 2678
rect 902 2663 905 2668
rect 934 2662 937 2738
rect 902 2658 905 2659
rect 966 2642 969 2648
rect 862 2552 865 2578
rect 874 2548 878 2551
rect 786 2538 790 2541
rect 758 2482 761 2488
rect 798 2482 801 2538
rect 770 2458 774 2461
rect 778 2458 785 2461
rect 650 2348 654 2351
rect 714 2348 718 2351
rect 678 2342 681 2348
rect 606 2301 609 2318
rect 606 2298 617 2301
rect 614 2263 617 2298
rect 686 2282 689 2348
rect 738 2338 742 2341
rect 646 2262 649 2278
rect 706 2268 710 2271
rect 738 2268 742 2271
rect 726 2262 729 2268
rect 686 2252 689 2258
rect 734 2242 737 2258
rect 574 2162 577 2168
rect 570 2158 574 2161
rect 606 2151 609 2178
rect 678 2152 681 2188
rect 726 2142 729 2147
rect 514 2138 518 2141
rect 534 2132 537 2138
rect 558 2102 561 2138
rect 542 2072 545 2098
rect 522 2058 526 2061
rect 494 2052 497 2058
rect 494 2032 497 2048
rect 526 2042 529 2048
rect 506 2038 510 2041
rect 406 1882 409 1938
rect 446 1872 449 1878
rect 470 1862 473 2018
rect 496 2003 498 2007
rect 502 2003 505 2007
rect 509 2003 512 2007
rect 518 1952 521 2018
rect 558 1992 561 2059
rect 530 1968 534 1971
rect 554 1958 558 1961
rect 574 1961 577 2118
rect 590 2082 593 2138
rect 678 2132 681 2138
rect 750 2132 753 2278
rect 758 2212 761 2418
rect 782 2342 785 2458
rect 798 2342 801 2347
rect 814 2332 817 2538
rect 834 2518 838 2521
rect 862 2492 865 2548
rect 886 2542 889 2608
rect 902 2552 905 2558
rect 926 2552 929 2558
rect 914 2548 918 2551
rect 874 2538 881 2541
rect 766 2321 769 2328
rect 766 2318 777 2321
rect 774 2162 777 2318
rect 798 2282 801 2328
rect 830 2312 833 2468
rect 838 2462 841 2488
rect 846 2472 849 2478
rect 862 2432 865 2468
rect 870 2462 873 2528
rect 878 2482 881 2538
rect 886 2492 889 2538
rect 894 2532 897 2548
rect 922 2538 926 2541
rect 886 2472 889 2478
rect 894 2468 902 2471
rect 878 2462 881 2468
rect 894 2452 897 2468
rect 910 2462 913 2528
rect 918 2472 921 2478
rect 942 2472 945 2538
rect 958 2522 961 2547
rect 974 2482 977 2718
rect 1000 2703 1002 2707
rect 1006 2703 1009 2707
rect 1013 2703 1016 2707
rect 1030 2672 1033 2738
rect 1078 2692 1081 2908
rect 1086 2892 1089 2898
rect 1098 2888 1102 2891
rect 1126 2792 1129 2948
rect 1134 2872 1137 2938
rect 1142 2892 1145 3058
rect 1166 2992 1169 3148
rect 1198 3092 1201 3168
rect 1238 3132 1241 3258
rect 1250 3148 1254 3151
rect 1238 3072 1241 3128
rect 1230 3002 1233 3059
rect 1182 2992 1185 2998
rect 1278 2992 1281 2998
rect 1286 2992 1289 3278
rect 1334 3262 1337 3268
rect 1310 3218 1318 3221
rect 1310 3152 1313 3218
rect 1358 3192 1361 3328
rect 1398 3292 1401 3388
rect 1414 3352 1417 3358
rect 1422 3332 1425 3458
rect 1430 3282 1433 3468
rect 1438 3452 1441 3458
rect 1446 3392 1449 3468
rect 1454 3462 1457 3518
rect 1506 3488 1510 3491
rect 1574 3482 1577 3548
rect 1646 3532 1649 3568
rect 1862 3552 1865 3558
rect 1686 3542 1689 3548
rect 1478 3462 1481 3468
rect 1494 3462 1497 3468
rect 1458 3448 1462 3451
rect 1494 3392 1497 3458
rect 1574 3452 1577 3459
rect 1602 3418 1606 3421
rect 1520 3403 1522 3407
rect 1526 3403 1529 3407
rect 1533 3403 1536 3407
rect 1542 3352 1545 3358
rect 1446 3302 1449 3347
rect 1478 3342 1481 3348
rect 1502 3322 1505 3338
rect 1526 3332 1529 3348
rect 1550 3342 1553 3388
rect 1558 3352 1561 3418
rect 1606 3352 1609 3408
rect 1586 3348 1590 3351
rect 1554 3338 1558 3341
rect 1566 3332 1569 3348
rect 1594 3338 1598 3341
rect 1494 3292 1497 3318
rect 1574 3312 1577 3338
rect 1422 3262 1425 3278
rect 1438 3272 1441 3288
rect 1518 3282 1521 3288
rect 1478 3272 1481 3278
rect 1486 3272 1489 3278
rect 1506 3268 1510 3271
rect 1370 3258 1374 3261
rect 1442 3258 1446 3261
rect 1466 3258 1470 3261
rect 1426 3248 1430 3251
rect 1334 3162 1337 3168
rect 1374 3152 1377 3248
rect 1406 3152 1409 3228
rect 1414 3212 1417 3218
rect 1414 3162 1417 3168
rect 1438 3152 1441 3238
rect 1462 3182 1465 3248
rect 1520 3203 1522 3207
rect 1526 3203 1529 3207
rect 1533 3203 1536 3207
rect 1478 3152 1481 3198
rect 1550 3192 1553 3258
rect 1550 3172 1553 3178
rect 1574 3152 1577 3208
rect 1582 3192 1585 3259
rect 1606 3218 1614 3221
rect 1606 3212 1609 3218
rect 1622 3211 1625 3508
rect 1638 3472 1641 3518
rect 1654 3512 1657 3518
rect 1686 3472 1689 3538
rect 1718 3532 1721 3547
rect 1782 3542 1785 3548
rect 1814 3542 1817 3547
rect 1882 3538 1886 3541
rect 1766 3463 1769 3478
rect 1782 3472 1785 3538
rect 1862 3532 1865 3538
rect 1902 3531 1905 3558
rect 1918 3552 1921 3558
rect 1914 3538 1918 3541
rect 1902 3528 1913 3531
rect 1846 3522 1849 3528
rect 1910 3492 1913 3528
rect 1942 3512 1945 3568
rect 1794 3488 1798 3491
rect 1898 3478 1902 3481
rect 1934 3472 1937 3478
rect 1898 3468 1902 3471
rect 1670 3452 1673 3459
rect 1942 3462 1945 3488
rect 1702 3412 1705 3418
rect 1634 3358 1638 3361
rect 1662 3352 1665 3358
rect 1670 3352 1673 3358
rect 1694 3352 1697 3368
rect 1802 3358 1806 3361
rect 1630 3232 1633 3348
rect 1690 3338 1694 3341
rect 1662 3292 1665 3338
rect 1678 3263 1681 3318
rect 1702 3312 1705 3318
rect 1650 3258 1654 3261
rect 1734 3262 1737 3348
rect 1762 3347 1766 3350
rect 1782 3342 1785 3348
rect 1822 3292 1825 3298
rect 1830 3292 1833 3458
rect 1862 3402 1865 3459
rect 1926 3442 1929 3458
rect 1950 3451 1953 3498
rect 1942 3448 1953 3451
rect 1958 3492 1961 3548
rect 1966 3542 1969 3658
rect 1982 3592 1985 3648
rect 2006 3642 2009 3648
rect 2014 3592 2017 3748
rect 2054 3742 2057 3747
rect 2024 3703 2026 3707
rect 2030 3703 2033 3707
rect 2037 3703 2040 3707
rect 2026 3688 2030 3691
rect 2078 3682 2081 3748
rect 2078 3672 2081 3678
rect 2086 3661 2089 3698
rect 2078 3658 2089 3661
rect 2022 3592 2025 3648
rect 1978 3548 1982 3551
rect 1978 3538 1982 3541
rect 1998 3532 2001 3558
rect 1974 3492 1977 3528
rect 2006 3502 2009 3558
rect 2022 3552 2025 3558
rect 2070 3552 2073 3588
rect 2058 3548 2062 3551
rect 2034 3538 2038 3541
rect 2042 3528 2046 3531
rect 1958 3472 1961 3488
rect 1998 3472 2001 3478
rect 1910 3412 1913 3438
rect 1910 3372 1913 3378
rect 1846 3342 1849 3348
rect 1806 3272 1809 3288
rect 1714 3238 1718 3241
rect 1630 3221 1633 3228
rect 1630 3218 1641 3221
rect 1614 3208 1625 3211
rect 1598 3152 1601 3158
rect 1614 3152 1617 3208
rect 1630 3172 1633 3178
rect 1586 3148 1590 3151
rect 1318 3122 1321 3138
rect 1334 3132 1337 3138
rect 1310 3118 1318 3121
rect 1294 3092 1297 3098
rect 1302 3062 1305 3118
rect 1310 3072 1313 3118
rect 1374 3081 1377 3148
rect 1366 3078 1377 3081
rect 1390 3081 1393 3118
rect 1390 3078 1401 3081
rect 1326 3072 1329 3078
rect 1350 3062 1353 3068
rect 1366 3062 1369 3078
rect 1398 3072 1401 3078
rect 1386 3068 1390 3071
rect 1374 3062 1377 3068
rect 1406 3062 1409 3128
rect 1438 3092 1441 3138
rect 1510 3132 1513 3148
rect 1486 3092 1489 3108
rect 1438 3072 1441 3088
rect 1454 3072 1457 3078
rect 1486 3072 1489 3088
rect 1326 3042 1329 3048
rect 1166 2912 1169 2988
rect 1366 2982 1369 3058
rect 1374 2971 1377 3058
rect 1458 3048 1462 3051
rect 1414 3042 1417 3048
rect 1382 3032 1385 3038
rect 1494 3002 1497 3118
rect 1518 3082 1521 3088
rect 1374 2968 1385 2971
rect 1382 2952 1385 2968
rect 1414 2952 1417 2968
rect 1422 2952 1425 2958
rect 1226 2948 1230 2951
rect 1222 2872 1225 2938
rect 1278 2892 1281 2908
rect 1342 2882 1345 2938
rect 1350 2902 1353 2947
rect 1398 2942 1401 2948
rect 1446 2942 1449 2998
rect 1466 2968 1470 2971
rect 1382 2912 1385 2938
rect 1406 2932 1409 2938
rect 1446 2902 1449 2938
rect 1382 2892 1385 2898
rect 1462 2892 1465 2928
rect 1370 2888 1374 2891
rect 1490 2888 1494 2891
rect 1294 2872 1297 2878
rect 1462 2872 1465 2878
rect 1158 2852 1161 2859
rect 1186 2788 1190 2791
rect 1122 2748 1126 2751
rect 1102 2732 1105 2738
rect 1086 2712 1089 2718
rect 1018 2659 1022 2661
rect 1014 2658 1022 2659
rect 1022 2592 1025 2598
rect 990 2542 993 2548
rect 1030 2542 1033 2668
rect 1118 2662 1121 2708
rect 1214 2692 1217 2859
rect 1222 2742 1225 2868
rect 1178 2688 1182 2691
rect 1222 2672 1225 2738
rect 1142 2662 1145 2668
rect 1222 2662 1225 2668
rect 1078 2562 1081 2618
rect 1074 2548 1078 2551
rect 1102 2542 1105 2548
rect 1118 2522 1121 2658
rect 1214 2642 1217 2658
rect 1222 2592 1225 2658
rect 1138 2568 1142 2571
rect 1146 2548 1150 2551
rect 1000 2503 1002 2507
rect 1006 2503 1009 2507
rect 1013 2503 1016 2507
rect 982 2482 985 2488
rect 1034 2478 1038 2481
rect 1010 2468 1014 2471
rect 930 2458 934 2461
rect 982 2452 985 2468
rect 1046 2462 1049 2488
rect 1102 2482 1105 2488
rect 1146 2478 1150 2481
rect 1070 2462 1073 2468
rect 906 2448 918 2451
rect 974 2422 977 2448
rect 866 2418 870 2421
rect 866 2388 870 2391
rect 922 2358 926 2361
rect 898 2348 902 2351
rect 926 2342 929 2348
rect 934 2332 937 2368
rect 966 2352 969 2378
rect 954 2348 958 2351
rect 866 2328 870 2331
rect 954 2328 958 2331
rect 982 2331 985 2438
rect 1078 2432 1081 2478
rect 1086 2472 1089 2478
rect 1094 2442 1097 2478
rect 1110 2472 1113 2478
rect 1122 2468 1126 2471
rect 1182 2463 1185 2468
rect 1122 2458 1126 2461
rect 1146 2458 1150 2461
rect 1182 2458 1185 2459
rect 998 2402 1001 2418
rect 990 2362 993 2368
rect 998 2362 1001 2378
rect 998 2352 1001 2358
rect 1014 2352 1017 2358
rect 1010 2338 1014 2341
rect 982 2328 990 2331
rect 878 2322 881 2328
rect 886 2302 889 2328
rect 942 2322 945 2328
rect 974 2322 977 2328
rect 886 2282 889 2298
rect 962 2288 966 2291
rect 982 2282 985 2318
rect 1000 2303 1002 2307
rect 1006 2303 1009 2307
rect 1013 2303 1016 2307
rect 1030 2282 1033 2418
rect 1062 2362 1065 2418
rect 1062 2342 1065 2347
rect 1078 2322 1081 2428
rect 1126 2392 1129 2428
rect 1158 2351 1161 2368
rect 1190 2352 1193 2468
rect 1094 2342 1097 2348
rect 1190 2342 1193 2348
rect 1086 2282 1089 2288
rect 1102 2282 1105 2288
rect 994 2278 998 2281
rect 798 2272 801 2278
rect 894 2272 897 2278
rect 878 2262 881 2268
rect 790 2252 793 2259
rect 790 2162 793 2168
rect 794 2148 798 2151
rect 690 2128 694 2131
rect 686 2112 689 2118
rect 590 2072 593 2078
rect 662 2072 665 2098
rect 694 2072 697 2078
rect 726 2072 729 2128
rect 750 2102 753 2128
rect 774 2092 777 2098
rect 798 2092 801 2148
rect 782 2082 785 2088
rect 814 2072 817 2078
rect 674 2068 678 2071
rect 622 2042 625 2048
rect 638 2022 641 2058
rect 654 2052 657 2058
rect 678 2032 681 2048
rect 710 2042 713 2059
rect 810 2058 814 2061
rect 822 2052 825 2178
rect 878 2162 881 2218
rect 830 2142 833 2158
rect 870 2152 873 2158
rect 902 2152 905 2278
rect 958 2272 961 2278
rect 922 2268 926 2271
rect 950 2242 953 2258
rect 910 2152 913 2238
rect 966 2182 969 2228
rect 874 2148 878 2151
rect 838 2142 841 2148
rect 846 2142 849 2148
rect 830 2132 833 2138
rect 966 2132 969 2178
rect 974 2132 977 2278
rect 1142 2272 1145 2338
rect 1206 2312 1209 2538
rect 1230 2392 1233 2858
rect 1238 2722 1241 2748
rect 1226 2388 1230 2391
rect 1206 2272 1209 2308
rect 1026 2268 1030 2271
rect 1038 2242 1041 2258
rect 1070 2252 1073 2258
rect 1134 2252 1137 2259
rect 1202 2238 1206 2241
rect 990 2142 993 2218
rect 998 2152 1001 2238
rect 1078 2202 1081 2218
rect 1062 2192 1065 2198
rect 1086 2142 1089 2148
rect 1094 2142 1097 2218
rect 1158 2162 1161 2168
rect 1146 2158 1150 2161
rect 1210 2158 1214 2161
rect 1110 2152 1113 2158
rect 1138 2148 1142 2151
rect 914 2128 918 2131
rect 994 2128 998 2131
rect 918 2092 921 2118
rect 982 2092 985 2118
rect 1000 2103 1002 2107
rect 1006 2103 1009 2107
rect 1013 2103 1016 2107
rect 1038 2092 1041 2138
rect 1094 2132 1097 2138
rect 1134 2132 1137 2138
rect 1114 2128 1118 2131
rect 850 2088 854 2091
rect 1078 2082 1081 2088
rect 970 2078 974 2081
rect 1010 2078 1014 2081
rect 1050 2078 1054 2081
rect 1098 2078 1102 2081
rect 910 2072 913 2078
rect 834 2068 838 2071
rect 986 2068 993 2071
rect 1034 2068 1038 2071
rect 886 2062 889 2068
rect 990 2062 993 2068
rect 1046 2062 1049 2068
rect 1070 2062 1073 2078
rect 1026 2058 1030 2061
rect 786 2038 790 2041
rect 802 2038 806 2041
rect 638 1992 641 2018
rect 606 1962 609 1978
rect 650 1968 654 1971
rect 630 1962 633 1968
rect 574 1958 582 1961
rect 614 1952 617 1958
rect 662 1952 665 1958
rect 538 1948 542 1951
rect 586 1948 590 1951
rect 478 1942 481 1947
rect 510 1942 513 1948
rect 566 1942 569 1948
rect 554 1938 558 1941
rect 586 1938 590 1941
rect 246 1752 249 1758
rect 254 1752 257 1758
rect 302 1752 305 1788
rect 310 1762 313 1828
rect 318 1772 321 1818
rect 334 1772 337 1818
rect 350 1792 353 1828
rect 390 1782 393 1818
rect 254 1742 257 1748
rect 234 1738 238 1741
rect 198 1682 201 1732
rect 198 1672 201 1678
rect 154 1668 158 1671
rect 26 1658 30 1661
rect 6 1642 9 1648
rect 6 1542 9 1548
rect 22 1542 25 1548
rect 22 1518 30 1521
rect 22 1462 25 1518
rect 62 1492 65 1548
rect 86 1542 89 1658
rect 118 1652 121 1659
rect 194 1658 198 1661
rect 166 1652 169 1658
rect 178 1638 182 1641
rect 94 1551 97 1628
rect 126 1572 129 1578
rect 30 1472 33 1478
rect 122 1468 126 1471
rect 6 1442 9 1448
rect 34 1378 38 1381
rect 22 1352 25 1368
rect 46 1362 49 1458
rect 62 1412 65 1418
rect 54 1382 57 1388
rect 70 1352 73 1398
rect 150 1392 153 1548
rect 166 1492 169 1618
rect 178 1548 182 1551
rect 182 1482 185 1528
rect 190 1522 193 1608
rect 206 1542 209 1688
rect 238 1682 241 1718
rect 226 1678 230 1681
rect 214 1672 217 1678
rect 214 1552 217 1618
rect 230 1582 233 1678
rect 246 1671 249 1738
rect 262 1732 265 1738
rect 278 1732 281 1748
rect 366 1742 369 1758
rect 374 1752 377 1768
rect 314 1738 318 1741
rect 286 1722 289 1738
rect 238 1668 249 1671
rect 238 1642 241 1668
rect 246 1642 249 1658
rect 238 1612 241 1638
rect 246 1592 249 1618
rect 254 1592 257 1718
rect 282 1688 286 1691
rect 274 1678 278 1681
rect 270 1662 273 1678
rect 286 1672 289 1678
rect 302 1662 305 1678
rect 286 1642 289 1658
rect 310 1652 313 1728
rect 310 1642 313 1648
rect 230 1562 233 1568
rect 206 1502 209 1538
rect 222 1492 225 1518
rect 206 1482 209 1488
rect 222 1482 225 1488
rect 158 1452 161 1458
rect 166 1391 169 1478
rect 230 1462 233 1488
rect 238 1472 241 1558
rect 246 1512 249 1588
rect 254 1552 257 1578
rect 294 1562 297 1608
rect 266 1548 270 1551
rect 298 1548 302 1551
rect 254 1492 257 1548
rect 274 1538 281 1541
rect 262 1492 265 1538
rect 158 1388 169 1391
rect 82 1368 86 1371
rect 50 1348 54 1351
rect 142 1351 145 1378
rect 6 1342 9 1348
rect 22 1262 25 1298
rect 30 1272 33 1278
rect 134 1272 137 1338
rect 158 1292 161 1388
rect 190 1362 193 1388
rect 174 1342 177 1358
rect 190 1282 193 1318
rect 198 1292 201 1358
rect 206 1352 209 1458
rect 270 1452 273 1508
rect 278 1492 281 1538
rect 306 1478 310 1481
rect 282 1468 286 1471
rect 318 1462 321 1708
rect 366 1692 369 1728
rect 330 1658 334 1661
rect 330 1638 334 1641
rect 342 1631 345 1668
rect 334 1628 345 1631
rect 350 1662 353 1688
rect 382 1672 385 1678
rect 334 1552 337 1628
rect 350 1611 353 1658
rect 390 1652 393 1678
rect 406 1672 409 1858
rect 438 1852 441 1858
rect 478 1852 481 1908
rect 534 1892 537 1938
rect 550 1872 553 1918
rect 442 1838 462 1841
rect 486 1841 489 1868
rect 530 1858 534 1861
rect 478 1838 489 1841
rect 422 1792 425 1838
rect 454 1752 457 1818
rect 434 1747 438 1750
rect 478 1751 481 1838
rect 558 1832 561 1868
rect 566 1862 569 1938
rect 598 1872 601 1918
rect 614 1872 617 1878
rect 618 1868 622 1871
rect 582 1852 585 1868
rect 630 1862 633 1948
rect 638 1872 641 1938
rect 646 1862 649 1868
rect 662 1862 665 1918
rect 670 1912 673 1958
rect 678 1952 681 1958
rect 686 1892 689 1968
rect 694 1952 697 1988
rect 702 1962 705 1968
rect 758 1952 761 2038
rect 822 2012 825 2048
rect 838 2042 841 2058
rect 878 2052 881 2058
rect 982 2052 985 2058
rect 1054 2052 1057 2058
rect 970 2048 974 2051
rect 894 2042 897 2048
rect 886 2032 889 2038
rect 898 1988 902 1991
rect 934 1982 937 2018
rect 1094 1982 1097 2058
rect 794 1968 798 1971
rect 994 1968 998 1971
rect 798 1962 801 1968
rect 1110 1952 1113 2118
rect 1126 2081 1129 2118
rect 1118 2078 1129 2081
rect 1118 2031 1121 2078
rect 1134 2071 1137 2128
rect 1130 2068 1137 2071
rect 1134 2052 1137 2058
rect 1150 2052 1153 2158
rect 1182 2152 1185 2158
rect 1222 2142 1225 2358
rect 1238 2262 1241 2718
rect 1262 2572 1265 2818
rect 1310 2772 1313 2859
rect 1446 2822 1449 2859
rect 1474 2768 1478 2771
rect 1270 2692 1273 2768
rect 1278 2762 1281 2768
rect 1310 2751 1313 2758
rect 1418 2748 1422 2751
rect 1310 2672 1313 2728
rect 1374 2722 1377 2728
rect 1406 2672 1409 2728
rect 1462 2692 1465 2708
rect 1334 2662 1337 2668
rect 1382 2662 1385 2668
rect 1322 2658 1326 2661
rect 1478 2662 1481 2668
rect 1334 2621 1337 2658
rect 1398 2652 1401 2659
rect 1366 2642 1369 2648
rect 1334 2618 1345 2621
rect 1342 2592 1345 2618
rect 1262 2482 1265 2568
rect 1274 2538 1278 2541
rect 1350 2491 1353 2638
rect 1494 2602 1497 2659
rect 1446 2592 1449 2598
rect 1502 2592 1505 3068
rect 1526 3062 1529 3148
rect 1622 3142 1625 3148
rect 1538 3138 1542 3141
rect 1550 3132 1553 3138
rect 1566 3122 1569 3138
rect 1550 3072 1553 3118
rect 1546 3068 1550 3071
rect 1558 3062 1561 3098
rect 1582 3062 1585 3138
rect 1606 3122 1609 3138
rect 1614 3132 1617 3138
rect 1590 3072 1593 3108
rect 1602 3088 1606 3091
rect 1522 3058 1526 3061
rect 1542 3052 1545 3058
rect 1562 3048 1566 3051
rect 1590 3011 1593 3058
rect 1638 3052 1641 3218
rect 1694 3162 1697 3168
rect 1658 3158 1662 3161
rect 1718 3152 1721 3168
rect 1774 3152 1777 3258
rect 1790 3252 1793 3259
rect 1878 3232 1881 3347
rect 1894 3332 1897 3338
rect 1918 3332 1921 3368
rect 1926 3302 1929 3358
rect 1902 3272 1905 3288
rect 1918 3272 1921 3278
rect 1934 3272 1937 3428
rect 1942 3392 1945 3448
rect 1958 3442 1961 3468
rect 1990 3462 1993 3468
rect 2002 3458 2006 3461
rect 1974 3442 1977 3458
rect 1950 3352 1953 3438
rect 1958 3362 1961 3368
rect 1954 3338 1958 3341
rect 1926 3262 1929 3268
rect 1886 3242 1889 3259
rect 1950 3252 1953 3258
rect 1974 3202 1977 3438
rect 1990 3332 1993 3348
rect 2014 3262 2017 3518
rect 2024 3503 2026 3507
rect 2030 3503 2033 3507
rect 2037 3503 2040 3507
rect 2054 3472 2057 3538
rect 2042 3468 2046 3471
rect 2030 3462 2033 3468
rect 2070 3462 2073 3548
rect 2078 3492 2081 3658
rect 2094 3602 2097 3659
rect 2126 3652 2129 3758
rect 2158 3742 2161 3768
rect 2170 3758 2174 3761
rect 2134 3682 2137 3728
rect 2142 3712 2145 3728
rect 2154 3678 2158 3681
rect 2134 3662 2137 3668
rect 2126 3632 2129 3648
rect 2142 3642 2145 3658
rect 2162 3638 2166 3641
rect 2174 3641 2177 3718
rect 2182 3702 2185 3728
rect 2198 3672 2201 3738
rect 2214 3732 2217 3818
rect 2230 3752 2233 3818
rect 2222 3742 2225 3748
rect 2238 3682 2241 3708
rect 2198 3662 2201 3668
rect 2218 3658 2222 3661
rect 2190 3642 2193 3658
rect 2198 3652 2201 3658
rect 2206 3642 2209 3648
rect 2174 3638 2182 3641
rect 2138 3618 2142 3621
rect 2194 3618 2198 3621
rect 2110 3592 2113 3608
rect 2194 3588 2198 3591
rect 2142 3562 2145 3568
rect 2130 3558 2134 3561
rect 2158 3552 2161 3558
rect 2106 3548 2110 3551
rect 2090 3538 2094 3541
rect 2086 3452 2089 3478
rect 2098 3458 2102 3461
rect 2098 3448 2102 3451
rect 2022 3332 2025 3347
rect 2054 3332 2057 3358
rect 2078 3352 2081 3448
rect 2118 3392 2121 3418
rect 2118 3372 2121 3378
rect 2102 3352 2105 3358
rect 2090 3348 2094 3351
rect 2114 3348 2118 3351
rect 2126 3351 2129 3548
rect 2166 3542 2169 3548
rect 2138 3538 2142 3541
rect 2134 3482 2137 3488
rect 2142 3482 2145 3538
rect 2146 3468 2150 3471
rect 2146 3458 2150 3461
rect 2158 3452 2161 3458
rect 2166 3392 2169 3528
rect 2174 3492 2177 3558
rect 2190 3522 2193 3548
rect 2214 3482 2217 3658
rect 2226 3638 2230 3641
rect 2238 3532 2241 3678
rect 2246 3512 2249 3818
rect 2266 3768 2270 3771
rect 2278 3752 2281 3758
rect 2262 3742 2265 3748
rect 2262 3702 2265 3728
rect 2262 3642 2265 3678
rect 2270 3662 2273 3748
rect 2286 3712 2289 3818
rect 2294 3682 2297 3718
rect 2302 3671 2305 3898
rect 2318 3842 2321 3918
rect 2406 3912 2409 3918
rect 2438 3892 2441 3918
rect 2494 3902 2497 3918
rect 2510 3882 2513 4118
rect 2518 4112 2521 4158
rect 2582 4152 2585 4218
rect 2590 4192 2593 4218
rect 2614 4182 2617 4218
rect 2610 4158 2614 4161
rect 2574 4132 2577 4138
rect 2598 4132 2601 4138
rect 2630 4132 2633 4248
rect 2698 4238 2702 4241
rect 2678 4232 2681 4238
rect 2582 4122 2585 4128
rect 2602 4118 2606 4121
rect 2526 4082 2529 4118
rect 2558 4082 2561 4098
rect 2598 4062 2601 4068
rect 2518 4042 2521 4048
rect 2534 4002 2537 4058
rect 2582 4022 2585 4058
rect 2590 4042 2593 4048
rect 2614 4042 2617 4118
rect 2622 4052 2625 4058
rect 2630 4052 2633 4128
rect 2646 4081 2649 4128
rect 2654 4102 2657 4218
rect 2662 4192 2665 4208
rect 2678 4172 2681 4228
rect 2710 4202 2713 4218
rect 2718 4212 2721 4248
rect 2774 4241 2777 4298
rect 2910 4292 2913 4318
rect 2858 4268 2862 4271
rect 2830 4262 2833 4268
rect 2786 4258 2790 4261
rect 2814 4252 2817 4258
rect 2838 4252 2841 4268
rect 2846 4252 2849 4258
rect 2774 4238 2782 4241
rect 2742 4232 2745 4238
rect 2790 4232 2793 4238
rect 2686 4162 2689 4168
rect 2678 4132 2681 4148
rect 2646 4078 2654 4081
rect 2638 4072 2641 4078
rect 2658 4068 2662 4071
rect 2622 4012 2625 4018
rect 2544 4003 2546 4007
rect 2550 4003 2553 4007
rect 2557 4003 2560 4007
rect 2534 3952 2537 3998
rect 2622 3972 2625 3978
rect 2598 3962 2601 3968
rect 2522 3948 2526 3951
rect 2554 3948 2558 3951
rect 2386 3878 2390 3881
rect 2434 3878 2438 3881
rect 2490 3878 2494 3881
rect 2442 3868 2446 3871
rect 2462 3862 2465 3868
rect 2362 3858 2366 3861
rect 2330 3838 2334 3841
rect 2342 3831 2345 3858
rect 2334 3828 2345 3831
rect 2310 3802 2313 3818
rect 2334 3792 2337 3828
rect 2342 3781 2345 3818
rect 2350 3812 2353 3848
rect 2358 3822 2361 3858
rect 2414 3852 2417 3858
rect 2374 3842 2377 3848
rect 2374 3782 2377 3788
rect 2342 3778 2353 3781
rect 2326 3772 2329 3778
rect 2310 3762 2313 3768
rect 2342 3762 2345 3768
rect 2314 3748 2318 3751
rect 2318 3682 2321 3718
rect 2326 3682 2329 3688
rect 2334 3682 2337 3718
rect 2342 3712 2345 3718
rect 2350 3712 2353 3778
rect 2398 3752 2401 3828
rect 2414 3792 2417 3808
rect 2422 3792 2425 3838
rect 2386 3748 2390 3751
rect 2398 3742 2401 3748
rect 2422 3742 2425 3748
rect 2358 3692 2361 3738
rect 2342 3682 2345 3688
rect 2394 3678 2398 3681
rect 2294 3668 2305 3671
rect 2282 3648 2286 3651
rect 2294 3642 2297 3668
rect 2302 3652 2305 3658
rect 2310 3652 2313 3668
rect 2350 3652 2353 3668
rect 2374 3652 2377 3678
rect 2430 3672 2433 3818
rect 2454 3752 2457 3858
rect 2470 3852 2473 3858
rect 2506 3848 2510 3851
rect 2466 3838 2470 3841
rect 2486 3812 2489 3838
rect 2518 3832 2521 3858
rect 2550 3842 2553 3938
rect 2582 3902 2585 3918
rect 2606 3892 2609 3948
rect 2614 3942 2617 3968
rect 2646 3962 2649 4018
rect 2670 4002 2673 4058
rect 2678 4032 2681 4128
rect 2718 4112 2721 4208
rect 2790 4192 2793 4218
rect 2798 4212 2801 4248
rect 2806 4222 2809 4248
rect 2850 4238 2854 4241
rect 2870 4241 2873 4288
rect 2910 4262 2913 4268
rect 2882 4258 2886 4261
rect 2870 4238 2878 4241
rect 2778 4188 2782 4191
rect 2798 4152 2801 4158
rect 2750 4112 2753 4147
rect 2766 4142 2769 4148
rect 2806 4142 2809 4178
rect 2830 4152 2833 4168
rect 2838 4142 2841 4228
rect 2846 4162 2849 4218
rect 2846 4152 2849 4158
rect 2862 4152 2865 4158
rect 2870 4142 2873 4158
rect 2878 4142 2881 4148
rect 2810 4118 2814 4121
rect 2686 4092 2689 4108
rect 2734 4072 2737 4078
rect 2754 4068 2758 4071
rect 2774 4062 2777 4068
rect 2846 4062 2849 4128
rect 2878 4122 2881 4128
rect 2886 4082 2889 4218
rect 2894 4212 2897 4248
rect 2918 4242 2921 4308
rect 2926 4282 2929 4328
rect 2934 4312 2937 4318
rect 2918 4192 2921 4228
rect 2926 4212 2929 4218
rect 2934 4192 2937 4268
rect 2950 4262 2953 4298
rect 2966 4292 2969 4328
rect 2982 4302 2985 4318
rect 2958 4252 2961 4278
rect 2982 4252 2985 4268
rect 2990 4262 2993 4288
rect 3006 4282 3009 4318
rect 3014 4272 3017 4278
rect 3038 4272 3041 4308
rect 3048 4303 3050 4307
rect 3054 4303 3057 4307
rect 3061 4303 3064 4307
rect 3078 4272 3081 4338
rect 3086 4302 3089 4348
rect 3234 4338 3238 4341
rect 3230 4292 3233 4318
rect 3238 4312 3241 4338
rect 3246 4322 3249 4358
rect 3254 4352 3257 4358
rect 3486 4352 3489 4358
rect 3558 4352 3561 4358
rect 3274 4348 3278 4351
rect 3418 4348 3422 4351
rect 3442 4348 3446 4351
rect 3474 4348 3478 4351
rect 3498 4348 3502 4351
rect 3514 4348 3518 4351
rect 3630 4351 3633 4398
rect 3622 4348 3633 4351
rect 3638 4352 3641 4358
rect 3670 4352 3673 4368
rect 3702 4352 3705 4398
rect 3766 4382 3769 4428
rect 3790 4402 3793 4428
rect 3830 4402 3833 4428
rect 3714 4358 3718 4361
rect 3750 4352 3753 4358
rect 3806 4352 3809 4398
rect 3862 4382 3865 4388
rect 3814 4352 3817 4358
rect 3738 4348 3742 4351
rect 3762 4348 3766 4351
rect 3786 4348 3790 4351
rect 3826 4348 3830 4351
rect 3262 4342 3265 4348
rect 3246 4292 3249 4318
rect 3270 4302 3273 4338
rect 3302 4322 3305 4328
rect 3334 4302 3337 4348
rect 3358 4342 3361 4348
rect 3366 4332 3369 4338
rect 3094 4282 3097 4288
rect 3142 4282 3145 4288
rect 3262 4282 3265 4298
rect 3390 4292 3393 4348
rect 3430 4341 3433 4348
rect 3430 4338 3441 4341
rect 3130 4278 3134 4281
rect 3330 4278 3334 4281
rect 3042 4248 3046 4251
rect 2942 4232 2945 4238
rect 2950 4232 2953 4248
rect 2966 4242 2969 4248
rect 3054 4222 3057 4268
rect 2942 4162 2945 4168
rect 2930 4158 2934 4161
rect 2898 4148 2902 4151
rect 2942 4142 2945 4148
rect 2894 4132 2897 4138
rect 2910 4092 2913 4128
rect 2942 4092 2945 4098
rect 2910 4062 2913 4088
rect 2826 4058 2830 4061
rect 2890 4058 2894 4061
rect 2922 4058 2926 4061
rect 2710 4052 2713 4058
rect 2698 4048 2702 4051
rect 2754 4048 2758 4051
rect 2778 4048 2782 4051
rect 2738 4038 2742 4041
rect 2786 4038 2790 4041
rect 2718 4032 2721 4038
rect 2798 4031 2801 4058
rect 2806 4042 2809 4048
rect 2814 4041 2817 4058
rect 2838 4042 2841 4048
rect 2814 4038 2822 4041
rect 2790 4028 2801 4031
rect 2630 3922 2633 3958
rect 2662 3932 2665 3938
rect 2670 3922 2673 3958
rect 2686 3942 2689 3968
rect 2694 3952 2697 3958
rect 2702 3952 2705 4018
rect 2574 3862 2577 3888
rect 2602 3858 2606 3861
rect 2562 3848 2566 3851
rect 2538 3828 2542 3831
rect 2446 3722 2449 3728
rect 2386 3658 2390 3661
rect 2410 3658 2414 3661
rect 2286 3612 2289 3628
rect 2286 3571 2289 3608
rect 2286 3568 2297 3571
rect 2294 3562 2297 3568
rect 2186 3478 2190 3481
rect 2142 3362 2145 3368
rect 2150 3362 2153 3378
rect 2174 3362 2177 3468
rect 2182 3431 2185 3448
rect 2190 3442 2193 3448
rect 2198 3432 2201 3478
rect 2214 3461 2217 3478
rect 2214 3458 2222 3461
rect 2246 3452 2249 3498
rect 2262 3492 2265 3547
rect 2302 3542 2305 3618
rect 2314 3588 2318 3591
rect 2314 3538 2318 3541
rect 2278 3532 2281 3538
rect 2302 3472 2305 3518
rect 2326 3492 2329 3648
rect 2254 3452 2257 3458
rect 2210 3448 2214 3451
rect 2234 3448 2238 3451
rect 2262 3442 2265 3468
rect 2234 3438 2238 3441
rect 2182 3428 2193 3431
rect 2190 3392 2193 3428
rect 2206 3422 2209 3428
rect 2238 3392 2241 3428
rect 2254 3372 2257 3418
rect 2278 3392 2281 3468
rect 2294 3462 2297 3468
rect 2290 3448 2294 3451
rect 2262 3362 2265 3368
rect 2310 3362 2313 3458
rect 2322 3448 2326 3451
rect 2334 3442 2337 3638
rect 2366 3632 2369 3648
rect 2386 3638 2390 3641
rect 2410 3638 2414 3641
rect 2422 3551 2425 3618
rect 2430 3562 2433 3588
rect 2438 3562 2441 3658
rect 2446 3582 2449 3678
rect 2462 3662 2465 3678
rect 2454 3652 2457 3658
rect 2478 3652 2481 3718
rect 2486 3652 2489 3808
rect 2544 3803 2546 3807
rect 2550 3803 2553 3807
rect 2557 3803 2560 3807
rect 2518 3762 2521 3768
rect 2530 3758 2534 3761
rect 2494 3742 2497 3758
rect 2538 3748 2542 3751
rect 2510 3742 2513 3748
rect 2574 3742 2577 3858
rect 2630 3852 2633 3918
rect 2638 3852 2641 3918
rect 2646 3872 2649 3888
rect 2678 3862 2681 3918
rect 2702 3912 2705 3948
rect 2598 3842 2601 3848
rect 2662 3842 2665 3858
rect 2678 3842 2681 3848
rect 2614 3832 2617 3838
rect 2642 3828 2646 3831
rect 2590 3752 2593 3818
rect 2622 3812 2625 3818
rect 2670 3802 2673 3818
rect 2538 3738 2542 3741
rect 2494 3662 2497 3668
rect 2474 3638 2478 3641
rect 2470 3612 2473 3628
rect 2462 3582 2465 3588
rect 2446 3562 2449 3578
rect 2458 3568 2462 3571
rect 2470 3562 2473 3608
rect 2378 3547 2382 3550
rect 2422 3548 2433 3551
rect 2430 3542 2433 3548
rect 2418 3538 2422 3541
rect 2418 3528 2422 3531
rect 2382 3511 2385 3528
rect 2382 3508 2393 3511
rect 2366 3482 2369 3498
rect 2342 3462 2345 3468
rect 2350 3462 2353 3478
rect 2366 3452 2369 3478
rect 2374 3462 2377 3468
rect 2338 3438 2342 3441
rect 2358 3392 2361 3448
rect 2382 3442 2385 3448
rect 2366 3362 2369 3368
rect 2122 3348 2129 3351
rect 2246 3358 2254 3361
rect 2098 3338 2102 3341
rect 2122 3338 2126 3341
rect 2134 3332 2137 3358
rect 2166 3352 2169 3358
rect 2174 3342 2177 3358
rect 2194 3348 2198 3351
rect 2182 3342 2185 3348
rect 2024 3303 2026 3307
rect 2030 3303 2033 3307
rect 2037 3303 2040 3307
rect 2054 3302 2057 3328
rect 2026 3288 2030 3291
rect 2094 3282 2097 3288
rect 2062 3272 2065 3278
rect 1982 3212 1985 3258
rect 2094 3252 2097 3259
rect 1950 3192 1953 3198
rect 1842 3168 1846 3171
rect 1658 3148 1662 3151
rect 1690 3148 1694 3151
rect 1730 3148 1734 3151
rect 1806 3151 1809 3158
rect 1918 3151 1921 3158
rect 1646 3122 1649 3138
rect 1686 3112 1689 3138
rect 1718 3112 1721 3138
rect 1694 3092 1697 3098
rect 1678 3072 1681 3078
rect 1726 3072 1729 3078
rect 1774 3072 1777 3148
rect 1990 3132 1993 3218
rect 2074 3168 2078 3171
rect 2082 3158 2086 3161
rect 2110 3152 2113 3328
rect 2126 3292 2129 3298
rect 2142 3182 2145 3208
rect 2166 3192 2169 3298
rect 2174 3282 2177 3338
rect 2190 3292 2193 3338
rect 2190 3282 2193 3288
rect 2010 3147 2014 3150
rect 2086 3148 2094 3151
rect 2086 3142 2089 3148
rect 2098 3138 2102 3141
rect 1790 3092 1793 3098
rect 1882 3088 1886 3091
rect 1918 3072 1921 3128
rect 1986 3088 1990 3091
rect 2014 3072 2017 3128
rect 2024 3103 2026 3107
rect 2030 3103 2033 3107
rect 2037 3103 2040 3107
rect 1758 3063 1761 3068
rect 1850 3059 1854 3062
rect 1582 3008 1593 3011
rect 1662 3012 1665 3059
rect 1520 3003 1522 3007
rect 1526 3003 1529 3007
rect 1533 3003 1536 3007
rect 1582 2992 1585 3008
rect 1530 2947 1534 2950
rect 1662 2951 1665 2978
rect 1758 2951 1761 3028
rect 1814 2952 1817 2968
rect 1846 2952 1849 3048
rect 1854 2992 1857 2998
rect 1870 2972 1873 3068
rect 1550 2942 1553 2948
rect 1738 2938 1742 2941
rect 1550 2872 1553 2938
rect 1520 2803 1522 2807
rect 1526 2803 1529 2807
rect 1533 2803 1536 2807
rect 1518 2751 1521 2768
rect 1550 2752 1553 2868
rect 1558 2852 1561 2859
rect 1558 2692 1561 2698
rect 1574 2672 1577 2898
rect 1590 2882 1593 2898
rect 1630 2882 1633 2898
rect 1662 2892 1665 2928
rect 1590 2872 1593 2878
rect 1662 2872 1665 2888
rect 1650 2868 1654 2871
rect 1598 2862 1601 2868
rect 1670 2862 1673 2908
rect 1678 2872 1681 2938
rect 1694 2912 1697 2918
rect 1774 2872 1777 2878
rect 1618 2858 1622 2861
rect 1642 2858 1646 2861
rect 1618 2848 1622 2851
rect 1650 2848 1654 2851
rect 1594 2748 1598 2751
rect 1614 2742 1617 2758
rect 1678 2752 1681 2768
rect 1582 2722 1585 2738
rect 1590 2732 1593 2738
rect 1590 2662 1593 2688
rect 1606 2652 1609 2718
rect 1614 2672 1617 2678
rect 1654 2672 1657 2678
rect 1622 2662 1625 2668
rect 1662 2662 1665 2748
rect 1686 2742 1689 2818
rect 1670 2692 1673 2698
rect 1642 2658 1646 2661
rect 1642 2648 1646 2651
rect 1520 2603 1522 2607
rect 1526 2603 1529 2607
rect 1533 2603 1536 2607
rect 1458 2588 1462 2591
rect 1542 2572 1545 2638
rect 1562 2588 1566 2591
rect 1598 2552 1601 2568
rect 1662 2552 1665 2578
rect 1350 2488 1358 2491
rect 1294 2463 1297 2468
rect 1294 2458 1297 2459
rect 1250 2438 1254 2441
rect 1254 2362 1257 2418
rect 1302 2372 1305 2468
rect 1322 2368 1326 2371
rect 1258 2348 1262 2351
rect 1262 2292 1265 2338
rect 1350 2292 1353 2488
rect 1374 2472 1377 2478
rect 1390 2452 1393 2459
rect 1398 2372 1401 2538
rect 1406 2432 1409 2548
rect 1518 2512 1521 2547
rect 1458 2488 1462 2491
rect 1470 2472 1473 2478
rect 1414 2361 1417 2368
rect 1410 2358 1417 2361
rect 1422 2352 1425 2418
rect 1486 2352 1489 2488
rect 1518 2482 1521 2498
rect 1534 2462 1537 2538
rect 1630 2532 1633 2547
rect 1646 2492 1649 2498
rect 1498 2458 1502 2461
rect 1510 2352 1513 2458
rect 1520 2403 1522 2407
rect 1526 2403 1529 2407
rect 1533 2403 1536 2407
rect 1542 2392 1545 2448
rect 1550 2412 1553 2418
rect 1358 2342 1361 2348
rect 1382 2342 1385 2348
rect 1366 2298 1374 2301
rect 1366 2292 1369 2298
rect 1382 2282 1385 2338
rect 1318 2272 1321 2278
rect 1382 2272 1385 2278
rect 1398 2263 1401 2268
rect 1250 2168 1254 2171
rect 1158 2132 1161 2138
rect 1198 2132 1201 2138
rect 1206 2132 1209 2138
rect 1230 2082 1233 2138
rect 1158 2042 1161 2078
rect 1202 2068 1206 2071
rect 1174 2062 1177 2068
rect 1222 2062 1225 2078
rect 1238 2062 1241 2078
rect 1262 2072 1265 2132
rect 1278 2082 1281 2228
rect 1310 2182 1313 2258
rect 1422 2222 1425 2348
rect 1446 2342 1449 2348
rect 1438 2312 1441 2318
rect 1438 2302 1441 2308
rect 1470 2282 1473 2288
rect 1478 2232 1481 2347
rect 1486 2272 1489 2298
rect 1550 2282 1553 2338
rect 1574 2302 1577 2468
rect 1634 2458 1638 2461
rect 1606 2352 1609 2438
rect 1662 2422 1665 2548
rect 1670 2502 1673 2668
rect 1678 2592 1681 2718
rect 1694 2672 1697 2758
rect 1726 2752 1729 2858
rect 1734 2792 1737 2848
rect 1730 2738 1734 2741
rect 1742 2732 1745 2868
rect 1766 2862 1769 2868
rect 1754 2848 1758 2851
rect 1750 2742 1753 2758
rect 1758 2752 1761 2768
rect 1782 2752 1785 2848
rect 1790 2762 1793 2888
rect 1798 2862 1801 2918
rect 1830 2892 1833 2918
rect 1846 2892 1849 2898
rect 1838 2882 1841 2888
rect 1806 2872 1809 2878
rect 1822 2872 1825 2878
rect 1834 2868 1838 2871
rect 1770 2748 1774 2751
rect 1790 2742 1793 2758
rect 1798 2752 1801 2778
rect 1806 2762 1809 2868
rect 1846 2752 1849 2868
rect 1902 2792 1905 2968
rect 1910 2922 1913 2948
rect 1918 2942 1921 3068
rect 1950 3052 1953 3059
rect 1966 2972 1969 3068
rect 2014 2942 2017 2947
rect 2030 2942 2033 3068
rect 2042 3059 2046 3062
rect 2062 3032 2065 3128
rect 2078 3072 2081 3128
rect 2094 3072 2097 3128
rect 2126 3111 2129 3158
rect 2142 3152 2145 3178
rect 2174 3172 2177 3278
rect 2190 3192 2193 3259
rect 2206 3232 2209 3358
rect 2230 3342 2233 3358
rect 2214 3312 2217 3328
rect 2222 3262 2225 3268
rect 2238 3261 2241 3348
rect 2246 3292 2249 3358
rect 2306 3348 2310 3351
rect 2338 3348 2342 3351
rect 2286 3342 2289 3348
rect 2278 3322 2281 3338
rect 2258 3318 2262 3321
rect 2278 3292 2281 3308
rect 2290 3288 2294 3291
rect 2250 3268 2254 3271
rect 2234 3258 2241 3261
rect 2258 3258 2262 3261
rect 2206 3202 2209 3228
rect 2214 3192 2217 3228
rect 2166 3152 2169 3168
rect 2142 3112 2145 3148
rect 2174 3142 2177 3168
rect 2162 3138 2166 3141
rect 2150 3132 2153 3138
rect 2182 3132 2185 3158
rect 2206 3142 2209 3168
rect 2126 3108 2137 3111
rect 2126 3092 2129 3098
rect 2106 3058 2110 3061
rect 2118 3022 2121 3038
rect 2134 3002 2137 3108
rect 2150 3082 2153 3128
rect 2158 3092 2161 3128
rect 2190 3122 2193 3128
rect 2154 3068 2158 3071
rect 2174 3062 2177 3108
rect 2222 3092 2225 3248
rect 2230 3182 2233 3258
rect 2246 3212 2249 3238
rect 2230 3162 2233 3168
rect 2238 3092 2241 3158
rect 2182 3072 2185 3078
rect 2214 3072 2217 3078
rect 2202 3058 2206 3061
rect 2142 2992 2145 3058
rect 2210 3048 2214 3051
rect 2218 3048 2222 3051
rect 2162 3038 2166 3041
rect 2158 2992 2161 3028
rect 2190 3002 2193 3038
rect 2166 2992 2169 2998
rect 2058 2938 2062 2941
rect 2122 2938 2126 2941
rect 2030 2932 2033 2938
rect 2134 2932 2137 2948
rect 2198 2942 2201 3048
rect 2238 3032 2241 3058
rect 2246 3022 2249 3208
rect 2254 3162 2257 3168
rect 2258 3148 2262 3151
rect 2254 3092 2257 3148
rect 2262 3102 2265 3138
rect 2254 3072 2257 3078
rect 2262 2982 2265 3058
rect 2262 2962 2265 2968
rect 2226 2947 2230 2950
rect 2270 2942 2273 3158
rect 2278 3152 2281 3248
rect 2310 3192 2313 3198
rect 2318 3152 2321 3338
rect 2342 3272 2345 3338
rect 2354 3328 2358 3331
rect 2374 3331 2377 3418
rect 2390 3352 2393 3508
rect 2414 3492 2417 3498
rect 2422 3482 2425 3488
rect 2438 3482 2441 3558
rect 2446 3542 2449 3548
rect 2478 3542 2481 3618
rect 2486 3592 2489 3648
rect 2502 3642 2505 3718
rect 2518 3652 2521 3738
rect 2538 3668 2542 3671
rect 2566 3662 2569 3698
rect 2590 3672 2593 3678
rect 2586 3658 2590 3661
rect 2554 3648 2558 3651
rect 2518 3632 2521 3648
rect 2530 3638 2534 3641
rect 2494 3612 2497 3618
rect 2544 3603 2546 3607
rect 2550 3603 2553 3607
rect 2557 3603 2560 3607
rect 2518 3592 2521 3598
rect 2486 3542 2489 3578
rect 2534 3572 2537 3578
rect 2506 3568 2510 3571
rect 2494 3562 2497 3568
rect 2546 3538 2550 3541
rect 2474 3518 2478 3521
rect 2486 3492 2489 3528
rect 2426 3468 2430 3471
rect 2458 3468 2462 3471
rect 2398 3392 2401 3468
rect 2414 3432 2417 3448
rect 2390 3342 2393 3348
rect 2370 3328 2377 3331
rect 2358 3302 2361 3328
rect 2370 3318 2374 3321
rect 2382 3292 2385 3338
rect 2390 3292 2393 3308
rect 2406 3272 2409 3278
rect 2350 3201 2353 3259
rect 2386 3248 2390 3251
rect 2398 3212 2401 3268
rect 2414 3252 2417 3428
rect 2438 3372 2441 3468
rect 2502 3462 2505 3478
rect 2446 3452 2449 3458
rect 2470 3442 2473 3458
rect 2482 3448 2486 3451
rect 2510 3451 2513 3538
rect 2526 3532 2529 3538
rect 2558 3532 2561 3538
rect 2566 3482 2569 3658
rect 2598 3652 2601 3768
rect 2606 3762 2609 3768
rect 2686 3762 2689 3908
rect 2710 3902 2713 3968
rect 2726 3941 2729 4018
rect 2750 3992 2753 4028
rect 2790 3982 2793 4028
rect 2798 4012 2801 4018
rect 2830 3982 2833 4018
rect 2826 3968 2830 3971
rect 2802 3958 2806 3961
rect 2734 3952 2737 3958
rect 2726 3938 2737 3941
rect 2722 3928 2726 3931
rect 2734 3922 2737 3938
rect 2742 3932 2745 3958
rect 2782 3942 2785 3948
rect 2838 3942 2841 3948
rect 2810 3938 2814 3941
rect 2774 3932 2777 3938
rect 2830 3932 2833 3938
rect 2802 3928 2806 3931
rect 2718 3902 2721 3918
rect 2702 3862 2705 3868
rect 2702 3792 2705 3838
rect 2702 3772 2705 3788
rect 2710 3782 2713 3898
rect 2718 3762 2721 3858
rect 2574 3642 2577 3648
rect 2526 3472 2529 3478
rect 2566 3462 2569 3478
rect 2502 3448 2513 3451
rect 2526 3452 2529 3458
rect 2486 3392 2489 3438
rect 2494 3422 2497 3448
rect 2486 3362 2489 3388
rect 2426 3268 2430 3271
rect 2438 3262 2441 3358
rect 2478 3342 2481 3348
rect 2450 3338 2454 3341
rect 2462 3302 2465 3328
rect 2502 3292 2505 3448
rect 2514 3438 2518 3441
rect 2544 3403 2546 3407
rect 2550 3403 2553 3407
rect 2557 3403 2560 3407
rect 2510 3362 2513 3398
rect 2522 3368 2526 3371
rect 2550 3362 2553 3388
rect 2566 3372 2569 3458
rect 2574 3442 2577 3638
rect 2598 3562 2601 3648
rect 2606 3632 2609 3718
rect 2622 3692 2625 3718
rect 2678 3672 2681 3718
rect 2686 3682 2689 3758
rect 2718 3751 2721 3758
rect 2714 3748 2721 3751
rect 2638 3662 2641 3668
rect 2654 3662 2657 3668
rect 2694 3662 2697 3748
rect 2702 3662 2705 3718
rect 2726 3692 2729 3878
rect 2750 3872 2753 3878
rect 2746 3858 2750 3861
rect 2742 3792 2745 3838
rect 2750 3792 2753 3848
rect 2758 3772 2761 3928
rect 2774 3842 2777 3848
rect 2782 3831 2785 3858
rect 2790 3842 2793 3848
rect 2798 3841 2801 3918
rect 2846 3912 2849 4058
rect 2898 4048 2902 4051
rect 2862 4022 2865 4048
rect 2862 3962 2865 4018
rect 2894 4002 2897 4018
rect 2890 3958 2894 3961
rect 2858 3928 2862 3931
rect 2798 3838 2806 3841
rect 2774 3828 2785 3831
rect 2774 3792 2777 3828
rect 2766 3772 2769 3788
rect 2774 3752 2777 3758
rect 2634 3648 2638 3651
rect 2638 3562 2641 3648
rect 2646 3642 2649 3648
rect 2662 3642 2665 3658
rect 2702 3642 2705 3648
rect 2686 3632 2689 3638
rect 2646 3562 2649 3568
rect 2654 3552 2657 3618
rect 2606 3532 2609 3538
rect 2582 3482 2585 3488
rect 2590 3441 2593 3518
rect 2622 3472 2625 3478
rect 2602 3458 2606 3461
rect 2626 3458 2630 3461
rect 2618 3448 2622 3451
rect 2590 3438 2598 3441
rect 2638 3441 2641 3518
rect 2654 3512 2657 3528
rect 2662 3482 2665 3588
rect 2670 3552 2673 3558
rect 2678 3542 2681 3618
rect 2694 3562 2697 3598
rect 2710 3572 2713 3678
rect 2726 3662 2729 3668
rect 2734 3651 2737 3728
rect 2742 3712 2745 3728
rect 2758 3672 2761 3678
rect 2774 3672 2777 3678
rect 2750 3662 2753 3668
rect 2726 3648 2737 3651
rect 2726 3622 2729 3648
rect 2742 3642 2745 3658
rect 2734 3632 2737 3638
rect 2686 3532 2689 3538
rect 2694 3492 2697 3518
rect 2662 3462 2665 3478
rect 2686 3462 2689 3468
rect 2710 3462 2713 3518
rect 2722 3468 2726 3471
rect 2654 3442 2657 3458
rect 2694 3452 2697 3458
rect 2734 3452 2737 3628
rect 2766 3552 2769 3618
rect 2774 3562 2777 3648
rect 2782 3572 2785 3818
rect 2798 3812 2801 3818
rect 2814 3792 2817 3858
rect 2822 3852 2825 3898
rect 2838 3862 2841 3868
rect 2830 3842 2833 3848
rect 2846 3842 2849 3858
rect 2854 3852 2857 3918
rect 2878 3862 2881 3868
rect 2886 3852 2889 3898
rect 2894 3881 2897 3918
rect 2910 3902 2913 4038
rect 2918 3992 2921 4058
rect 2930 4038 2934 4041
rect 2930 4018 2934 4021
rect 2930 3947 2934 3950
rect 2894 3878 2905 3881
rect 2894 3862 2897 3868
rect 2902 3852 2905 3878
rect 2910 3872 2913 3878
rect 2918 3862 2921 3908
rect 2942 3862 2945 3868
rect 2870 3842 2873 3848
rect 2806 3762 2809 3768
rect 2846 3752 2849 3828
rect 2854 3802 2857 3818
rect 2878 3792 2881 3818
rect 2858 3788 2862 3791
rect 2862 3772 2865 3778
rect 2894 3762 2897 3848
rect 2934 3762 2937 3818
rect 2950 3762 2953 4198
rect 2990 4172 2993 4218
rect 2974 4152 2977 4168
rect 2966 4102 2969 4148
rect 2998 4142 3001 4168
rect 2998 4072 3001 4138
rect 2994 4058 2998 4061
rect 2958 3952 2961 4038
rect 3022 4031 3025 4148
rect 3038 4142 3041 4148
rect 3078 4142 3081 4268
rect 3102 4262 3105 4278
rect 3174 4262 3177 4268
rect 3118 4182 3121 4218
rect 3142 4161 3145 4168
rect 3130 4148 3134 4151
rect 3154 4148 3158 4151
rect 3038 4132 3041 4138
rect 3048 4103 3050 4107
rect 3054 4103 3057 4107
rect 3061 4103 3064 4107
rect 3070 4082 3073 4098
rect 3078 4092 3081 4118
rect 3086 4082 3089 4128
rect 3070 4062 3073 4078
rect 3022 4028 3033 4031
rect 3030 3992 3033 4028
rect 3038 3992 3041 4058
rect 3046 4042 3049 4048
rect 3086 3992 3089 4078
rect 3094 4042 3097 4138
rect 3102 4102 3105 4138
rect 3166 4132 3169 4138
rect 3190 4132 3193 4138
rect 3198 4132 3201 4258
rect 3238 4172 3241 4248
rect 3246 4192 3249 4198
rect 3234 4168 3238 4171
rect 3246 4152 3249 4178
rect 3254 4162 3257 4268
rect 3262 4222 3265 4278
rect 3358 4262 3361 4288
rect 3438 4282 3441 4338
rect 3446 4322 3449 4348
rect 3486 4342 3489 4348
rect 3446 4292 3449 4298
rect 3314 4258 3318 4261
rect 3222 4142 3225 4148
rect 3254 4141 3257 4158
rect 3246 4138 3257 4141
rect 3174 4082 3177 4088
rect 3198 4082 3201 4128
rect 3130 4058 3134 4061
rect 3174 3992 3177 4068
rect 3186 4058 3190 4061
rect 3202 4058 3206 4061
rect 2994 3988 2998 3991
rect 3022 3952 3025 3968
rect 3094 3952 3097 3988
rect 3142 3962 3145 3968
rect 3162 3938 3169 3941
rect 3126 3932 3129 3938
rect 3006 3902 3009 3918
rect 3048 3903 3050 3907
rect 3054 3903 3057 3907
rect 3061 3903 3064 3907
rect 3142 3902 3145 3918
rect 3006 3892 3009 3898
rect 2982 3862 2985 3878
rect 3022 3862 3025 3868
rect 3006 3832 3009 3858
rect 3030 3852 3033 3888
rect 3038 3862 3041 3868
rect 3102 3862 3105 3868
rect 3074 3848 3078 3851
rect 3046 3842 3049 3848
rect 3066 3838 3070 3841
rect 2962 3768 2966 3771
rect 2890 3758 2894 3761
rect 2850 3748 2854 3751
rect 2878 3742 2881 3748
rect 2934 3742 2937 3748
rect 2974 3742 2977 3818
rect 3014 3782 3017 3838
rect 3026 3768 3030 3771
rect 3038 3762 3041 3818
rect 2986 3758 2990 3761
rect 3010 3758 3014 3761
rect 3014 3752 3017 3758
rect 2826 3738 2830 3741
rect 2914 3738 2918 3741
rect 3018 3738 3022 3741
rect 2790 3661 2793 3738
rect 2886 3732 2889 3738
rect 2942 3732 2945 3738
rect 2826 3728 2830 3731
rect 2914 3728 2918 3731
rect 2798 3722 2801 3728
rect 2926 3722 2929 3728
rect 2806 3702 2809 3718
rect 2902 3712 2905 3718
rect 2790 3658 2798 3661
rect 2790 3642 2793 3648
rect 2806 3642 2809 3678
rect 2830 3662 2833 3668
rect 2814 3642 2817 3648
rect 2786 3548 2790 3551
rect 2798 3541 2801 3638
rect 2822 3632 2825 3648
rect 2834 3638 2838 3641
rect 2834 3618 2838 3621
rect 2846 3592 2849 3668
rect 2854 3572 2857 3678
rect 2862 3642 2865 3708
rect 2902 3682 2905 3688
rect 2890 3678 2894 3681
rect 2906 3668 2910 3671
rect 2870 3652 2873 3658
rect 2926 3642 2929 3708
rect 2934 3641 2937 3658
rect 2942 3652 2945 3698
rect 2966 3692 2969 3738
rect 2998 3722 3001 3738
rect 3042 3728 3046 3731
rect 2970 3678 2974 3681
rect 2990 3672 2993 3718
rect 3014 3692 3017 3718
rect 3048 3703 3050 3707
rect 3054 3703 3057 3707
rect 3061 3703 3064 3707
rect 3062 3682 3065 3688
rect 2950 3662 2953 3668
rect 2966 3642 2969 3648
rect 2934 3638 2945 3641
rect 2862 3582 2865 3638
rect 2810 3558 2814 3561
rect 2842 3548 2846 3551
rect 2794 3538 2801 3541
rect 2666 3448 2670 3451
rect 2638 3438 2646 3441
rect 2690 3438 2694 3441
rect 2606 3392 2609 3418
rect 2614 3372 2617 3438
rect 2622 3392 2625 3438
rect 2586 3358 2590 3361
rect 2510 3302 2513 3348
rect 2526 3292 2529 3338
rect 2534 3292 2537 3338
rect 2550 3312 2553 3318
rect 2466 3288 2470 3291
rect 2558 3282 2561 3328
rect 2474 3268 2478 3271
rect 2494 3268 2502 3271
rect 2562 3268 2566 3271
rect 2462 3262 2465 3268
rect 2466 3248 2470 3251
rect 2454 3242 2457 3248
rect 2410 3238 2414 3241
rect 2494 3212 2497 3268
rect 2574 3262 2577 3338
rect 2590 3331 2593 3358
rect 2598 3352 2601 3358
rect 2606 3352 2609 3368
rect 2630 3362 2633 3378
rect 2646 3362 2649 3388
rect 2654 3382 2657 3418
rect 2666 3388 2670 3391
rect 2678 3362 2681 3408
rect 2686 3342 2689 3418
rect 2702 3392 2705 3448
rect 2722 3438 2726 3441
rect 2734 3352 2737 3398
rect 2742 3392 2745 3458
rect 2758 3441 2761 3518
rect 2754 3438 2761 3441
rect 2774 3442 2777 3518
rect 2782 3462 2785 3498
rect 2806 3462 2809 3518
rect 2798 3452 2801 3458
rect 2814 3452 2817 3518
rect 2822 3512 2825 3528
rect 2862 3482 2865 3508
rect 2822 3462 2825 3468
rect 2830 3452 2833 3478
rect 2838 3462 2841 3468
rect 2786 3448 2790 3451
rect 2846 3442 2849 3448
rect 2810 3438 2814 3441
rect 2758 3412 2761 3418
rect 2782 3392 2785 3418
rect 2750 3372 2753 3378
rect 2746 3368 2750 3371
rect 2778 3368 2782 3371
rect 2778 3358 2782 3361
rect 2738 3348 2742 3351
rect 2790 3342 2793 3358
rect 2822 3352 2825 3398
rect 2838 3391 2841 3418
rect 2854 3392 2857 3448
rect 2862 3422 2865 3478
rect 2870 3462 2873 3618
rect 2882 3568 2886 3571
rect 2890 3548 2894 3551
rect 2918 3532 2921 3538
rect 2878 3482 2881 3528
rect 2910 3492 2913 3518
rect 2918 3512 2921 3528
rect 2878 3472 2881 3478
rect 2894 3452 2897 3478
rect 2902 3462 2905 3468
rect 2926 3462 2929 3498
rect 2934 3472 2937 3618
rect 2942 3592 2945 3638
rect 2990 3592 2993 3598
rect 2998 3582 3001 3658
rect 2950 3572 2953 3578
rect 2942 3522 2945 3548
rect 2966 3532 2969 3538
rect 2966 3462 2969 3518
rect 2878 3442 2881 3448
rect 2910 3442 2913 3458
rect 2922 3448 2926 3451
rect 2934 3432 2937 3458
rect 2942 3442 2945 3448
rect 2958 3442 2961 3448
rect 2974 3442 2977 3578
rect 2982 3552 2985 3578
rect 3006 3572 3009 3638
rect 3014 3622 3017 3628
rect 3022 3612 3025 3678
rect 3030 3668 3038 3671
rect 3030 3592 3033 3668
rect 3038 3652 3041 3658
rect 3054 3642 3057 3648
rect 3070 3642 3073 3838
rect 3086 3832 3089 3858
rect 3110 3852 3113 3888
rect 3118 3862 3121 3868
rect 3126 3842 3129 3898
rect 3166 3892 3169 3938
rect 3182 3901 3185 4058
rect 3214 4052 3217 4138
rect 3226 4128 3230 4131
rect 3246 4092 3249 4138
rect 3262 4131 3265 4218
rect 3278 4192 3281 4228
rect 3270 4162 3273 4168
rect 3278 4152 3281 4178
rect 3286 4172 3289 4258
rect 3298 4248 3302 4251
rect 3338 4248 3342 4251
rect 3298 4238 3302 4241
rect 3310 4222 3313 4248
rect 3358 4242 3361 4248
rect 3302 4172 3305 4178
rect 3286 4142 3289 4158
rect 3310 4152 3313 4168
rect 3306 4148 3310 4151
rect 3254 4128 3265 4131
rect 3306 4138 3310 4141
rect 3234 4078 3238 4081
rect 3222 4052 3225 4058
rect 3198 4042 3201 4048
rect 3226 4038 3230 4041
rect 3174 3898 3185 3901
rect 3174 3892 3177 3898
rect 3142 3882 3145 3888
rect 3206 3872 3209 3938
rect 3086 3742 3089 3828
rect 3118 3762 3121 3818
rect 3094 3752 3097 3758
rect 3126 3752 3129 3758
rect 3142 3752 3145 3758
rect 3114 3748 3118 3751
rect 3194 3748 3198 3751
rect 3214 3751 3217 3998
rect 3238 3942 3241 4068
rect 3254 4062 3257 4128
rect 3262 4062 3265 4068
rect 3254 3962 3257 4058
rect 3262 4052 3265 4058
rect 3270 3992 3273 4138
rect 3278 4062 3281 4078
rect 3302 4072 3305 4108
rect 3310 4092 3313 4128
rect 3318 4081 3321 4158
rect 3326 4152 3329 4238
rect 3366 4191 3369 4268
rect 3374 4252 3377 4258
rect 3398 4252 3401 4278
rect 3430 4272 3433 4278
rect 3410 4258 3414 4261
rect 3382 4242 3385 4248
rect 3362 4188 3369 4191
rect 3374 4192 3377 4218
rect 3350 4162 3353 4168
rect 3358 4162 3361 4188
rect 3334 4112 3337 4148
rect 3350 4092 3353 4148
rect 3374 4142 3377 4148
rect 3366 4082 3369 4088
rect 3310 4078 3321 4081
rect 3302 4062 3305 4068
rect 3226 3938 3230 3941
rect 3254 3882 3257 3958
rect 3266 3948 3270 3951
rect 3290 3948 3294 3951
rect 3302 3942 3305 4058
rect 3310 4042 3313 4078
rect 3318 4052 3321 4068
rect 3326 4062 3329 4068
rect 3318 3952 3321 4048
rect 3334 3972 3337 4018
rect 3342 3992 3345 4058
rect 3358 3962 3361 4078
rect 3390 4062 3393 4138
rect 3398 4092 3401 4238
rect 3414 4162 3417 4258
rect 3422 4232 3425 4268
rect 3454 4262 3457 4268
rect 3446 4212 3449 4248
rect 3462 4232 3465 4268
rect 3470 4192 3473 4338
rect 3502 4332 3505 4348
rect 3478 4282 3481 4308
rect 3486 4292 3489 4298
rect 3518 4292 3521 4298
rect 3534 4272 3537 4338
rect 3542 4312 3545 4348
rect 3486 4252 3489 4268
rect 3502 4262 3505 4268
rect 3482 4248 3486 4251
rect 3478 4232 3481 4238
rect 3502 4192 3505 4248
rect 3510 4222 3513 4248
rect 3510 4192 3513 4208
rect 3450 4158 3454 4161
rect 3494 4152 3497 4178
rect 3526 4162 3529 4268
rect 3534 4252 3537 4268
rect 3542 4262 3545 4308
rect 3598 4302 3601 4348
rect 3622 4332 3625 4348
rect 3634 4338 3638 4341
rect 3634 4318 3638 4321
rect 3594 4288 3598 4291
rect 3614 4282 3617 4318
rect 3626 4288 3630 4291
rect 3646 4282 3649 4328
rect 3654 4282 3657 4348
rect 3698 4338 3702 4341
rect 3662 4332 3665 4338
rect 3678 4292 3681 4338
rect 3726 4332 3729 4338
rect 3686 4302 3689 4318
rect 3710 4292 3713 4308
rect 3670 4272 3673 4288
rect 3626 4268 3630 4271
rect 3658 4268 3662 4271
rect 3662 4262 3665 4268
rect 3642 4258 3649 4261
rect 3606 4252 3609 4258
rect 3558 4152 3561 4248
rect 3568 4203 3570 4207
rect 3574 4203 3577 4207
rect 3581 4203 3584 4207
rect 3434 4138 3438 4141
rect 3426 4128 3430 4131
rect 3434 4118 3438 4121
rect 3446 4082 3449 4148
rect 3474 4138 3478 4141
rect 3454 4092 3457 4138
rect 3486 4132 3489 4148
rect 3486 4122 3489 4128
rect 3450 4078 3454 4081
rect 3382 3992 3385 4058
rect 3406 3972 3409 4068
rect 3438 4058 3446 4061
rect 3438 3992 3441 4058
rect 3414 3982 3417 3988
rect 3338 3948 3342 3951
rect 3322 3938 3329 3941
rect 3314 3928 3318 3931
rect 3326 3882 3329 3938
rect 3214 3748 3222 3751
rect 3150 3742 3153 3748
rect 3166 3742 3169 3748
rect 3094 3702 3097 3718
rect 3102 3682 3105 3738
rect 3082 3658 3086 3661
rect 3110 3652 3113 3668
rect 3118 3662 3121 3738
rect 3130 3728 3134 3731
rect 3174 3692 3177 3718
rect 3214 3712 3217 3728
rect 3222 3722 3225 3748
rect 3134 3662 3137 3668
rect 3154 3658 3158 3661
rect 3166 3652 3169 3658
rect 3082 3648 3086 3651
rect 3150 3642 3153 3648
rect 3122 3638 3126 3641
rect 2994 3568 2998 3571
rect 3010 3558 3014 3561
rect 3014 3552 3017 3558
rect 2986 3548 2990 3551
rect 3046 3532 3049 3538
rect 3054 3532 3057 3638
rect 3174 3632 3177 3668
rect 3190 3652 3193 3668
rect 3182 3642 3185 3648
rect 3206 3642 3209 3678
rect 3230 3672 3233 3858
rect 3294 3852 3297 3859
rect 3274 3758 3278 3761
rect 3246 3742 3249 3748
rect 3254 3732 3257 3758
rect 3266 3748 3270 3751
rect 3270 3742 3273 3748
rect 3310 3742 3313 3868
rect 3350 3842 3353 3958
rect 3382 3952 3385 3958
rect 3374 3942 3377 3948
rect 3358 3932 3361 3938
rect 3382 3872 3385 3948
rect 3390 3902 3393 3968
rect 3406 3952 3409 3968
rect 3422 3962 3425 3968
rect 3406 3942 3409 3948
rect 3430 3942 3433 3958
rect 3438 3942 3441 3948
rect 3446 3911 3449 3968
rect 3454 3922 3457 4068
rect 3462 3932 3465 3978
rect 3478 3952 3481 4078
rect 3494 3992 3497 4148
rect 3502 4142 3505 4148
rect 3518 4128 3526 4131
rect 3502 4062 3505 4118
rect 3518 4092 3521 4128
rect 3514 4078 3518 4081
rect 3526 4072 3529 4128
rect 3550 4072 3553 4108
rect 3558 4092 3561 4098
rect 3566 4082 3569 4148
rect 3574 4132 3577 4138
rect 3582 4122 3585 4148
rect 3638 4132 3641 4168
rect 3574 4102 3577 4118
rect 3506 4058 3510 4061
rect 3510 3952 3513 3988
rect 3542 3952 3545 4048
rect 3550 3982 3553 4068
rect 3590 4062 3593 4128
rect 3630 4092 3633 4118
rect 3646 4092 3649 4258
rect 3654 4252 3657 4258
rect 3670 4152 3673 4258
rect 3678 4252 3681 4258
rect 3678 4152 3681 4168
rect 3678 4122 3681 4128
rect 3686 4112 3689 4118
rect 3598 4072 3601 4088
rect 3562 4058 3566 4061
rect 3586 4058 3590 4061
rect 3618 4058 3622 4061
rect 3602 4048 3606 4051
rect 3574 4042 3577 4048
rect 3630 4042 3633 4088
rect 3646 4082 3649 4088
rect 3650 4068 3654 4071
rect 3662 4062 3665 4098
rect 3682 4088 3686 4091
rect 3682 4078 3686 4081
rect 3662 4052 3665 4058
rect 3568 4003 3570 4007
rect 3574 4003 3577 4007
rect 3581 4003 3584 4007
rect 3566 3962 3569 3978
rect 3590 3972 3593 4038
rect 3554 3958 3561 3961
rect 3470 3942 3473 3948
rect 3518 3922 3521 3938
rect 3526 3932 3529 3948
rect 3550 3932 3553 3938
rect 3446 3908 3457 3911
rect 3454 3892 3457 3908
rect 3426 3878 3430 3881
rect 3426 3868 3430 3871
rect 3438 3870 3441 3878
rect 3398 3852 3401 3868
rect 3462 3862 3465 3888
rect 3494 3872 3497 3918
rect 3410 3858 3414 3861
rect 3514 3858 3518 3861
rect 3386 3818 3390 3821
rect 3414 3762 3417 3768
rect 3442 3758 3446 3761
rect 3326 3751 3329 3758
rect 3398 3752 3401 3758
rect 3406 3752 3409 3758
rect 3450 3748 3454 3751
rect 3518 3751 3521 3758
rect 3542 3752 3545 3868
rect 3558 3832 3561 3958
rect 3566 3882 3569 3958
rect 3582 3952 3585 3958
rect 3606 3952 3609 3958
rect 3582 3912 3585 3948
rect 3590 3942 3593 3948
rect 3614 3942 3617 3978
rect 3622 3962 3625 4018
rect 3646 3962 3649 4048
rect 3622 3942 3625 3948
rect 3630 3922 3633 3948
rect 3646 3922 3649 3958
rect 3654 3942 3657 3948
rect 3662 3932 3665 3938
rect 3670 3932 3673 4058
rect 3694 3982 3697 4258
rect 3702 4241 3705 4278
rect 3738 4268 3742 4271
rect 3710 4252 3713 4258
rect 3702 4238 3713 4241
rect 3710 4222 3713 4238
rect 3726 4142 3729 4258
rect 3742 4252 3745 4258
rect 3750 4232 3753 4348
rect 3794 4338 3798 4341
rect 3758 4312 3761 4338
rect 3774 4292 3777 4338
rect 3806 4332 3809 4348
rect 3822 4322 3825 4338
rect 3838 4332 3841 4338
rect 3846 4321 3849 4348
rect 3870 4332 3873 4348
rect 3878 4342 3881 4428
rect 3894 4352 3897 4428
rect 3918 4402 3921 4428
rect 3942 4402 3945 4428
rect 3966 4402 3969 4428
rect 3890 4348 3894 4351
rect 3838 4318 3849 4321
rect 3758 4262 3761 4268
rect 3782 4262 3785 4298
rect 3830 4282 3833 4298
rect 3838 4282 3841 4318
rect 3878 4292 3881 4298
rect 3886 4292 3889 4318
rect 3770 4258 3774 4261
rect 3758 4202 3761 4258
rect 3790 4252 3793 4268
rect 3818 4258 3822 4261
rect 3798 4252 3801 4258
rect 3762 4158 3766 4161
rect 3730 4138 3734 4141
rect 3714 4128 3718 4131
rect 3702 4032 3705 4058
rect 3714 4038 3718 4041
rect 3726 4032 3729 4058
rect 3734 4052 3737 4078
rect 3746 4068 3750 4071
rect 3750 4052 3753 4058
rect 3734 4022 3737 4048
rect 3758 4041 3761 4138
rect 3766 4132 3769 4148
rect 3766 4092 3769 4128
rect 3774 4072 3777 4138
rect 3782 4102 3785 4148
rect 3782 4082 3785 4098
rect 3798 4092 3801 4158
rect 3814 4152 3817 4208
rect 3822 4142 3825 4228
rect 3830 4152 3833 4158
rect 3814 4122 3817 4128
rect 3822 4112 3825 4138
rect 3770 4068 3774 4071
rect 3782 4062 3785 4078
rect 3802 4068 3806 4071
rect 3814 4062 3817 4078
rect 3838 4062 3841 4278
rect 3878 4271 3881 4288
rect 3874 4268 3881 4271
rect 3846 4232 3849 4268
rect 3866 4258 3870 4261
rect 3854 4212 3857 4258
rect 3870 4182 3873 4218
rect 3878 4212 3881 4268
rect 3894 4271 3897 4338
rect 3890 4268 3897 4271
rect 3902 4272 3905 4398
rect 3918 4362 3921 4368
rect 3926 4352 3929 4358
rect 3934 4342 3937 4378
rect 3942 4362 3945 4368
rect 3942 4342 3945 4348
rect 3918 4302 3921 4338
rect 3950 4331 3953 4398
rect 3982 4392 3985 4428
rect 4006 4402 4009 4428
rect 4022 4402 4025 4428
rect 3974 4362 3977 4368
rect 3990 4362 3993 4398
rect 4038 4372 4041 4428
rect 4062 4402 4065 4428
rect 4046 4382 4049 4388
rect 4022 4362 4025 4368
rect 3962 4358 3966 4361
rect 4062 4352 4065 4358
rect 3970 4348 3974 4351
rect 4002 4348 4006 4351
rect 4006 4342 4009 4348
rect 3942 4328 3953 4331
rect 3994 4338 3998 4341
rect 3922 4268 3929 4271
rect 3846 4092 3849 4118
rect 3854 4062 3857 4138
rect 3870 4132 3873 4168
rect 3862 4072 3865 4118
rect 3870 4082 3873 4128
rect 3834 4058 3838 4061
rect 3806 4052 3809 4058
rect 3870 4052 3873 4068
rect 3878 4062 3881 4198
rect 3886 4192 3889 4268
rect 3910 4252 3913 4258
rect 3894 4192 3897 4228
rect 3910 4162 3913 4168
rect 3894 4132 3897 4148
rect 3918 4142 3921 4258
rect 3926 4192 3929 4268
rect 3942 4252 3945 4328
rect 3958 4262 3961 4268
rect 3942 4202 3945 4248
rect 3966 4242 3969 4338
rect 3974 4272 3977 4298
rect 3982 4282 3985 4328
rect 4046 4322 4049 4348
rect 4054 4332 4057 4338
rect 4078 4322 4081 4338
rect 4090 4328 4094 4331
rect 4102 4322 4105 4428
rect 4126 4402 4129 4428
rect 4118 4352 4121 4378
rect 4142 4352 4145 4428
rect 4198 4372 4201 4378
rect 4214 4362 4217 4428
rect 4230 4382 4233 4428
rect 4342 4402 4345 4428
rect 4346 4398 4353 4401
rect 4154 4358 4158 4361
rect 4218 4358 4222 4361
rect 4146 4348 4150 4351
rect 4178 4348 4182 4351
rect 4218 4348 4222 4351
rect 4110 4332 4113 4348
rect 4198 4342 4201 4348
rect 4126 4332 4129 4338
rect 4142 4332 4145 4338
rect 4182 4322 4185 4338
rect 4046 4292 4049 4298
rect 3994 4288 3998 4291
rect 4038 4272 4041 4288
rect 4054 4282 4057 4308
rect 4062 4282 4065 4318
rect 3998 4262 4001 4268
rect 3974 4232 3977 4258
rect 3974 4202 3977 4228
rect 3950 4162 3953 4168
rect 3966 4162 3969 4168
rect 3974 4162 3977 4178
rect 3998 4151 4001 4178
rect 3994 4148 4001 4151
rect 4006 4152 4009 4258
rect 4014 4252 4017 4258
rect 4014 4192 4017 4208
rect 3950 4142 3953 4148
rect 3938 4138 3945 4141
rect 3926 4122 3929 4128
rect 3918 4082 3921 4108
rect 3890 4068 3894 4071
rect 3926 4062 3929 4108
rect 3770 4048 3774 4051
rect 3794 4048 3798 4051
rect 3758 4038 3769 4041
rect 3726 3962 3729 4018
rect 3766 3992 3769 4038
rect 3690 3938 3694 3941
rect 3570 3868 3574 3871
rect 3582 3862 3585 3898
rect 3602 3868 3609 3871
rect 3586 3858 3590 3861
rect 3594 3848 3598 3851
rect 3606 3822 3609 3868
rect 3568 3803 3570 3807
rect 3574 3803 3577 3807
rect 3581 3803 3584 3807
rect 3358 3732 3361 3748
rect 3462 3742 3465 3748
rect 3606 3742 3609 3778
rect 3410 3738 3414 3741
rect 3434 3738 3438 3741
rect 3294 3712 3297 3728
rect 3390 3712 3393 3718
rect 3214 3662 3217 3668
rect 3222 3652 3225 3658
rect 3214 3632 3217 3638
rect 3078 3592 3081 3628
rect 3222 3622 3225 3648
rect 3238 3642 3241 3698
rect 3262 3662 3265 3708
rect 3358 3682 3361 3698
rect 3430 3682 3433 3718
rect 3310 3662 3313 3668
rect 3338 3658 3342 3661
rect 3246 3631 3249 3658
rect 3294 3652 3297 3658
rect 3238 3628 3249 3631
rect 3254 3632 3257 3648
rect 3366 3642 3369 3648
rect 3102 3592 3105 3618
rect 3110 3562 3113 3578
rect 3062 3522 3065 3528
rect 3014 3502 3017 3518
rect 3048 3503 3050 3507
rect 3054 3503 3057 3507
rect 3061 3503 3064 3507
rect 3078 3482 3081 3558
rect 3086 3532 3089 3558
rect 3110 3552 3113 3558
rect 3126 3542 3129 3548
rect 3110 3531 3113 3538
rect 3134 3531 3137 3538
rect 3110 3528 3137 3531
rect 3094 3522 3097 3528
rect 3038 3472 3041 3478
rect 3010 3468 3014 3471
rect 2994 3458 2998 3461
rect 3034 3458 3038 3461
rect 2966 3432 2969 3438
rect 2886 3422 2889 3428
rect 2990 3422 2993 3448
rect 2998 3442 3001 3448
rect 3026 3438 3030 3441
rect 2838 3388 2846 3391
rect 2846 3372 2849 3378
rect 2830 3362 2833 3368
rect 2886 3362 2889 3398
rect 2902 3352 2905 3418
rect 2914 3368 2918 3371
rect 2926 3362 2929 3378
rect 2934 3362 2937 3418
rect 2974 3362 2977 3408
rect 2998 3372 3001 3378
rect 2962 3358 2966 3361
rect 3002 3358 3006 3361
rect 2850 3348 2854 3351
rect 2994 3348 2998 3351
rect 2806 3342 2809 3348
rect 2698 3338 2705 3341
rect 2590 3328 2601 3331
rect 2506 3248 2510 3251
rect 2538 3248 2542 3251
rect 2590 3242 2593 3318
rect 2598 3262 2601 3328
rect 2630 3312 2633 3318
rect 2654 3292 2657 3338
rect 2678 3292 2681 3338
rect 2690 3328 2694 3331
rect 2702 3292 2705 3338
rect 2970 3338 2974 3341
rect 2710 3312 2713 3328
rect 2766 3292 2769 3338
rect 2786 3318 2790 3321
rect 2814 3292 2817 3338
rect 2834 3318 2838 3321
rect 2846 3292 2849 3308
rect 2854 3292 2857 3338
rect 2874 3328 2878 3331
rect 2878 3322 2881 3328
rect 2886 3312 2889 3318
rect 2894 3292 2897 3308
rect 2902 3302 2905 3338
rect 2910 3332 2913 3338
rect 2918 3321 2921 3338
rect 2910 3318 2921 3321
rect 2910 3292 2913 3318
rect 2934 3312 2937 3318
rect 2926 3292 2929 3298
rect 2950 3292 2953 3338
rect 2958 3332 2961 3338
rect 3002 3318 3006 3321
rect 3014 3311 3017 3428
rect 3046 3392 3049 3448
rect 3034 3338 3041 3341
rect 3026 3328 3030 3331
rect 3006 3308 3017 3311
rect 3006 3292 3009 3308
rect 3030 3292 3033 3318
rect 3038 3292 3041 3338
rect 3054 3322 3057 3468
rect 3102 3462 3105 3468
rect 3086 3452 3089 3458
rect 3094 3452 3097 3458
rect 3110 3442 3113 3518
rect 3142 3472 3145 3618
rect 3238 3602 3241 3628
rect 3278 3622 3281 3628
rect 3246 3612 3249 3618
rect 3150 3562 3153 3568
rect 3190 3562 3193 3578
rect 3230 3562 3233 3568
rect 3150 3542 3153 3548
rect 3178 3538 3182 3541
rect 3150 3502 3153 3518
rect 3130 3458 3134 3461
rect 3162 3458 3166 3461
rect 3190 3452 3193 3558
rect 3222 3522 3225 3528
rect 3198 3452 3201 3518
rect 3210 3468 3214 3471
rect 3222 3462 3225 3488
rect 3122 3448 3126 3451
rect 3154 3448 3158 3451
rect 3218 3448 3222 3451
rect 3174 3442 3177 3448
rect 3230 3442 3233 3518
rect 3246 3492 3249 3538
rect 3254 3522 3257 3528
rect 3258 3468 3262 3471
rect 3270 3451 3273 3618
rect 3286 3562 3289 3568
rect 3310 3562 3313 3568
rect 3282 3538 3286 3541
rect 3318 3522 3321 3538
rect 3286 3472 3289 3518
rect 3282 3458 3286 3461
rect 3270 3448 3278 3451
rect 3294 3442 3297 3498
rect 3310 3442 3313 3518
rect 3318 3442 3321 3468
rect 3326 3462 3329 3588
rect 3334 3582 3337 3618
rect 3334 3562 3337 3568
rect 3374 3552 3377 3558
rect 3342 3542 3345 3548
rect 3358 3522 3361 3528
rect 3338 3518 3342 3521
rect 3358 3472 3361 3518
rect 3382 3492 3385 3668
rect 3414 3662 3417 3668
rect 3438 3662 3441 3718
rect 3450 3668 3454 3671
rect 3462 3662 3465 3738
rect 3534 3732 3537 3738
rect 3486 3702 3489 3728
rect 3486 3682 3489 3698
rect 3494 3692 3497 3698
rect 3534 3672 3537 3728
rect 3442 3658 3457 3661
rect 3546 3658 3550 3661
rect 3406 3642 3409 3648
rect 3406 3582 3409 3588
rect 3390 3562 3393 3568
rect 3398 3552 3401 3558
rect 3414 3542 3417 3658
rect 3442 3648 3446 3651
rect 3438 3562 3441 3608
rect 3426 3558 3430 3561
rect 3394 3538 3398 3541
rect 3430 3538 3438 3541
rect 3422 3531 3425 3538
rect 3414 3528 3425 3531
rect 3414 3492 3417 3528
rect 3430 3492 3433 3538
rect 3434 3468 3438 3471
rect 3374 3462 3377 3468
rect 3346 3458 3350 3461
rect 3390 3452 3393 3468
rect 3330 3448 3334 3451
rect 3146 3438 3150 3441
rect 3202 3438 3206 3441
rect 3354 3438 3358 3441
rect 3062 3322 3065 3348
rect 3048 3303 3050 3307
rect 3054 3303 3057 3307
rect 3061 3303 3064 3307
rect 2630 3282 2633 3288
rect 2974 3282 2977 3288
rect 2642 3268 2646 3271
rect 2914 3268 2918 3271
rect 2614 3262 2617 3268
rect 2544 3203 2546 3207
rect 2550 3203 2553 3207
rect 2557 3203 2560 3207
rect 2350 3198 2358 3201
rect 2366 3192 2369 3198
rect 2438 3162 2441 3168
rect 2462 3162 2465 3168
rect 2486 3162 2489 3168
rect 2510 3162 2513 3168
rect 2538 3158 2542 3161
rect 2290 3148 2294 3151
rect 2278 3092 2281 3108
rect 2294 3102 2297 3138
rect 2302 3132 2305 3138
rect 2318 3102 2321 3138
rect 2286 3098 2294 3101
rect 2286 3072 2289 3098
rect 2294 3062 2297 3088
rect 2318 3072 2321 3088
rect 2314 3068 2318 3071
rect 2302 3058 2310 3061
rect 2282 3048 2286 3051
rect 2294 3042 2297 3048
rect 2302 3031 2305 3058
rect 2294 3028 2305 3031
rect 2294 2992 2297 3028
rect 2310 3002 2313 3038
rect 2318 2992 2321 3028
rect 2334 2982 2337 3148
rect 2342 3132 2345 3158
rect 2398 3152 2401 3158
rect 2362 3148 2366 3151
rect 2386 3148 2390 3151
rect 2342 3092 2345 3108
rect 2374 3092 2377 3138
rect 2382 3072 2385 3098
rect 2362 3058 2366 3061
rect 2310 2972 2313 2978
rect 2150 2938 2158 2941
rect 2282 2938 2286 2941
rect 2150 2932 2153 2938
rect 1942 2892 1945 2898
rect 1950 2872 1953 2918
rect 2024 2903 2026 2907
rect 2030 2903 2033 2907
rect 2037 2903 2040 2907
rect 1910 2852 1913 2859
rect 1906 2778 1910 2781
rect 1926 2772 1929 2868
rect 2022 2862 2025 2868
rect 2006 2832 2009 2859
rect 1810 2748 1814 2751
rect 1822 2742 1825 2748
rect 1862 2742 1865 2758
rect 1886 2752 1889 2758
rect 1742 2722 1745 2728
rect 1758 2712 1761 2738
rect 1790 2722 1793 2738
rect 1702 2682 1705 2688
rect 1798 2682 1801 2688
rect 1766 2663 1769 2668
rect 1698 2658 1702 2661
rect 1734 2572 1737 2658
rect 1782 2592 1785 2598
rect 1794 2588 1798 2591
rect 1730 2548 1734 2551
rect 1678 2462 1681 2468
rect 1686 2452 1689 2458
rect 1662 2392 1665 2398
rect 1654 2362 1657 2368
rect 1702 2352 1705 2358
rect 1550 2272 1553 2278
rect 1590 2272 1593 2298
rect 1578 2268 1582 2271
rect 1466 2218 1470 2221
rect 1286 2152 1289 2178
rect 1294 2072 1297 2078
rect 1246 2062 1249 2068
rect 1258 2058 1262 2061
rect 1302 2052 1305 2058
rect 1318 2052 1321 2168
rect 1422 2162 1425 2168
rect 1438 2162 1441 2168
rect 1426 2158 1430 2161
rect 1466 2158 1470 2161
rect 1334 2142 1337 2147
rect 1414 2132 1417 2158
rect 1478 2142 1481 2218
rect 1520 2203 1522 2207
rect 1526 2203 1529 2207
rect 1533 2203 1536 2207
rect 1502 2152 1505 2158
rect 1442 2138 1446 2141
rect 1458 2138 1462 2141
rect 1458 2128 1462 2131
rect 1498 2128 1502 2131
rect 1326 2062 1329 2068
rect 1274 2048 1278 2051
rect 1326 2042 1329 2048
rect 1306 2038 1310 2041
rect 1118 2028 1129 2031
rect 1118 1972 1121 2018
rect 1126 1952 1129 2028
rect 1134 1952 1137 2018
rect 734 1922 737 1947
rect 758 1942 761 1948
rect 814 1942 817 1948
rect 830 1932 833 1947
rect 906 1938 910 1941
rect 974 1932 977 1938
rect 734 1892 737 1918
rect 770 1888 774 1891
rect 710 1863 713 1868
rect 634 1858 638 1861
rect 496 1803 498 1807
rect 502 1803 505 1807
rect 509 1803 512 1807
rect 486 1762 489 1768
rect 550 1751 553 1768
rect 582 1762 585 1798
rect 590 1772 593 1778
rect 598 1772 601 1858
rect 606 1852 609 1858
rect 622 1842 625 1848
rect 638 1842 641 1848
rect 678 1822 681 1858
rect 710 1778 718 1781
rect 478 1748 489 1751
rect 438 1672 441 1688
rect 366 1642 369 1648
rect 390 1632 393 1648
rect 342 1608 353 1611
rect 334 1512 337 1548
rect 342 1542 345 1608
rect 374 1582 377 1618
rect 398 1612 401 1618
rect 350 1532 353 1578
rect 374 1552 377 1568
rect 386 1558 390 1561
rect 390 1552 393 1558
rect 398 1552 401 1588
rect 374 1542 377 1548
rect 366 1532 369 1538
rect 398 1532 401 1538
rect 342 1522 345 1528
rect 350 1492 353 1498
rect 366 1492 369 1508
rect 382 1492 385 1518
rect 334 1482 337 1488
rect 282 1458 286 1461
rect 262 1442 265 1448
rect 286 1442 289 1448
rect 222 1392 225 1428
rect 214 1322 217 1368
rect 230 1352 233 1368
rect 262 1352 265 1408
rect 226 1278 230 1281
rect 154 1268 158 1271
rect 178 1268 182 1271
rect 6 1242 9 1248
rect 30 1182 33 1188
rect 54 1172 57 1178
rect 46 1152 49 1158
rect 70 1152 73 1178
rect 78 1162 81 1168
rect 110 1152 113 1268
rect 206 1262 209 1278
rect 230 1262 233 1268
rect 118 1192 121 1259
rect 186 1258 190 1261
rect 218 1258 222 1261
rect 166 1252 169 1258
rect 246 1252 249 1318
rect 278 1282 281 1358
rect 294 1351 297 1438
rect 318 1372 321 1458
rect 326 1352 329 1478
rect 350 1472 353 1488
rect 390 1482 393 1488
rect 406 1482 409 1668
rect 426 1648 430 1651
rect 454 1642 457 1738
rect 414 1532 417 1578
rect 422 1562 425 1618
rect 442 1558 446 1561
rect 454 1542 457 1558
rect 462 1552 465 1558
rect 422 1532 425 1538
rect 438 1492 441 1538
rect 450 1528 454 1531
rect 470 1522 473 1548
rect 478 1511 481 1658
rect 470 1508 481 1511
rect 486 1562 489 1748
rect 534 1672 537 1738
rect 582 1691 585 1758
rect 594 1748 598 1751
rect 638 1751 641 1758
rect 710 1752 713 1778
rect 726 1772 729 1888
rect 742 1862 745 1878
rect 758 1772 761 1778
rect 730 1768 734 1771
rect 718 1762 721 1768
rect 722 1748 726 1751
rect 574 1688 585 1691
rect 498 1659 502 1662
rect 538 1658 542 1661
rect 566 1642 569 1658
rect 574 1652 577 1688
rect 622 1672 625 1738
rect 670 1732 673 1748
rect 670 1692 673 1718
rect 606 1663 609 1668
rect 718 1662 721 1748
rect 734 1671 737 1768
rect 742 1692 745 1748
rect 766 1732 769 1878
rect 782 1852 785 1908
rect 902 1892 905 1898
rect 822 1872 825 1878
rect 806 1862 809 1868
rect 838 1863 841 1868
rect 870 1862 873 1868
rect 918 1862 921 1868
rect 934 1863 937 1898
rect 958 1872 961 1918
rect 1000 1903 1002 1907
rect 1006 1903 1009 1907
rect 1013 1903 1016 1907
rect 1022 1892 1025 1938
rect 1046 1932 1049 1948
rect 1062 1931 1065 1948
rect 1074 1938 1078 1941
rect 1062 1928 1070 1931
rect 1074 1928 1078 1931
rect 1054 1922 1057 1928
rect 1086 1901 1089 1948
rect 1126 1932 1129 1948
rect 1158 1942 1161 2038
rect 1334 2022 1337 2128
rect 1398 2122 1401 2128
rect 1406 2102 1409 2118
rect 1358 2072 1361 2088
rect 1382 2072 1385 2098
rect 1402 2088 1406 2091
rect 1422 2082 1425 2118
rect 1406 2072 1409 2078
rect 1346 2068 1350 2071
rect 1366 2062 1369 2068
rect 1438 2063 1441 2108
rect 1518 2092 1521 2098
rect 1342 2052 1345 2058
rect 1390 2052 1393 2058
rect 1370 2048 1374 2051
rect 1222 2002 1225 2018
rect 1174 1962 1177 1968
rect 1138 1938 1142 1941
rect 1138 1928 1142 1931
rect 1150 1922 1153 1928
rect 1094 1912 1097 1918
rect 1086 1898 1097 1901
rect 1030 1872 1033 1878
rect 958 1862 961 1868
rect 790 1852 793 1858
rect 782 1792 785 1848
rect 794 1838 798 1841
rect 838 1792 841 1848
rect 842 1768 846 1771
rect 862 1762 865 1818
rect 850 1748 854 1751
rect 894 1751 897 1758
rect 766 1682 769 1728
rect 798 1702 801 1748
rect 806 1742 809 1748
rect 830 1742 833 1748
rect 726 1668 737 1671
rect 690 1658 694 1661
rect 698 1638 702 1641
rect 496 1603 498 1607
rect 502 1603 505 1607
rect 509 1603 512 1607
rect 558 1592 561 1638
rect 686 1632 689 1638
rect 718 1631 721 1648
rect 726 1642 729 1668
rect 854 1662 857 1748
rect 910 1692 913 1838
rect 918 1752 921 1858
rect 1046 1822 1049 1859
rect 1094 1832 1097 1898
rect 1110 1892 1113 1898
rect 1118 1882 1121 1888
rect 1158 1882 1161 1908
rect 1118 1872 1121 1878
rect 994 1818 998 1821
rect 958 1792 961 1808
rect 994 1748 998 1751
rect 1010 1748 1014 1751
rect 1022 1732 1025 1768
rect 1030 1752 1033 1758
rect 1046 1742 1049 1758
rect 1054 1732 1057 1768
rect 1134 1762 1137 1818
rect 1122 1758 1126 1761
rect 1094 1752 1097 1758
rect 1086 1742 1089 1748
rect 1110 1742 1113 1748
rect 1090 1738 1094 1741
rect 1078 1732 1081 1738
rect 970 1728 974 1731
rect 1114 1728 1118 1731
rect 862 1662 865 1688
rect 974 1682 977 1718
rect 1000 1703 1002 1707
rect 1006 1703 1009 1707
rect 1013 1703 1016 1707
rect 1018 1688 1022 1691
rect 1126 1682 1129 1758
rect 1142 1712 1145 1738
rect 1158 1732 1161 1798
rect 1166 1772 1169 1948
rect 1190 1942 1193 1998
rect 1230 1952 1233 1958
rect 1202 1948 1206 1951
rect 1258 1948 1262 1951
rect 1214 1942 1217 1948
rect 1286 1942 1289 2018
rect 1366 1962 1369 2018
rect 1398 1992 1401 2038
rect 1430 1992 1433 1998
rect 1334 1951 1337 1958
rect 1366 1952 1369 1958
rect 1454 1952 1457 2068
rect 1462 1952 1465 2088
rect 1510 2082 1513 2088
rect 1470 2062 1473 2068
rect 1534 2062 1537 2118
rect 1550 2062 1553 2068
rect 1502 2022 1505 2028
rect 1520 2003 1522 2007
rect 1526 2003 1529 2007
rect 1533 2003 1536 2007
rect 1514 1958 1518 1961
rect 1514 1948 1518 1951
rect 1234 1938 1238 1941
rect 1250 1938 1254 1941
rect 1222 1922 1225 1938
rect 1270 1932 1273 1938
rect 1294 1932 1297 1938
rect 1406 1932 1409 1938
rect 1174 1852 1177 1918
rect 1182 1882 1185 1888
rect 1166 1762 1169 1768
rect 1134 1692 1137 1698
rect 1158 1692 1161 1708
rect 1174 1692 1177 1848
rect 1182 1792 1185 1838
rect 1190 1792 1193 1868
rect 1198 1862 1201 1918
rect 1206 1882 1209 1908
rect 1254 1872 1257 1908
rect 1262 1872 1265 1928
rect 1278 1872 1281 1928
rect 1286 1922 1289 1928
rect 1198 1802 1201 1858
rect 1230 1852 1233 1858
rect 1246 1852 1249 1858
rect 1218 1828 1222 1831
rect 1254 1772 1257 1868
rect 1274 1858 1278 1861
rect 1182 1752 1185 1758
rect 1254 1752 1257 1768
rect 1262 1752 1265 1858
rect 1294 1852 1297 1878
rect 1290 1848 1294 1851
rect 1270 1762 1273 1818
rect 1278 1762 1281 1768
rect 1302 1752 1305 1918
rect 1310 1872 1313 1878
rect 1326 1872 1329 1878
rect 1334 1852 1337 1918
rect 1382 1882 1385 1888
rect 1370 1878 1374 1881
rect 1350 1862 1353 1878
rect 1378 1868 1382 1871
rect 1406 1862 1409 1888
rect 1454 1882 1457 1948
rect 1470 1922 1473 1938
rect 1486 1932 1489 1948
rect 1506 1938 1510 1941
rect 1494 1922 1497 1938
rect 1534 1932 1537 1938
rect 1550 1932 1553 1948
rect 1558 1942 1561 2218
rect 1590 2142 1593 2268
rect 1606 2262 1609 2348
rect 1694 2342 1697 2348
rect 1726 2342 1729 2538
rect 1742 2492 1745 2508
rect 1806 2482 1809 2738
rect 1830 2722 1833 2738
rect 1830 2662 1833 2668
rect 1846 2602 1849 2728
rect 1894 2722 1897 2728
rect 1862 2663 1865 2718
rect 1894 2682 1897 2688
rect 1910 2572 1913 2768
rect 1926 2572 1929 2758
rect 1974 2751 1977 2778
rect 1990 2742 1993 2748
rect 1974 2663 1977 2688
rect 1990 2672 1993 2678
rect 2006 2572 2009 2808
rect 2022 2752 2025 2858
rect 2046 2782 2049 2908
rect 2054 2892 2057 2898
rect 2086 2862 2089 2868
rect 2118 2863 2121 2928
rect 2150 2882 2153 2888
rect 2182 2862 2185 2868
rect 2090 2778 2094 2781
rect 2134 2752 2137 2858
rect 2022 2742 2025 2748
rect 2154 2747 2158 2750
rect 2086 2732 2089 2738
rect 1962 2558 1966 2561
rect 1946 2548 1950 2551
rect 1834 2538 1838 2541
rect 1854 2532 1857 2547
rect 1886 2542 1889 2548
rect 1910 2542 1913 2548
rect 1938 2538 1942 2541
rect 1838 2492 1841 2528
rect 1758 2392 1761 2478
rect 1870 2472 1873 2538
rect 1774 2462 1777 2468
rect 1802 2459 1806 2462
rect 1870 2462 1873 2468
rect 1798 2372 1801 2418
rect 1894 2372 1897 2518
rect 1926 2491 1929 2518
rect 1926 2488 1937 2491
rect 1902 2452 1905 2459
rect 1934 2452 1937 2488
rect 1950 2462 1953 2548
rect 1982 2542 1985 2548
rect 2014 2542 2017 2728
rect 2024 2703 2026 2707
rect 2030 2703 2033 2707
rect 2037 2703 2040 2707
rect 2026 2688 2030 2691
rect 2054 2562 2057 2698
rect 2114 2688 2118 2691
rect 2102 2672 2105 2678
rect 2086 2622 2089 2659
rect 2110 2572 2113 2608
rect 2086 2552 2089 2558
rect 2142 2552 2145 2588
rect 1970 2538 1974 2541
rect 1986 2538 1990 2541
rect 2122 2538 2126 2541
rect 2146 2538 2150 2541
rect 1942 2371 1945 2458
rect 1934 2368 1945 2371
rect 1790 2342 1793 2348
rect 1646 2292 1649 2338
rect 1750 2292 1753 2318
rect 1670 2272 1673 2278
rect 1790 2272 1793 2338
rect 1798 2262 1801 2368
rect 1918 2351 1921 2358
rect 1822 2302 1825 2347
rect 1846 2292 1849 2298
rect 1886 2292 1889 2328
rect 1918 2282 1921 2328
rect 1886 2262 1889 2278
rect 1918 2263 1921 2268
rect 1686 2172 1689 2259
rect 1854 2182 1857 2218
rect 1774 2172 1777 2178
rect 1726 2152 1729 2158
rect 1698 2148 1702 2151
rect 1778 2148 1782 2151
rect 1854 2151 1857 2158
rect 1934 2152 1937 2368
rect 1950 2362 1953 2368
rect 1950 2292 1953 2328
rect 1958 2191 1961 2518
rect 1974 2502 1977 2528
rect 1974 2482 1977 2498
rect 1990 2451 1993 2518
rect 1998 2462 2001 2538
rect 2024 2503 2026 2507
rect 2030 2503 2033 2507
rect 2037 2503 2040 2507
rect 2094 2502 2097 2538
rect 2026 2488 2030 2491
rect 2050 2488 2054 2491
rect 2038 2482 2041 2488
rect 2078 2462 2081 2468
rect 1986 2448 1993 2451
rect 1950 2188 1961 2191
rect 1670 2142 1673 2148
rect 1686 2142 1689 2148
rect 1698 2138 1702 2141
rect 1654 2092 1657 2118
rect 1622 2082 1625 2088
rect 1670 2082 1673 2138
rect 1678 2132 1681 2138
rect 1570 2078 1574 2081
rect 1602 2078 1606 2081
rect 1590 2062 1593 2068
rect 1570 2058 1574 2061
rect 1574 2032 1577 2048
rect 1598 1972 1601 2078
rect 1678 2072 1681 2128
rect 1710 2122 1713 2148
rect 1730 2138 1734 2141
rect 1718 2132 1721 2138
rect 1742 2102 1745 2148
rect 1750 2112 1753 2148
rect 1778 2138 1782 2141
rect 1758 2132 1761 2138
rect 1698 2068 1702 2071
rect 1630 2032 1633 2068
rect 1638 2062 1641 2068
rect 1646 2022 1649 2068
rect 1662 2052 1665 2068
rect 1686 2062 1689 2068
rect 1670 2052 1673 2058
rect 1710 2052 1713 2098
rect 1662 2022 1665 2048
rect 1710 2042 1713 2048
rect 1718 2022 1721 2028
rect 1646 1982 1649 2018
rect 1614 1962 1617 1968
rect 1678 1962 1681 1968
rect 1642 1958 1646 1961
rect 1650 1948 1654 1951
rect 1622 1944 1625 1948
rect 1570 1938 1574 1941
rect 1638 1942 1641 1948
rect 1666 1938 1670 1941
rect 1614 1932 1617 1938
rect 1586 1928 1590 1931
rect 1562 1918 1566 1921
rect 1422 1872 1425 1878
rect 1346 1858 1350 1861
rect 1406 1852 1409 1858
rect 1418 1848 1422 1851
rect 1346 1838 1350 1841
rect 1182 1732 1185 1748
rect 1246 1742 1249 1748
rect 1190 1721 1193 1738
rect 1198 1732 1201 1738
rect 1254 1732 1257 1738
rect 1190 1718 1201 1721
rect 1198 1692 1201 1718
rect 1222 1712 1225 1718
rect 1278 1692 1281 1748
rect 1326 1742 1329 1748
rect 1342 1742 1345 1818
rect 1366 1772 1369 1818
rect 1454 1792 1457 1848
rect 1306 1738 1310 1741
rect 1358 1732 1361 1758
rect 1338 1728 1342 1731
rect 1286 1692 1289 1718
rect 1310 1692 1313 1718
rect 1166 1688 1174 1691
rect 1166 1682 1169 1688
rect 1222 1682 1225 1688
rect 1242 1678 1246 1681
rect 1306 1678 1310 1681
rect 1054 1672 1057 1678
rect 1174 1672 1177 1678
rect 1206 1672 1209 1678
rect 1154 1668 1158 1671
rect 1258 1668 1262 1671
rect 926 1662 929 1668
rect 718 1628 729 1631
rect 726 1622 729 1628
rect 514 1578 518 1581
rect 594 1578 598 1581
rect 618 1578 622 1581
rect 486 1512 489 1558
rect 502 1542 505 1548
rect 534 1532 537 1568
rect 542 1552 545 1558
rect 558 1522 561 1548
rect 402 1468 406 1471
rect 350 1362 353 1458
rect 362 1448 366 1451
rect 390 1372 393 1378
rect 390 1362 393 1368
rect 310 1342 313 1348
rect 326 1332 329 1338
rect 294 1292 297 1318
rect 302 1282 305 1308
rect 322 1278 326 1281
rect 254 1262 257 1268
rect 270 1252 273 1278
rect 278 1262 281 1278
rect 334 1272 337 1278
rect 286 1262 289 1268
rect 326 1262 329 1268
rect 306 1258 310 1261
rect 342 1252 345 1268
rect 246 1241 249 1248
rect 246 1238 257 1241
rect 170 1178 174 1181
rect 142 1151 145 1158
rect 6 1142 9 1148
rect 22 1122 25 1148
rect 30 1072 33 1078
rect 46 1062 49 1068
rect 54 1062 57 1088
rect 110 1072 113 1148
rect 238 1151 241 1228
rect 158 1142 161 1148
rect 206 1142 209 1148
rect 26 1058 30 1061
rect 6 1042 9 1048
rect 94 951 97 988
rect 6 942 9 948
rect 110 942 113 1068
rect 118 1063 121 1088
rect 118 1058 121 1059
rect 134 961 137 1118
rect 150 1072 153 1088
rect 230 1072 233 1138
rect 254 1072 257 1238
rect 270 1172 273 1248
rect 334 1192 337 1218
rect 342 1202 345 1248
rect 286 1162 289 1178
rect 298 1158 302 1161
rect 270 1082 273 1138
rect 318 1132 321 1138
rect 302 1112 305 1118
rect 270 1072 273 1078
rect 158 992 161 1058
rect 214 1012 217 1059
rect 246 1052 249 1058
rect 206 962 209 998
rect 246 972 249 978
rect 134 958 142 961
rect 202 948 206 951
rect 218 948 222 951
rect 218 938 222 941
rect 126 932 129 938
rect 186 928 190 931
rect 6 872 9 878
rect 22 862 25 928
rect 94 872 97 928
rect 30 852 33 868
rect 134 862 137 868
rect 150 862 153 868
rect 118 822 121 859
rect 70 751 73 798
rect 134 762 137 768
rect 146 758 150 761
rect 166 752 169 928
rect 182 882 185 918
rect 230 892 233 938
rect 222 872 225 878
rect 210 868 214 871
rect 238 852 241 868
rect 246 862 249 878
rect 254 872 257 1068
rect 294 1062 297 1098
rect 306 1068 310 1071
rect 274 1058 278 1061
rect 314 1058 318 1061
rect 302 1051 305 1058
rect 298 1048 305 1051
rect 278 1002 281 1048
rect 326 1002 329 1168
rect 334 1162 337 1188
rect 350 1172 353 1358
rect 378 1348 382 1351
rect 414 1342 417 1478
rect 430 1472 433 1478
rect 358 1322 361 1338
rect 366 1282 369 1308
rect 422 1282 425 1458
rect 446 1442 449 1448
rect 462 1422 465 1428
rect 438 1392 441 1398
rect 462 1392 465 1418
rect 434 1358 438 1361
rect 470 1352 473 1508
rect 566 1502 569 1538
rect 574 1532 577 1558
rect 630 1552 633 1558
rect 586 1548 590 1551
rect 594 1538 598 1541
rect 550 1472 553 1478
rect 582 1462 585 1528
rect 534 1452 537 1459
rect 602 1458 606 1461
rect 566 1452 569 1458
rect 614 1452 617 1548
rect 622 1462 625 1468
rect 594 1448 598 1451
rect 570 1438 574 1441
rect 478 1362 481 1418
rect 496 1403 498 1407
rect 502 1403 505 1407
rect 509 1403 512 1407
rect 558 1392 561 1438
rect 478 1352 481 1358
rect 574 1352 577 1358
rect 470 1342 473 1348
rect 542 1342 545 1348
rect 554 1338 561 1341
rect 362 1278 366 1281
rect 378 1268 382 1271
rect 366 1262 369 1268
rect 418 1258 422 1261
rect 430 1251 433 1318
rect 438 1292 441 1318
rect 494 1292 497 1338
rect 558 1332 561 1338
rect 470 1262 473 1268
rect 478 1262 481 1278
rect 446 1252 449 1258
rect 542 1252 545 1258
rect 550 1252 553 1288
rect 558 1272 561 1328
rect 582 1322 585 1358
rect 590 1292 593 1448
rect 614 1442 617 1448
rect 602 1378 606 1381
rect 598 1342 601 1348
rect 590 1272 593 1278
rect 598 1262 601 1338
rect 606 1332 609 1338
rect 614 1312 617 1318
rect 654 1312 657 1459
rect 662 1432 665 1547
rect 670 1472 673 1538
rect 718 1532 721 1618
rect 726 1592 729 1618
rect 718 1492 721 1518
rect 670 1342 673 1468
rect 734 1462 737 1658
rect 750 1592 753 1658
rect 766 1652 769 1659
rect 882 1658 886 1661
rect 842 1638 846 1641
rect 874 1638 878 1641
rect 742 1572 745 1578
rect 758 1551 761 1598
rect 754 1548 761 1551
rect 766 1552 769 1558
rect 774 1552 777 1608
rect 830 1592 833 1618
rect 838 1602 841 1618
rect 870 1612 873 1618
rect 894 1612 897 1648
rect 910 1602 913 1618
rect 958 1592 961 1659
rect 782 1572 785 1578
rect 966 1572 969 1668
rect 1270 1662 1273 1678
rect 1318 1672 1321 1678
rect 1286 1662 1289 1668
rect 982 1592 985 1608
rect 882 1568 886 1571
rect 790 1552 793 1558
rect 822 1551 825 1558
rect 918 1551 921 1568
rect 806 1532 809 1538
rect 902 1532 905 1538
rect 758 1472 761 1478
rect 866 1468 870 1471
rect 806 1462 809 1468
rect 718 1372 721 1378
rect 734 1371 737 1418
rect 726 1368 737 1371
rect 678 1351 681 1358
rect 710 1352 713 1358
rect 726 1352 729 1368
rect 694 1332 697 1338
rect 622 1292 625 1298
rect 734 1292 737 1358
rect 742 1342 745 1438
rect 782 1372 785 1418
rect 762 1348 766 1351
rect 774 1342 777 1358
rect 702 1262 705 1268
rect 718 1262 721 1268
rect 430 1248 438 1251
rect 406 1172 409 1248
rect 514 1228 518 1231
rect 496 1203 498 1207
rect 502 1203 505 1207
rect 509 1203 512 1207
rect 406 1151 409 1158
rect 446 1152 449 1198
rect 542 1192 545 1238
rect 566 1231 569 1258
rect 578 1238 582 1241
rect 566 1228 577 1231
rect 566 1192 569 1218
rect 574 1212 577 1228
rect 454 1152 457 1168
rect 478 1162 481 1168
rect 598 1162 601 1248
rect 606 1242 609 1258
rect 614 1162 617 1238
rect 678 1232 681 1258
rect 654 1162 657 1168
rect 466 1158 470 1161
rect 558 1152 561 1158
rect 438 1142 441 1148
rect 470 1142 473 1148
rect 398 1122 401 1138
rect 346 1118 350 1121
rect 334 1052 337 1118
rect 342 1042 345 1118
rect 414 1092 417 1108
rect 438 1072 441 1138
rect 446 1092 449 1138
rect 478 1102 481 1148
rect 542 1142 545 1148
rect 566 1142 569 1158
rect 582 1152 585 1158
rect 574 1142 577 1148
rect 518 1138 526 1141
rect 478 1092 481 1098
rect 458 1078 462 1081
rect 486 1072 489 1118
rect 418 1068 422 1071
rect 354 1058 358 1061
rect 358 1022 361 1028
rect 326 992 329 998
rect 310 962 313 968
rect 262 892 265 948
rect 278 932 281 958
rect 358 952 361 958
rect 290 948 294 951
rect 310 942 313 948
rect 322 938 326 941
rect 286 932 289 938
rect 366 932 369 1068
rect 434 1058 438 1061
rect 382 1032 385 1038
rect 390 1032 393 1058
rect 374 1012 377 1018
rect 390 992 393 1018
rect 390 962 393 988
rect 398 962 401 1048
rect 406 982 409 1048
rect 422 982 425 988
rect 386 948 390 951
rect 382 932 385 938
rect 270 902 273 928
rect 270 882 273 898
rect 222 762 225 828
rect 138 748 142 751
rect 178 748 182 751
rect 146 738 150 741
rect 166 732 169 748
rect 222 742 225 748
rect 178 738 182 741
rect 202 738 206 741
rect 230 732 233 788
rect 254 752 257 868
rect 286 862 289 868
rect 302 792 305 859
rect 358 852 361 918
rect 378 858 382 861
rect 370 838 374 841
rect 318 792 321 798
rect 302 772 305 778
rect 322 768 326 771
rect 282 758 286 761
rect 334 752 337 828
rect 390 761 393 918
rect 386 758 393 761
rect 6 692 9 718
rect 22 662 25 688
rect 70 662 73 728
rect 102 722 105 728
rect 126 672 129 688
rect 90 659 94 662
rect 6 642 9 648
rect 30 622 33 648
rect 22 618 30 621
rect 22 552 25 618
rect 30 572 33 578
rect 70 572 73 658
rect 134 652 137 718
rect 142 692 145 728
rect 182 722 185 728
rect 150 702 153 718
rect 142 662 145 668
rect 138 648 142 651
rect 142 582 145 648
rect 158 642 161 648
rect 166 622 169 658
rect 174 652 177 708
rect 182 692 185 718
rect 198 662 201 728
rect 230 722 233 728
rect 206 672 209 678
rect 214 672 217 698
rect 222 662 225 688
rect 246 662 249 668
rect 234 658 238 661
rect 182 652 185 658
rect 190 652 193 658
rect 174 551 177 578
rect 114 548 118 551
rect 6 542 9 548
rect 198 502 201 658
rect 242 648 246 651
rect 254 642 257 748
rect 262 742 265 748
rect 302 732 305 748
rect 314 738 318 741
rect 342 712 345 758
rect 362 748 366 751
rect 354 738 358 741
rect 270 662 273 678
rect 286 642 289 648
rect 254 592 257 618
rect 262 572 265 638
rect 254 562 257 568
rect 278 562 281 618
rect 278 552 281 558
rect 206 542 209 548
rect 6 442 9 448
rect 22 362 25 458
rect 54 452 57 459
rect 78 372 81 378
rect 34 348 38 351
rect 6 322 9 338
rect 22 332 25 338
rect 46 332 49 358
rect 74 348 78 351
rect 30 322 33 328
rect 6 242 9 248
rect 22 192 25 258
rect 38 152 41 268
rect 54 263 57 318
rect 86 272 89 458
rect 126 452 129 488
rect 162 458 166 461
rect 190 452 193 459
rect 222 452 225 468
rect 254 462 257 548
rect 294 542 297 688
rect 306 658 310 661
rect 322 648 326 651
rect 326 551 329 558
rect 310 542 313 548
rect 238 452 241 458
rect 122 438 126 441
rect 230 432 233 448
rect 238 432 241 438
rect 118 362 121 368
rect 126 362 129 368
rect 126 342 129 348
rect 98 338 102 341
rect 118 272 121 318
rect 126 282 129 318
rect 142 272 145 368
rect 222 362 225 378
rect 194 348 198 351
rect 226 348 230 351
rect 174 342 177 348
rect 238 342 241 348
rect 246 342 249 388
rect 254 352 257 438
rect 262 412 265 488
rect 270 462 273 498
rect 278 472 281 478
rect 286 461 289 518
rect 294 492 297 538
rect 334 502 337 658
rect 342 652 345 708
rect 362 658 366 661
rect 346 638 350 641
rect 318 462 321 468
rect 278 458 289 461
rect 298 458 302 461
rect 334 461 337 498
rect 334 458 342 461
rect 270 422 273 428
rect 262 352 265 408
rect 278 362 281 458
rect 286 442 289 448
rect 294 432 297 448
rect 302 442 305 448
rect 350 442 353 638
rect 358 632 361 638
rect 366 632 369 648
rect 374 641 377 718
rect 390 642 393 658
rect 398 652 401 958
rect 406 942 409 948
rect 430 882 433 1058
rect 438 952 441 1048
rect 446 952 449 1018
rect 496 1003 498 1007
rect 502 1003 505 1007
rect 509 1003 512 1007
rect 454 972 457 978
rect 482 968 486 971
rect 470 952 473 958
rect 494 952 497 968
rect 506 958 510 961
rect 438 912 441 948
rect 450 938 457 941
rect 446 932 449 938
rect 446 892 449 898
rect 430 762 433 878
rect 406 722 409 738
rect 414 712 417 748
rect 422 722 425 728
rect 406 672 409 698
rect 414 692 417 708
rect 438 702 441 868
rect 446 752 449 758
rect 454 742 457 938
rect 494 932 497 938
rect 518 932 521 1138
rect 530 1128 534 1131
rect 526 1062 529 1078
rect 550 1052 553 1058
rect 574 992 577 1138
rect 598 1092 601 1158
rect 638 1152 641 1158
rect 646 1152 649 1158
rect 670 1152 673 1158
rect 610 1138 614 1141
rect 614 1112 617 1138
rect 622 1122 625 1138
rect 654 1101 657 1118
rect 670 1112 673 1138
rect 678 1112 681 1228
rect 710 1192 713 1208
rect 718 1172 721 1178
rect 698 1158 702 1161
rect 714 1148 718 1151
rect 646 1098 657 1101
rect 582 1072 585 1088
rect 598 1062 601 1068
rect 598 972 601 1058
rect 614 1042 617 1059
rect 550 942 553 947
rect 462 751 465 908
rect 550 872 553 928
rect 482 858 486 861
rect 506 859 510 862
rect 496 803 498 807
rect 502 803 505 807
rect 509 803 512 807
rect 470 752 473 758
rect 462 748 470 751
rect 530 748 534 751
rect 454 712 457 718
rect 478 682 481 748
rect 498 738 502 741
rect 398 642 401 648
rect 374 638 382 641
rect 390 602 393 618
rect 390 582 393 588
rect 358 552 361 558
rect 406 522 409 668
rect 478 662 481 668
rect 518 662 521 668
rect 526 652 529 658
rect 534 642 537 678
rect 542 671 545 848
rect 550 842 553 858
rect 558 852 561 958
rect 598 912 601 968
rect 622 942 625 988
rect 646 962 649 1098
rect 682 1088 686 1091
rect 654 972 657 978
rect 662 972 665 1078
rect 694 1062 697 1148
rect 702 1092 705 1148
rect 682 1058 686 1061
rect 694 1052 697 1058
rect 634 948 638 951
rect 614 922 617 938
rect 598 872 601 908
rect 566 842 569 858
rect 574 842 577 848
rect 566 782 569 788
rect 558 762 561 768
rect 574 752 577 758
rect 550 682 553 718
rect 558 712 561 738
rect 574 712 577 738
rect 582 712 585 728
rect 542 668 553 671
rect 542 642 545 658
rect 550 652 553 668
rect 422 551 425 598
rect 462 591 465 618
rect 496 603 498 607
rect 502 603 505 607
rect 509 603 512 607
rect 454 588 465 591
rect 526 592 529 638
rect 582 621 585 668
rect 590 652 593 658
rect 614 652 617 918
rect 622 862 625 898
rect 646 812 649 878
rect 662 852 665 968
rect 670 952 673 1048
rect 702 1042 705 1078
rect 726 1072 729 1218
rect 734 1192 737 1198
rect 742 1172 745 1338
rect 782 1272 785 1358
rect 814 1312 817 1468
rect 878 1462 881 1488
rect 918 1482 921 1488
rect 926 1482 929 1568
rect 886 1472 889 1478
rect 902 1462 905 1478
rect 926 1452 929 1478
rect 966 1471 969 1528
rect 962 1468 969 1471
rect 982 1462 985 1578
rect 994 1558 998 1561
rect 1006 1542 1009 1548
rect 1046 1542 1049 1548
rect 1054 1542 1057 1548
rect 990 1472 993 1538
rect 1002 1528 1006 1531
rect 1000 1503 1002 1507
rect 1006 1503 1009 1507
rect 1013 1503 1016 1507
rect 998 1472 1001 1478
rect 1018 1468 1022 1471
rect 998 1452 1001 1458
rect 898 1448 902 1451
rect 962 1448 966 1451
rect 986 1448 990 1451
rect 934 1442 937 1448
rect 834 1418 838 1421
rect 838 1342 841 1348
rect 846 1342 849 1348
rect 894 1342 897 1388
rect 910 1372 913 1418
rect 926 1352 929 1378
rect 942 1362 945 1448
rect 950 1382 953 1418
rect 982 1392 985 1438
rect 946 1358 950 1361
rect 966 1352 969 1388
rect 974 1362 977 1368
rect 926 1332 929 1348
rect 1014 1342 1017 1388
rect 1022 1352 1025 1358
rect 1030 1351 1033 1518
rect 1054 1512 1057 1528
rect 1062 1501 1065 1598
rect 1070 1522 1073 1659
rect 1210 1658 1214 1661
rect 1078 1562 1081 1578
rect 1118 1562 1121 1588
rect 1078 1552 1081 1558
rect 1118 1542 1121 1548
rect 1086 1532 1089 1538
rect 1054 1498 1065 1501
rect 1038 1452 1041 1458
rect 1046 1452 1049 1458
rect 1042 1438 1046 1441
rect 1038 1362 1041 1368
rect 1026 1348 1033 1351
rect 938 1338 942 1341
rect 994 1338 998 1341
rect 1034 1338 1038 1341
rect 906 1328 913 1331
rect 946 1328 950 1331
rect 790 1272 793 1278
rect 838 1272 841 1328
rect 866 1318 870 1321
rect 846 1262 849 1298
rect 862 1292 865 1308
rect 870 1282 873 1288
rect 854 1272 857 1278
rect 894 1262 897 1298
rect 910 1292 913 1328
rect 910 1282 913 1288
rect 942 1282 945 1318
rect 958 1302 961 1318
rect 990 1292 993 1338
rect 1046 1332 1049 1418
rect 1054 1352 1057 1498
rect 1070 1442 1073 1468
rect 1078 1462 1081 1518
rect 1110 1472 1113 1518
rect 1126 1492 1129 1648
rect 1142 1602 1145 1658
rect 1254 1652 1257 1658
rect 1326 1652 1329 1688
rect 1350 1681 1353 1718
rect 1374 1691 1377 1788
rect 1462 1781 1465 1858
rect 1478 1792 1481 1918
rect 1534 1892 1537 1908
rect 1630 1892 1633 1918
rect 1694 1892 1697 1948
rect 1702 1942 1705 2018
rect 1726 1992 1729 2068
rect 1734 2052 1737 2078
rect 1766 2072 1769 2088
rect 1742 2052 1745 2058
rect 1550 1872 1553 1878
rect 1638 1872 1641 1878
rect 1502 1842 1505 1868
rect 1566 1863 1569 1868
rect 1686 1862 1689 1868
rect 1634 1858 1638 1861
rect 1454 1778 1465 1781
rect 1422 1752 1425 1758
rect 1390 1742 1393 1747
rect 1342 1678 1353 1681
rect 1366 1688 1377 1691
rect 1342 1672 1345 1678
rect 1366 1672 1369 1688
rect 1446 1682 1449 1748
rect 1454 1722 1457 1778
rect 1502 1752 1505 1838
rect 1520 1803 1522 1807
rect 1526 1803 1529 1807
rect 1533 1803 1536 1807
rect 1566 1792 1569 1808
rect 1354 1668 1358 1671
rect 1134 1532 1137 1588
rect 1146 1558 1150 1561
rect 1202 1558 1206 1561
rect 1158 1552 1161 1558
rect 1198 1542 1201 1558
rect 1214 1542 1217 1548
rect 1222 1542 1225 1548
rect 1270 1542 1273 1558
rect 1294 1542 1297 1618
rect 1186 1538 1190 1541
rect 1158 1532 1161 1538
rect 1202 1528 1206 1531
rect 1242 1518 1246 1521
rect 1134 1472 1137 1478
rect 1098 1458 1102 1461
rect 1106 1458 1110 1461
rect 1098 1448 1102 1451
rect 1122 1438 1129 1441
rect 1102 1362 1105 1368
rect 1062 1342 1065 1348
rect 1000 1303 1002 1307
rect 1006 1303 1009 1307
rect 1013 1303 1016 1307
rect 1022 1272 1025 1298
rect 1046 1282 1049 1298
rect 906 1268 910 1271
rect 950 1262 953 1268
rect 1022 1262 1025 1268
rect 1054 1252 1057 1268
rect 914 1248 918 1251
rect 878 1242 881 1248
rect 810 1218 814 1221
rect 742 1082 745 1168
rect 758 1162 761 1168
rect 754 1148 758 1151
rect 786 1148 790 1151
rect 766 1142 769 1148
rect 806 1092 809 1208
rect 882 1168 886 1171
rect 918 1151 921 1168
rect 974 1162 977 1218
rect 982 1192 985 1218
rect 990 1162 993 1168
rect 830 1132 833 1148
rect 854 1142 857 1148
rect 902 1142 905 1148
rect 838 1063 841 1088
rect 854 1072 857 1138
rect 902 1092 905 1128
rect 942 1072 945 1118
rect 914 1068 918 1071
rect 954 1068 958 1071
rect 746 1059 750 1062
rect 694 1032 697 1038
rect 702 952 705 958
rect 670 872 673 948
rect 742 942 745 948
rect 790 942 793 1038
rect 854 972 857 1068
rect 958 1052 961 1058
rect 926 1042 929 1048
rect 910 992 913 1028
rect 870 982 873 988
rect 806 951 809 958
rect 678 882 681 888
rect 798 872 801 908
rect 854 902 857 968
rect 918 962 921 1018
rect 898 958 902 961
rect 922 958 926 961
rect 934 952 937 1048
rect 958 992 961 1048
rect 974 1042 977 1158
rect 990 1071 993 1158
rect 1006 1152 1009 1218
rect 1014 1162 1017 1168
rect 1000 1103 1002 1107
rect 1006 1103 1009 1107
rect 1013 1103 1016 1107
rect 1022 1082 1025 1238
rect 1030 1142 1033 1158
rect 1038 1152 1041 1248
rect 1062 1242 1065 1338
rect 1070 1332 1073 1348
rect 1078 1342 1081 1358
rect 1110 1352 1113 1358
rect 1126 1352 1129 1438
rect 1134 1432 1137 1468
rect 1142 1392 1145 1518
rect 1310 1482 1313 1618
rect 1326 1572 1329 1648
rect 1318 1542 1321 1558
rect 1326 1532 1329 1538
rect 1226 1478 1230 1481
rect 1150 1472 1153 1478
rect 1174 1462 1177 1468
rect 1186 1458 1190 1461
rect 1202 1458 1206 1461
rect 1150 1452 1153 1458
rect 1170 1448 1174 1451
rect 1186 1448 1190 1451
rect 1198 1442 1201 1448
rect 1158 1362 1161 1418
rect 1214 1412 1217 1478
rect 1246 1462 1249 1478
rect 1270 1472 1273 1478
rect 1318 1472 1321 1518
rect 1334 1492 1337 1618
rect 1342 1552 1345 1598
rect 1358 1572 1361 1618
rect 1366 1602 1369 1668
rect 1414 1662 1417 1668
rect 1386 1628 1390 1631
rect 1446 1622 1449 1659
rect 1366 1562 1369 1578
rect 1406 1572 1409 1578
rect 1362 1548 1366 1551
rect 1342 1542 1345 1548
rect 1350 1532 1353 1548
rect 1374 1532 1377 1568
rect 1394 1548 1398 1551
rect 1414 1542 1417 1558
rect 1398 1532 1401 1538
rect 1350 1492 1353 1528
rect 1326 1472 1329 1478
rect 1374 1472 1377 1528
rect 1430 1502 1433 1538
rect 1382 1472 1385 1488
rect 1438 1482 1441 1488
rect 1430 1472 1433 1478
rect 1282 1468 1286 1471
rect 1258 1438 1262 1441
rect 1170 1368 1174 1371
rect 1178 1358 1182 1361
rect 1210 1358 1214 1361
rect 1134 1352 1137 1358
rect 1154 1348 1158 1351
rect 1178 1348 1182 1351
rect 1202 1348 1206 1351
rect 1086 1342 1089 1348
rect 1078 1311 1081 1338
rect 1086 1322 1089 1338
rect 1094 1332 1097 1338
rect 1126 1332 1129 1338
rect 1158 1332 1161 1338
rect 1114 1328 1118 1331
rect 1070 1308 1081 1311
rect 1070 1292 1073 1308
rect 1082 1278 1086 1281
rect 1082 1268 1086 1271
rect 1094 1202 1097 1268
rect 1102 1262 1105 1318
rect 1190 1292 1193 1328
rect 1110 1282 1113 1288
rect 1118 1282 1121 1288
rect 1126 1272 1129 1288
rect 1198 1282 1201 1348
rect 1214 1302 1217 1318
rect 1178 1268 1182 1271
rect 1118 1172 1121 1198
rect 1142 1192 1145 1258
rect 1182 1242 1185 1248
rect 1154 1238 1158 1241
rect 1198 1202 1201 1268
rect 1206 1262 1209 1268
rect 1222 1252 1225 1408
rect 1246 1372 1249 1418
rect 1270 1412 1273 1448
rect 1286 1392 1289 1468
rect 1298 1458 1302 1461
rect 1314 1458 1318 1461
rect 1298 1448 1302 1451
rect 1230 1342 1233 1368
rect 1242 1358 1246 1361
rect 1238 1352 1241 1358
rect 1254 1352 1257 1358
rect 1254 1322 1257 1338
rect 1238 1302 1241 1318
rect 1254 1278 1257 1298
rect 1262 1292 1265 1358
rect 1282 1338 1286 1341
rect 1294 1331 1297 1358
rect 1310 1342 1313 1418
rect 1326 1392 1329 1448
rect 1338 1358 1342 1361
rect 1358 1342 1361 1348
rect 1374 1341 1377 1458
rect 1382 1362 1385 1368
rect 1390 1362 1393 1368
rect 1370 1338 1377 1341
rect 1398 1342 1401 1418
rect 1454 1362 1457 1618
rect 1478 1542 1481 1638
rect 1494 1612 1497 1748
rect 1502 1742 1505 1748
rect 1574 1731 1577 1778
rect 1594 1768 1598 1771
rect 1582 1762 1585 1768
rect 1610 1758 1614 1761
rect 1602 1748 1606 1751
rect 1630 1751 1633 1828
rect 1638 1772 1641 1778
rect 1686 1772 1689 1848
rect 1686 1752 1689 1768
rect 1626 1748 1633 1751
rect 1582 1732 1585 1738
rect 1574 1728 1582 1731
rect 1534 1672 1537 1688
rect 1550 1672 1553 1678
rect 1598 1672 1601 1678
rect 1606 1672 1609 1718
rect 1578 1658 1582 1661
rect 1522 1648 1526 1651
rect 1520 1603 1522 1607
rect 1526 1603 1529 1607
rect 1533 1603 1536 1607
rect 1550 1572 1553 1658
rect 1614 1642 1617 1658
rect 1622 1642 1625 1658
rect 1614 1622 1617 1628
rect 1630 1612 1633 1748
rect 1654 1702 1657 1748
rect 1662 1732 1665 1738
rect 1674 1718 1678 1721
rect 1686 1712 1689 1738
rect 1694 1692 1697 1818
rect 1702 1792 1705 1938
rect 1710 1862 1713 1978
rect 1726 1952 1729 1988
rect 1750 1952 1753 2068
rect 1786 2059 1790 2062
rect 1758 1992 1761 2038
rect 1806 2022 1809 2128
rect 1830 2062 1833 2148
rect 1950 2151 1953 2188
rect 1850 2088 1854 2091
rect 1886 2082 1889 2118
rect 1886 2062 1889 2068
rect 1918 2063 1921 2078
rect 1934 2072 1937 2138
rect 1966 2082 1969 2358
rect 1974 2352 1977 2358
rect 1998 2352 2001 2418
rect 2074 2347 2078 2350
rect 1990 2312 1993 2328
rect 1982 2262 1985 2278
rect 1998 2202 2001 2318
rect 2024 2303 2026 2307
rect 2030 2303 2033 2307
rect 2037 2303 2040 2307
rect 2014 2252 2017 2259
rect 2030 2142 2033 2268
rect 2046 2151 2049 2298
rect 2070 2272 2073 2338
rect 2094 2262 2097 2408
rect 2102 2371 2105 2518
rect 2126 2472 2129 2508
rect 2142 2472 2145 2478
rect 2110 2463 2113 2468
rect 2150 2462 2153 2538
rect 2102 2368 2113 2371
rect 2110 2362 2113 2368
rect 2114 2348 2118 2351
rect 2130 2348 2134 2351
rect 2150 2342 2153 2418
rect 2158 2362 2161 2718
rect 2174 2572 2177 2798
rect 2198 2791 2201 2938
rect 2350 2932 2353 3038
rect 2230 2902 2233 2928
rect 2254 2918 2262 2921
rect 2230 2872 2233 2898
rect 2242 2888 2246 2891
rect 2214 2863 2217 2868
rect 2194 2788 2201 2791
rect 2254 2782 2257 2918
rect 2262 2791 2265 2838
rect 2262 2788 2273 2791
rect 2182 2682 2185 2688
rect 2182 2652 2185 2659
rect 2198 2572 2201 2778
rect 2214 2682 2217 2698
rect 2222 2682 2225 2738
rect 2254 2732 2257 2747
rect 2270 2742 2273 2788
rect 2286 2752 2289 2928
rect 2302 2912 2305 2928
rect 2350 2891 2353 2928
rect 2346 2888 2353 2891
rect 2326 2862 2329 2868
rect 2310 2852 2313 2859
rect 2262 2682 2265 2698
rect 2286 2682 2289 2738
rect 2238 2662 2241 2668
rect 2234 2628 2238 2631
rect 2238 2592 2241 2598
rect 2214 2562 2217 2568
rect 2238 2552 2241 2568
rect 2166 2452 2169 2518
rect 2174 2502 2177 2538
rect 2182 2482 2185 2498
rect 2178 2468 2182 2471
rect 2174 2352 2177 2358
rect 2150 2312 2153 2328
rect 2182 2322 2185 2458
rect 2190 2452 2193 2518
rect 2198 2342 2201 2538
rect 2246 2522 2249 2678
rect 2286 2662 2289 2668
rect 2258 2648 2262 2651
rect 2246 2501 2249 2518
rect 2238 2498 2249 2501
rect 2206 2462 2209 2498
rect 2206 2452 2209 2458
rect 2222 2352 2225 2448
rect 2158 2302 2161 2318
rect 2198 2312 2201 2328
rect 2206 2312 2209 2328
rect 2158 2272 2161 2278
rect 2154 2228 2158 2231
rect 2166 2191 2169 2308
rect 2198 2262 2201 2298
rect 2230 2292 2233 2348
rect 2206 2272 2209 2278
rect 2214 2272 2217 2278
rect 2238 2272 2241 2498
rect 2246 2452 2249 2488
rect 2262 2481 2265 2528
rect 2270 2492 2273 2538
rect 2254 2478 2265 2481
rect 2254 2462 2257 2478
rect 2262 2462 2265 2468
rect 2246 2442 2249 2448
rect 2246 2362 2249 2368
rect 2278 2362 2281 2518
rect 2286 2502 2289 2618
rect 2294 2572 2297 2778
rect 2358 2772 2361 3048
rect 2382 2942 2385 2947
rect 2366 2902 2369 2938
rect 2398 2932 2401 3118
rect 2406 3092 2409 3158
rect 2414 3152 2417 3158
rect 2478 3142 2481 3148
rect 2574 3142 2577 3208
rect 2598 3152 2601 3178
rect 2606 3162 2609 3258
rect 2614 3242 2617 3248
rect 2622 3212 2625 3268
rect 2662 3252 2665 3268
rect 2670 3262 2673 3268
rect 2710 3262 2713 3268
rect 2718 3262 2721 3268
rect 2750 3262 2753 3268
rect 2642 3248 2646 3251
rect 2682 3248 2686 3251
rect 2710 3251 2713 3258
rect 2710 3248 2721 3251
rect 2622 3152 2625 3158
rect 2458 3138 2462 3141
rect 2506 3138 2510 3141
rect 2618 3138 2622 3141
rect 2430 3132 2433 3138
rect 2526 3132 2529 3138
rect 2466 3118 2470 3121
rect 2482 3118 2486 3121
rect 2414 3112 2417 3118
rect 2414 3072 2417 3078
rect 2438 3072 2441 3118
rect 2494 3092 2497 3128
rect 2502 3118 2510 3121
rect 2538 3118 2542 3121
rect 2482 3068 2486 3071
rect 2418 3058 2422 3061
rect 2406 3012 2409 3038
rect 2414 2962 2417 2968
rect 2430 2952 2433 3068
rect 2454 3062 2457 3068
rect 2438 3042 2441 3048
rect 2462 3041 2465 3058
rect 2474 3048 2478 3051
rect 2502 3051 2505 3118
rect 2510 3082 2513 3108
rect 2526 3072 2529 3078
rect 2514 3068 2518 3071
rect 2494 3048 2505 3051
rect 2514 3048 2518 3051
rect 2462 3038 2473 3041
rect 2470 2972 2473 3038
rect 2458 2948 2462 2951
rect 2486 2942 2489 2948
rect 2374 2862 2377 2868
rect 2382 2772 2385 2928
rect 2414 2912 2417 2918
rect 2430 2912 2433 2938
rect 2438 2922 2441 2928
rect 2446 2922 2449 2928
rect 2398 2841 2401 2908
rect 2434 2888 2438 2891
rect 2422 2862 2425 2868
rect 2406 2852 2409 2859
rect 2398 2838 2409 2841
rect 2406 2772 2409 2838
rect 2438 2772 2441 2868
rect 2454 2842 2457 2938
rect 2478 2932 2481 2938
rect 2474 2858 2478 2861
rect 2302 2758 2334 2761
rect 2302 2742 2305 2758
rect 2330 2748 2334 2751
rect 2310 2742 2313 2748
rect 2318 2712 2321 2748
rect 2346 2738 2350 2741
rect 2386 2738 2390 2741
rect 2410 2738 2414 2741
rect 2310 2682 2313 2698
rect 2302 2652 2305 2658
rect 2302 2592 2305 2628
rect 2318 2572 2321 2708
rect 2334 2672 2337 2738
rect 2334 2662 2337 2668
rect 2350 2662 2353 2718
rect 2366 2692 2369 2738
rect 2402 2718 2406 2721
rect 2374 2702 2377 2718
rect 2386 2688 2390 2691
rect 2310 2532 2313 2548
rect 2318 2542 2321 2548
rect 2294 2521 2297 2528
rect 2294 2518 2305 2521
rect 2294 2482 2297 2508
rect 2302 2462 2305 2518
rect 2302 2402 2305 2458
rect 2318 2392 2321 2418
rect 2342 2412 2345 2658
rect 2354 2648 2358 2651
rect 2382 2632 2385 2658
rect 2422 2612 2425 2658
rect 2430 2652 2433 2718
rect 2438 2712 2441 2728
rect 2446 2712 2449 2748
rect 2358 2562 2361 2608
rect 2358 2552 2361 2558
rect 2390 2551 2393 2588
rect 2426 2558 2430 2561
rect 2446 2552 2449 2708
rect 2454 2692 2457 2838
rect 2478 2762 2481 2828
rect 2494 2782 2497 3048
rect 2510 2962 2513 3048
rect 2502 2952 2505 2958
rect 2514 2948 2518 2951
rect 2510 2932 2513 2938
rect 2526 2892 2529 3068
rect 2550 3062 2553 3138
rect 2582 3102 2585 3118
rect 2598 3092 2601 3138
rect 2618 3128 2625 3131
rect 2562 3068 2566 3071
rect 2610 3068 2614 3071
rect 2598 3062 2601 3068
rect 2534 3032 2537 3038
rect 2544 3003 2546 3007
rect 2550 3003 2553 3007
rect 2557 3003 2560 3007
rect 2566 2992 2569 3058
rect 2534 2942 2537 2948
rect 2542 2892 2545 2958
rect 2574 2951 2577 3058
rect 2602 3048 2606 3051
rect 2590 3042 2593 3048
rect 2570 2948 2577 2951
rect 2566 2942 2569 2948
rect 2566 2872 2569 2938
rect 2590 2932 2593 2978
rect 2622 2972 2625 3128
rect 2630 3092 2633 3158
rect 2630 3052 2633 3088
rect 2638 2972 2641 3238
rect 2694 3212 2697 3248
rect 2678 3162 2681 3208
rect 2710 3192 2713 3238
rect 2646 3158 2654 3161
rect 2666 3158 2670 3161
rect 2646 3142 2649 3148
rect 2646 3112 2649 3138
rect 2650 3068 2654 3071
rect 2662 3061 2665 3138
rect 2670 3092 2673 3138
rect 2678 3132 2681 3138
rect 2694 3112 2697 3138
rect 2694 3098 2702 3101
rect 2678 3072 2681 3078
rect 2658 3058 2665 3061
rect 2646 2972 2649 3058
rect 2674 3048 2678 3051
rect 2662 2962 2665 3048
rect 2694 2972 2697 3098
rect 2702 3042 2705 3058
rect 2710 3052 2713 3118
rect 2718 3092 2721 3248
rect 2742 3222 2745 3258
rect 2766 3252 2769 3268
rect 2726 3152 2729 3198
rect 2734 3162 2737 3208
rect 2742 3142 2745 3218
rect 2750 3142 2753 3218
rect 2798 3202 2801 3258
rect 2806 3222 2809 3268
rect 2822 3242 2825 3248
rect 2822 3192 2825 3208
rect 2774 3162 2777 3168
rect 2782 3162 2785 3168
rect 2806 3142 2809 3148
rect 2738 3118 2742 3121
rect 2750 3112 2753 3138
rect 2734 3102 2737 3108
rect 2726 3042 2729 3048
rect 2734 2992 2737 3098
rect 2758 3092 2761 3138
rect 2798 3132 2801 3138
rect 2770 3118 2774 3121
rect 2774 3092 2777 3108
rect 2750 3061 2753 3068
rect 2750 3058 2761 3061
rect 2746 3048 2750 3051
rect 2758 3022 2761 3058
rect 2758 2992 2761 3018
rect 2766 2981 2769 3068
rect 2758 2978 2769 2981
rect 2686 2942 2689 2948
rect 2602 2938 2606 2941
rect 2626 2938 2630 2941
rect 2666 2938 2670 2941
rect 2614 2872 2617 2918
rect 2630 2872 2633 2878
rect 2502 2863 2505 2868
rect 2518 2782 2521 2868
rect 2566 2862 2569 2868
rect 2606 2862 2609 2868
rect 2534 2852 2537 2858
rect 2544 2803 2546 2807
rect 2550 2803 2553 2807
rect 2557 2803 2560 2807
rect 2574 2802 2577 2858
rect 2598 2842 2601 2858
rect 2622 2852 2625 2858
rect 2610 2848 2614 2851
rect 2542 2772 2545 2778
rect 2614 2762 2617 2768
rect 2462 2742 2465 2748
rect 2486 2742 2489 2758
rect 2622 2752 2625 2848
rect 2638 2832 2641 2918
rect 2654 2871 2657 2918
rect 2670 2912 2673 2918
rect 2670 2892 2673 2898
rect 2654 2868 2665 2871
rect 2650 2858 2654 2861
rect 2662 2762 2665 2868
rect 2678 2862 2681 2868
rect 2670 2842 2673 2848
rect 2694 2762 2697 2918
rect 2710 2881 2713 2938
rect 2718 2892 2721 2958
rect 2710 2878 2721 2881
rect 2702 2832 2705 2858
rect 2710 2812 2713 2868
rect 2706 2758 2710 2761
rect 2598 2742 2601 2748
rect 2646 2742 2649 2748
rect 2694 2742 2697 2748
rect 2718 2742 2721 2878
rect 2726 2862 2729 2868
rect 2734 2852 2737 2948
rect 2750 2892 2753 2958
rect 2758 2952 2761 2978
rect 2766 2952 2769 2958
rect 2758 2942 2761 2948
rect 2758 2922 2761 2928
rect 2774 2892 2777 3048
rect 2754 2868 2758 2871
rect 2774 2852 2777 2868
rect 2730 2848 2734 2851
rect 2762 2848 2766 2851
rect 2782 2841 2785 3118
rect 2814 3082 2817 3188
rect 2830 3102 2833 3268
rect 2870 3262 2873 3268
rect 2846 3242 2849 3248
rect 2854 3212 2857 3248
rect 2838 3162 2841 3168
rect 2862 3162 2865 3218
rect 2878 3192 2881 3268
rect 2922 3248 2926 3251
rect 2894 3242 2897 3248
rect 2870 3141 2873 3148
rect 2886 3142 2889 3148
rect 2870 3138 2878 3141
rect 2838 3092 2841 3128
rect 2846 3122 2849 3128
rect 2862 3092 2865 3138
rect 2874 3128 2878 3131
rect 2886 3122 2889 3138
rect 2894 3111 2897 3238
rect 2902 3192 2905 3208
rect 2918 3162 2921 3168
rect 2934 3162 2937 3278
rect 2986 3268 2990 3271
rect 3058 3268 3062 3271
rect 2942 3262 2945 3268
rect 2966 3262 2969 3268
rect 2990 3252 2993 3258
rect 2946 3248 2950 3251
rect 2966 3162 2969 3208
rect 2990 3152 2993 3198
rect 3006 3192 3009 3248
rect 3014 3242 3017 3268
rect 3026 3248 3030 3251
rect 3038 3212 3041 3248
rect 3022 3162 3025 3168
rect 3070 3162 3073 3358
rect 3086 3342 3089 3348
rect 3078 3262 3081 3268
rect 3086 3262 3089 3338
rect 3094 3282 3097 3338
rect 3102 3292 3105 3418
rect 3118 3362 3121 3378
rect 3134 3362 3137 3418
rect 3166 3382 3169 3418
rect 3190 3362 3193 3388
rect 3154 3358 3158 3361
rect 3170 3358 3174 3361
rect 3110 3352 3113 3358
rect 3126 3322 3129 3328
rect 3098 3268 3102 3271
rect 3086 3242 3089 3258
rect 3110 3252 3113 3318
rect 3126 3292 3129 3308
rect 3134 3292 3137 3338
rect 3142 3312 3145 3338
rect 3158 3301 3161 3318
rect 3166 3312 3169 3318
rect 3182 3312 3185 3338
rect 3202 3328 3206 3331
rect 3158 3298 3169 3301
rect 3150 3272 3153 3278
rect 3134 3252 3137 3258
rect 3122 3248 3126 3251
rect 3102 3162 3105 3168
rect 3110 3162 3113 3208
rect 2938 3138 2942 3141
rect 3050 3138 3054 3141
rect 2886 3108 2897 3111
rect 2846 3082 2849 3088
rect 2854 3082 2857 3088
rect 2790 3042 2793 3058
rect 2790 2952 2793 3038
rect 2802 2958 2806 2961
rect 2790 2892 2793 2948
rect 2806 2932 2809 2938
rect 2814 2902 2817 3078
rect 2822 3032 2825 3068
rect 2878 3062 2881 3068
rect 2886 3052 2889 3108
rect 2894 3092 2897 3098
rect 2910 3072 2913 3078
rect 2898 3068 2902 3071
rect 2914 3058 2918 3061
rect 2910 3048 2918 3051
rect 2838 3042 2841 3048
rect 2862 3042 2865 3048
rect 2838 2972 2841 3028
rect 2886 2972 2889 2998
rect 2834 2938 2838 2941
rect 2774 2838 2785 2841
rect 2734 2772 2737 2838
rect 2774 2772 2777 2838
rect 2806 2832 2809 2858
rect 2814 2762 2817 2858
rect 2822 2772 2825 2928
rect 2838 2862 2841 2868
rect 2846 2852 2849 2918
rect 2862 2872 2865 2938
rect 2862 2862 2865 2868
rect 2838 2772 2841 2848
rect 2846 2762 2849 2768
rect 2766 2752 2769 2758
rect 2722 2738 2726 2741
rect 2738 2738 2742 2741
rect 2478 2702 2481 2718
rect 2482 2688 2486 2691
rect 2542 2672 2545 2718
rect 2574 2712 2577 2728
rect 2454 2572 2457 2659
rect 2518 2612 2521 2658
rect 2550 2652 2553 2659
rect 2544 2603 2546 2607
rect 2550 2603 2553 2607
rect 2557 2603 2560 2607
rect 2566 2602 2569 2658
rect 2582 2652 2585 2668
rect 2466 2558 2470 2561
rect 2466 2548 2470 2551
rect 2542 2551 2545 2588
rect 2590 2562 2593 2718
rect 2614 2712 2617 2718
rect 2622 2712 2625 2728
rect 2662 2702 2665 2718
rect 2670 2712 2673 2728
rect 2606 2672 2609 2678
rect 2630 2662 2633 2698
rect 2606 2552 2609 2558
rect 2662 2552 2665 2558
rect 2442 2538 2446 2541
rect 2358 2522 2361 2528
rect 2354 2488 2358 2491
rect 2390 2482 2393 2528
rect 2390 2452 2393 2459
rect 2422 2442 2425 2538
rect 2558 2532 2561 2538
rect 2510 2492 2513 2528
rect 2582 2481 2585 2518
rect 2630 2512 2633 2528
rect 2638 2512 2641 2528
rect 2578 2478 2585 2481
rect 2518 2472 2521 2478
rect 2590 2472 2593 2478
rect 2458 2468 2462 2471
rect 2578 2468 2582 2471
rect 2634 2468 2638 2471
rect 2502 2462 2505 2468
rect 2306 2358 2310 2361
rect 2254 2352 2257 2358
rect 2278 2342 2281 2348
rect 2318 2342 2321 2388
rect 2330 2358 2334 2361
rect 2342 2342 2345 2388
rect 2374 2362 2377 2368
rect 2410 2358 2414 2361
rect 2402 2348 2409 2351
rect 2394 2338 2398 2341
rect 2298 2328 2302 2331
rect 2362 2328 2366 2331
rect 2246 2312 2249 2318
rect 2262 2282 2265 2288
rect 2178 2248 2182 2251
rect 2158 2188 2169 2191
rect 2214 2192 2217 2268
rect 2242 2248 2246 2251
rect 1998 2132 2001 2138
rect 1986 2078 1990 2081
rect 2014 2063 2017 2118
rect 2024 2103 2026 2107
rect 2030 2103 2033 2107
rect 2037 2103 2040 2107
rect 2094 2072 2097 2118
rect 1986 2058 1990 2061
rect 2098 2058 2102 2061
rect 1830 2042 1833 2058
rect 1822 1992 1825 1998
rect 1758 1972 1761 1988
rect 1854 1982 1857 2018
rect 1774 1952 1777 1958
rect 1738 1948 1742 1951
rect 1798 1942 1801 1958
rect 1854 1952 1857 1968
rect 1726 1882 1729 1888
rect 1718 1851 1721 1868
rect 1710 1848 1721 1851
rect 1734 1852 1737 1938
rect 1766 1872 1769 1878
rect 1782 1872 1785 1938
rect 1794 1928 1798 1931
rect 1806 1872 1809 1878
rect 1746 1868 1750 1871
rect 1786 1868 1790 1871
rect 1798 1862 1801 1868
rect 1814 1862 1817 1948
rect 1834 1938 1838 1941
rect 1822 1932 1825 1938
rect 1746 1858 1750 1861
rect 1710 1732 1713 1848
rect 1758 1841 1761 1858
rect 1774 1852 1777 1858
rect 1738 1838 1761 1841
rect 1782 1812 1785 1858
rect 1814 1852 1817 1858
rect 1834 1849 1838 1851
rect 1834 1848 1841 1849
rect 1846 1832 1849 1948
rect 1862 1942 1865 2028
rect 1894 1972 1897 2008
rect 1894 1962 1897 1968
rect 1934 1952 1937 1968
rect 1874 1938 1878 1941
rect 1866 1928 1870 1931
rect 1886 1912 1889 1948
rect 1906 1938 1910 1941
rect 1938 1938 1942 1941
rect 1886 1882 1889 1888
rect 1870 1862 1873 1878
rect 1858 1858 1862 1861
rect 1718 1752 1721 1768
rect 1726 1732 1729 1788
rect 1758 1772 1761 1798
rect 1742 1762 1745 1768
rect 1738 1748 1750 1751
rect 1786 1748 1790 1751
rect 1774 1732 1777 1738
rect 1798 1732 1801 1748
rect 1822 1742 1825 1768
rect 1830 1732 1833 1748
rect 1854 1732 1857 1768
rect 1878 1732 1881 1868
rect 1886 1772 1889 1878
rect 1894 1862 1897 1918
rect 1918 1882 1921 1918
rect 1934 1892 1937 1928
rect 1918 1862 1921 1868
rect 1898 1848 1902 1851
rect 1910 1792 1913 1818
rect 1926 1812 1929 1848
rect 1934 1801 1937 1878
rect 1942 1872 1945 1918
rect 1950 1902 1953 2018
rect 2046 1992 2049 2038
rect 2054 2012 2057 2018
rect 2102 2002 2105 2058
rect 2086 1972 2089 1978
rect 2002 1968 2006 1971
rect 1958 1952 1961 1968
rect 2062 1962 2065 1968
rect 1974 1882 1977 1918
rect 1982 1912 1985 1958
rect 2050 1948 2054 1951
rect 2006 1941 2009 1948
rect 2002 1938 2009 1941
rect 2070 1942 2073 1958
rect 2090 1948 2094 1951
rect 1998 1922 2001 1938
rect 2110 1932 2113 2168
rect 2158 2151 2161 2188
rect 2230 2182 2233 2248
rect 2254 2182 2257 2248
rect 2126 2082 2129 2148
rect 2190 2142 2193 2178
rect 2222 2162 2225 2178
rect 2246 2162 2249 2178
rect 2206 2152 2209 2158
rect 2270 2152 2273 2158
rect 2226 2148 2230 2151
rect 2278 2142 2281 2268
rect 2302 2252 2305 2318
rect 2326 2262 2329 2288
rect 2334 2281 2337 2318
rect 2350 2302 2353 2318
rect 2406 2312 2409 2348
rect 2422 2342 2425 2438
rect 2454 2382 2457 2418
rect 2478 2362 2481 2448
rect 2474 2348 2481 2351
rect 2446 2342 2449 2348
rect 2450 2338 2454 2341
rect 2466 2328 2470 2331
rect 2394 2288 2398 2291
rect 2334 2278 2345 2281
rect 2334 2262 2337 2268
rect 2342 2252 2345 2278
rect 2382 2272 2385 2278
rect 2362 2268 2366 2271
rect 2398 2252 2401 2278
rect 2406 2262 2409 2308
rect 2310 2242 2313 2248
rect 2478 2232 2481 2348
rect 2510 2342 2513 2468
rect 2578 2458 2582 2461
rect 2530 2448 2534 2451
rect 2602 2448 2606 2451
rect 2638 2442 2641 2458
rect 2544 2403 2546 2407
rect 2550 2403 2553 2407
rect 2557 2403 2560 2407
rect 2582 2351 2585 2358
rect 2654 2352 2657 2528
rect 2670 2482 2673 2648
rect 2678 2562 2681 2708
rect 2702 2662 2705 2738
rect 2726 2712 2729 2718
rect 2718 2652 2721 2668
rect 2726 2662 2729 2668
rect 2686 2572 2689 2618
rect 2750 2582 2753 2678
rect 2766 2632 2769 2748
rect 2802 2738 2806 2741
rect 2826 2738 2830 2741
rect 2810 2718 2814 2721
rect 2758 2572 2761 2578
rect 2746 2548 2750 2551
rect 2682 2538 2686 2541
rect 2742 2532 2745 2548
rect 2678 2462 2681 2518
rect 2750 2492 2753 2528
rect 2774 2491 2777 2718
rect 2830 2702 2833 2718
rect 2846 2682 2849 2718
rect 2854 2663 2857 2858
rect 2862 2752 2865 2858
rect 2870 2772 2873 2918
rect 2886 2912 2889 2928
rect 2886 2882 2889 2898
rect 2902 2892 2905 3028
rect 2910 2992 2913 3048
rect 2926 3041 2929 3128
rect 2934 3092 2937 3128
rect 2942 3062 2945 3118
rect 2918 3038 2929 3041
rect 2910 2952 2913 2958
rect 2910 2872 2913 2948
rect 2886 2782 2889 2868
rect 2910 2852 2913 2868
rect 2918 2772 2921 3038
rect 2934 3032 2937 3048
rect 2950 2972 2953 3128
rect 2974 3092 2977 3138
rect 2982 3132 2985 3138
rect 3014 3092 3017 3138
rect 3030 3102 3033 3128
rect 3030 3082 3033 3088
rect 3038 3072 3041 3138
rect 3086 3122 3089 3138
rect 3048 3103 3050 3107
rect 3054 3103 3057 3107
rect 3061 3103 3064 3107
rect 2974 3052 2977 3068
rect 2974 3042 2977 3048
rect 2974 2962 2977 3038
rect 2930 2958 2934 2961
rect 2982 2942 2985 2948
rect 2958 2922 2961 2938
rect 2958 2872 2961 2908
rect 2966 2882 2969 2918
rect 2946 2858 2950 2861
rect 2926 2792 2929 2848
rect 2942 2832 2945 2858
rect 2950 2842 2953 2848
rect 2966 2772 2969 2858
rect 2974 2852 2977 2938
rect 2982 2872 2985 2878
rect 2982 2842 2985 2868
rect 2990 2841 2993 3068
rect 2998 3062 3001 3068
rect 3022 3062 3025 3068
rect 3010 3048 3014 3051
rect 3034 3048 3038 3051
rect 3014 3042 3017 3048
rect 3046 3042 3049 3048
rect 3022 2962 3025 2968
rect 3030 2962 3033 3038
rect 3038 2942 3041 3028
rect 3054 2972 3057 3088
rect 3070 3082 3073 3118
rect 3094 3092 3097 3108
rect 3082 3068 3086 3071
rect 3062 3062 3065 3068
rect 3094 2972 3097 3078
rect 3102 2992 3105 3118
rect 3110 3062 3113 3068
rect 3118 3051 3121 3248
rect 3134 3212 3137 3248
rect 3158 3212 3161 3268
rect 3150 3162 3153 3168
rect 3158 3162 3161 3178
rect 3166 3172 3169 3298
rect 3178 3268 3182 3271
rect 3214 3262 3217 3358
rect 3222 3302 3225 3418
rect 3230 3342 3233 3428
rect 3286 3362 3289 3418
rect 3310 3362 3313 3408
rect 3298 3358 3302 3361
rect 3326 3361 3329 3418
rect 3350 3362 3353 3418
rect 3398 3402 3401 3468
rect 3414 3452 3417 3468
rect 3430 3432 3433 3468
rect 3358 3362 3361 3368
rect 3326 3358 3337 3361
rect 3238 3352 3241 3358
rect 3274 3348 3278 3351
rect 3310 3348 3326 3351
rect 3262 3342 3265 3348
rect 3310 3342 3313 3348
rect 3322 3338 3326 3341
rect 3246 3322 3249 3328
rect 3230 3292 3233 3308
rect 3254 3292 3257 3338
rect 3174 3242 3177 3248
rect 3198 3242 3201 3258
rect 3214 3192 3217 3248
rect 3222 3222 3225 3278
rect 3246 3272 3249 3278
rect 3230 3252 3233 3258
rect 3254 3252 3257 3258
rect 3222 3192 3225 3218
rect 3182 3162 3185 3178
rect 3126 3092 3129 3138
rect 3134 3128 3142 3131
rect 3114 3048 3126 3051
rect 3118 2972 3121 3038
rect 3134 2972 3137 3128
rect 3166 3122 3169 3128
rect 3174 3092 3177 3138
rect 3186 3128 3190 3131
rect 3198 3092 3201 3138
rect 3214 3082 3217 3118
rect 3222 3092 3225 3178
rect 3230 3152 3233 3198
rect 3254 3162 3257 3168
rect 3238 3152 3241 3158
rect 3254 3142 3257 3148
rect 3158 3072 3161 3078
rect 3174 3052 3177 3078
rect 3202 3068 3206 3071
rect 3214 3071 3217 3078
rect 3230 3072 3233 3088
rect 3214 3068 3225 3071
rect 3182 3062 3185 3068
rect 3206 3058 3214 3061
rect 3146 3048 3150 3051
rect 3194 3048 3198 3051
rect 3142 3002 3145 3018
rect 3182 2972 3185 3048
rect 3206 2972 3209 3058
rect 3222 3052 3225 3068
rect 3230 2992 3233 3068
rect 3238 3062 3241 3118
rect 3246 3092 3249 3138
rect 3254 3052 3257 3118
rect 3242 3048 3246 3051
rect 3262 2972 3265 3328
rect 3286 3292 3289 3338
rect 3322 3328 3326 3331
rect 3302 3302 3305 3318
rect 3310 3292 3313 3318
rect 3334 3301 3337 3358
rect 3366 3352 3369 3368
rect 3406 3362 3409 3388
rect 3398 3352 3401 3358
rect 3374 3342 3377 3348
rect 3406 3342 3409 3358
rect 3430 3342 3433 3348
rect 3326 3298 3337 3301
rect 3298 3268 3302 3271
rect 3278 3262 3281 3268
rect 3290 3248 3294 3251
rect 3314 3248 3318 3251
rect 3278 3162 3281 3168
rect 3326 3162 3329 3298
rect 3342 3291 3345 3338
rect 3350 3322 3353 3328
rect 3338 3288 3345 3291
rect 3342 3272 3345 3278
rect 3350 3252 3353 3278
rect 3358 3162 3361 3318
rect 3366 3262 3369 3338
rect 3366 3232 3369 3258
rect 3374 3152 3377 3338
rect 3382 3332 3385 3338
rect 3390 3282 3393 3288
rect 3286 3142 3289 3148
rect 3302 3142 3305 3148
rect 3350 3142 3353 3148
rect 3362 3138 3366 3141
rect 3310 3132 3313 3138
rect 3270 3092 3273 3118
rect 3294 3112 3297 3118
rect 3286 3082 3289 3098
rect 3274 3068 3278 3071
rect 3294 3062 3297 3068
rect 3326 3062 3329 3078
rect 3270 3042 3273 3048
rect 3270 2972 3273 2988
rect 3286 2972 3289 2998
rect 3090 2938 3094 2941
rect 3122 2938 3134 2941
rect 3170 2938 3174 2941
rect 2998 2932 3001 2938
rect 3006 2932 3009 2938
rect 3030 2932 3033 2938
rect 3014 2872 3017 2928
rect 3002 2848 3006 2851
rect 2990 2838 3001 2841
rect 2934 2762 2937 2768
rect 2946 2758 2953 2761
rect 2938 2748 2942 2751
rect 2862 2742 2865 2748
rect 2890 2738 2894 2741
rect 2886 2712 2889 2728
rect 2902 2672 2905 2718
rect 2822 2652 2825 2658
rect 2886 2652 2889 2668
rect 2906 2658 2910 2661
rect 2790 2542 2793 2548
rect 2774 2488 2785 2491
rect 2758 2472 2761 2478
rect 2774 2472 2777 2478
rect 2678 2351 2681 2418
rect 2710 2352 2713 2358
rect 2598 2342 2601 2348
rect 2490 2338 2494 2341
rect 2530 2338 2534 2341
rect 2518 2272 2521 2288
rect 2534 2282 2537 2298
rect 2566 2292 2569 2338
rect 2650 2328 2654 2331
rect 2714 2318 2718 2321
rect 2502 2263 2505 2268
rect 2366 2162 2369 2178
rect 2314 2158 2318 2161
rect 2370 2158 2374 2161
rect 2286 2152 2289 2158
rect 2326 2152 2329 2158
rect 2398 2152 2401 2178
rect 2422 2162 2425 2218
rect 2430 2152 2433 2228
rect 2438 2192 2441 2218
rect 2454 2162 2457 2168
rect 2438 2152 2441 2158
rect 2306 2148 2310 2151
rect 2350 2142 2353 2148
rect 2454 2142 2457 2148
rect 2462 2142 2465 2148
rect 2510 2142 2513 2218
rect 2534 2212 2537 2278
rect 2544 2203 2546 2207
rect 2550 2203 2553 2207
rect 2557 2203 2560 2207
rect 2566 2152 2569 2288
rect 2614 2272 2617 2318
rect 2630 2282 2633 2288
rect 2630 2262 2633 2268
rect 2594 2258 2598 2261
rect 2574 2252 2577 2258
rect 2614 2252 2617 2258
rect 2602 2248 2606 2251
rect 2606 2222 2609 2228
rect 2606 2212 2609 2218
rect 2598 2151 2601 2158
rect 2630 2152 2633 2208
rect 2638 2142 2641 2258
rect 2654 2232 2657 2278
rect 2666 2268 2670 2271
rect 2678 2252 2681 2288
rect 2686 2272 2689 2298
rect 2726 2292 2729 2468
rect 2758 2452 2761 2458
rect 2738 2448 2742 2451
rect 2774 2392 2777 2468
rect 2782 2452 2785 2488
rect 2790 2462 2793 2468
rect 2798 2462 2801 2548
rect 2806 2482 2809 2648
rect 2822 2551 2825 2568
rect 2838 2512 2841 2648
rect 2858 2568 2870 2571
rect 2858 2558 2862 2561
rect 2874 2548 2878 2551
rect 2822 2482 2825 2498
rect 2854 2482 2857 2508
rect 2878 2482 2881 2538
rect 2758 2362 2761 2368
rect 2782 2352 2785 2358
rect 2754 2348 2758 2351
rect 2734 2342 2737 2348
rect 2798 2342 2801 2388
rect 2806 2362 2809 2478
rect 2854 2452 2857 2459
rect 2902 2422 2905 2618
rect 2910 2552 2913 2658
rect 2918 2652 2921 2738
rect 2926 2682 2929 2698
rect 2950 2692 2953 2758
rect 2958 2752 2961 2768
rect 2858 2358 2862 2361
rect 2814 2352 2817 2358
rect 2834 2348 2838 2351
rect 2746 2338 2750 2341
rect 2838 2322 2841 2338
rect 2742 2312 2745 2318
rect 2766 2292 2769 2308
rect 2754 2278 2758 2281
rect 2734 2262 2737 2268
rect 2682 2248 2686 2251
rect 2706 2248 2710 2251
rect 2758 2242 2761 2268
rect 2774 2252 2777 2298
rect 2782 2272 2785 2278
rect 2806 2262 2809 2318
rect 2818 2278 2822 2281
rect 2838 2262 2841 2318
rect 2854 2302 2857 2358
rect 2870 2352 2873 2368
rect 2878 2342 2881 2398
rect 2898 2358 2902 2361
rect 2898 2348 2902 2351
rect 2862 2291 2865 2298
rect 2858 2288 2865 2291
rect 2890 2278 2894 2281
rect 2810 2258 2822 2261
rect 2786 2248 2790 2251
rect 2862 2242 2865 2268
rect 2894 2262 2897 2268
rect 2874 2258 2878 2261
rect 2882 2258 2886 2261
rect 2882 2248 2886 2251
rect 2886 2242 2889 2248
rect 2810 2238 2814 2241
rect 2758 2232 2761 2238
rect 2670 2162 2673 2218
rect 2658 2158 2662 2161
rect 2690 2158 2694 2161
rect 2682 2148 2686 2151
rect 2654 2142 2657 2148
rect 2202 2138 2206 2141
rect 2282 2138 2286 2141
rect 2314 2138 2318 2141
rect 2402 2138 2406 2141
rect 2682 2138 2686 2141
rect 2714 2138 2718 2141
rect 2230 2122 2233 2138
rect 2162 2078 2166 2081
rect 2170 2078 2177 2081
rect 2174 2072 2177 2078
rect 2222 2072 2225 2078
rect 2122 2059 2126 2062
rect 2162 2048 2166 2051
rect 2202 2048 2206 2051
rect 2190 2041 2193 2048
rect 2222 2041 2225 2058
rect 2190 2038 2225 2041
rect 2118 1942 2121 1958
rect 2154 1948 2158 1951
rect 2134 1942 2137 1948
rect 2010 1928 2014 1931
rect 2110 1922 2113 1928
rect 2024 1903 2026 1907
rect 2030 1903 2033 1907
rect 2037 1903 2040 1907
rect 2142 1902 2145 1918
rect 2158 1912 2161 1948
rect 2182 1932 2185 1938
rect 1926 1798 1937 1801
rect 1898 1768 1902 1771
rect 1926 1762 1929 1798
rect 1942 1792 1945 1828
rect 1934 1772 1937 1788
rect 1950 1762 1953 1878
rect 1962 1788 1966 1791
rect 1898 1748 1926 1751
rect 1882 1728 1886 1731
rect 1694 1672 1697 1688
rect 1702 1672 1705 1698
rect 1718 1672 1721 1728
rect 1758 1672 1761 1718
rect 1486 1542 1489 1548
rect 1466 1528 1470 1531
rect 1494 1522 1497 1558
rect 1514 1538 1518 1541
rect 1462 1462 1465 1468
rect 1470 1462 1473 1518
rect 1502 1502 1505 1518
rect 1478 1441 1481 1498
rect 1518 1472 1521 1538
rect 1534 1532 1537 1568
rect 1550 1542 1553 1568
rect 1574 1562 1577 1568
rect 1558 1532 1561 1548
rect 1606 1542 1609 1598
rect 1614 1552 1617 1608
rect 1638 1602 1641 1668
rect 1658 1638 1662 1641
rect 1638 1552 1641 1558
rect 1658 1548 1662 1551
rect 1606 1532 1609 1538
rect 1546 1528 1550 1531
rect 1538 1478 1542 1481
rect 1506 1468 1510 1471
rect 1486 1462 1489 1468
rect 1530 1458 1534 1461
rect 1474 1438 1481 1441
rect 1486 1422 1489 1448
rect 1550 1422 1553 1468
rect 1558 1462 1561 1468
rect 1566 1462 1569 1518
rect 1582 1472 1585 1498
rect 1606 1492 1609 1508
rect 1622 1472 1625 1498
rect 1410 1338 1414 1341
rect 1290 1328 1297 1331
rect 1314 1328 1318 1331
rect 1286 1272 1289 1278
rect 1286 1262 1289 1268
rect 1230 1252 1233 1258
rect 1294 1222 1297 1328
rect 1306 1318 1310 1321
rect 1366 1281 1369 1338
rect 1418 1328 1422 1331
rect 1358 1278 1369 1281
rect 1302 1262 1305 1278
rect 1310 1252 1313 1258
rect 1322 1238 1326 1241
rect 1326 1202 1329 1218
rect 1334 1172 1337 1278
rect 1358 1272 1361 1278
rect 1178 1168 1182 1171
rect 1266 1168 1270 1171
rect 1086 1162 1089 1168
rect 1118 1162 1121 1168
rect 1066 1158 1070 1161
rect 1098 1158 1102 1161
rect 1058 1148 1062 1151
rect 1082 1148 1086 1151
rect 1066 1138 1070 1141
rect 1098 1138 1102 1141
rect 990 1068 998 1071
rect 1022 1070 1025 1078
rect 986 1058 990 1061
rect 998 1052 1001 1068
rect 1030 1032 1033 1138
rect 1118 1132 1121 1138
rect 1126 1122 1129 1158
rect 1138 1148 1142 1151
rect 1158 1142 1161 1158
rect 1206 1142 1209 1148
rect 1230 1142 1233 1158
rect 1298 1148 1302 1151
rect 1146 1138 1150 1141
rect 1218 1138 1222 1141
rect 1238 1132 1241 1148
rect 1246 1142 1249 1148
rect 1318 1142 1321 1148
rect 1294 1132 1297 1138
rect 1038 1092 1041 1118
rect 1214 1112 1217 1128
rect 1302 1121 1305 1128
rect 1294 1118 1305 1121
rect 1050 1088 1054 1091
rect 1062 1072 1065 1078
rect 1070 1072 1073 1078
rect 1118 1072 1121 1098
rect 1138 1088 1142 1091
rect 1126 1082 1129 1088
rect 1158 1082 1161 1098
rect 1174 1072 1177 1078
rect 1190 1072 1193 1078
rect 1218 1068 1222 1071
rect 1042 1048 1046 1051
rect 1142 1032 1145 1068
rect 1230 1062 1233 1118
rect 1194 1058 1198 1061
rect 974 1002 977 1018
rect 1062 992 1065 1028
rect 1090 1018 1094 1021
rect 1018 958 1022 961
rect 950 952 953 958
rect 974 952 977 958
rect 922 948 926 951
rect 954 938 958 941
rect 994 938 998 941
rect 878 932 881 938
rect 990 932 993 938
rect 878 892 881 918
rect 886 872 889 918
rect 934 872 937 878
rect 950 872 953 898
rect 746 868 750 871
rect 694 862 697 868
rect 726 862 729 868
rect 966 863 969 888
rect 714 858 718 861
rect 818 859 822 862
rect 702 842 705 848
rect 734 842 737 848
rect 694 832 697 838
rect 726 832 729 838
rect 758 812 761 818
rect 630 752 633 768
rect 638 752 641 758
rect 646 752 649 808
rect 678 762 681 768
rect 774 762 777 818
rect 910 812 913 818
rect 702 752 705 758
rect 674 748 678 751
rect 622 741 625 748
rect 622 738 633 741
rect 698 738 702 741
rect 630 692 633 738
rect 574 618 585 621
rect 454 552 457 588
rect 574 542 577 618
rect 638 562 641 708
rect 662 702 665 718
rect 658 688 662 691
rect 654 652 657 678
rect 670 662 673 688
rect 710 682 713 758
rect 750 752 753 758
rect 870 752 873 808
rect 950 752 953 858
rect 974 852 977 928
rect 982 892 985 918
rect 1000 903 1002 907
rect 1006 903 1009 907
rect 1013 903 1016 907
rect 1030 872 1033 918
rect 1038 842 1041 928
rect 1046 892 1049 968
rect 1074 958 1078 961
rect 1054 902 1057 948
rect 1078 942 1081 948
rect 1126 942 1129 978
rect 1150 962 1153 1058
rect 1174 1052 1177 1058
rect 1214 1022 1217 1048
rect 1182 962 1185 1018
rect 1198 1002 1201 1018
rect 1138 958 1142 961
rect 1054 872 1057 898
rect 1102 822 1105 918
rect 1118 892 1121 898
rect 1134 882 1137 918
rect 1150 902 1153 958
rect 1166 952 1169 958
rect 1158 942 1161 948
rect 1214 942 1217 958
rect 1222 942 1225 948
rect 1230 942 1233 1018
rect 1238 952 1241 1108
rect 1294 1092 1297 1118
rect 1302 1092 1305 1098
rect 1334 1092 1337 1138
rect 1342 1112 1345 1258
rect 1358 1252 1361 1258
rect 1366 1251 1369 1268
rect 1374 1262 1377 1298
rect 1366 1248 1374 1251
rect 1354 1158 1358 1161
rect 1354 1148 1358 1151
rect 1358 1122 1361 1128
rect 1262 1082 1265 1088
rect 1358 1082 1361 1088
rect 1314 1068 1318 1071
rect 1270 1052 1273 1068
rect 1270 962 1273 1048
rect 1278 1022 1281 1058
rect 1294 1052 1297 1058
rect 1302 1042 1305 1048
rect 1142 882 1145 888
rect 1146 868 1150 871
rect 1110 862 1113 868
rect 1078 802 1081 818
rect 734 742 737 748
rect 754 738 758 741
rect 746 718 750 721
rect 678 662 681 668
rect 702 662 705 668
rect 710 662 713 678
rect 754 658 758 661
rect 670 641 673 658
rect 730 648 734 651
rect 670 638 681 641
rect 670 632 673 638
rect 650 628 654 631
rect 654 592 657 598
rect 654 582 657 588
rect 662 562 665 568
rect 486 492 489 518
rect 510 512 513 538
rect 574 532 577 538
rect 534 482 537 532
rect 590 512 593 547
rect 542 492 545 508
rect 558 492 561 508
rect 390 472 393 478
rect 478 472 481 478
rect 534 472 537 478
rect 558 472 561 488
rect 626 478 630 481
rect 638 472 641 558
rect 678 544 681 638
rect 686 542 689 648
rect 750 642 753 648
rect 742 632 745 638
rect 742 562 745 608
rect 758 602 761 658
rect 694 552 697 558
rect 734 552 737 558
rect 746 548 750 551
rect 670 472 673 488
rect 366 462 369 468
rect 354 438 358 441
rect 326 402 329 418
rect 286 392 289 398
rect 350 392 353 428
rect 374 422 377 448
rect 406 432 409 459
rect 478 442 481 468
rect 326 372 329 378
rect 354 368 358 371
rect 270 342 273 348
rect 258 338 262 341
rect 174 332 177 338
rect 198 332 201 338
rect 150 262 153 318
rect 166 312 169 328
rect 206 302 209 318
rect 214 312 217 328
rect 294 292 297 348
rect 302 302 305 358
rect 310 342 313 368
rect 342 352 345 358
rect 366 352 369 418
rect 374 362 377 398
rect 406 352 409 388
rect 322 348 326 351
rect 402 338 406 341
rect 158 272 161 278
rect 214 272 217 278
rect 286 272 289 278
rect 238 268 262 271
rect 206 262 209 268
rect 238 262 241 268
rect 294 262 297 268
rect 302 262 305 298
rect 310 272 313 298
rect 318 282 321 338
rect 386 328 390 331
rect 402 318 406 321
rect 326 292 329 308
rect 374 272 377 278
rect 10 118 14 121
rect 22 62 25 118
rect 38 92 41 148
rect 54 122 57 259
rect 130 258 134 261
rect 162 258 166 261
rect 266 258 270 261
rect 246 252 249 258
rect 310 252 313 258
rect 186 248 190 251
rect 122 238 126 241
rect 70 151 73 198
rect 150 192 153 218
rect 98 188 102 191
rect 86 142 89 148
rect 134 142 137 148
rect 94 72 97 78
rect 134 72 137 138
rect 118 62 121 68
rect 150 63 153 188
rect 198 162 201 248
rect 238 242 241 248
rect 274 238 278 241
rect 230 232 233 238
rect 210 228 214 231
rect 222 202 225 218
rect 166 151 169 158
rect 182 72 185 78
rect 198 62 201 158
rect 206 152 209 178
rect 238 172 241 178
rect 246 172 249 238
rect 318 222 321 268
rect 382 262 385 298
rect 354 258 358 261
rect 370 248 374 251
rect 334 232 337 248
rect 354 238 358 241
rect 218 168 222 171
rect 222 152 225 158
rect 238 152 241 158
rect 230 92 233 148
rect 262 142 265 178
rect 294 172 297 218
rect 218 88 222 91
rect 262 82 265 138
rect 278 62 281 68
rect 310 63 313 208
rect 342 172 345 238
rect 358 202 361 218
rect 366 162 369 188
rect 382 172 385 218
rect 390 182 393 288
rect 406 272 409 298
rect 406 252 409 258
rect 422 252 425 368
rect 462 352 465 388
rect 474 358 478 361
rect 486 352 489 408
rect 496 403 498 407
rect 502 403 505 407
rect 509 403 512 407
rect 518 362 521 458
rect 558 382 561 468
rect 566 462 569 468
rect 570 458 577 461
rect 610 458 622 461
rect 574 371 577 458
rect 622 452 625 458
rect 638 452 641 468
rect 646 452 649 458
rect 610 448 614 451
rect 582 442 585 448
rect 594 438 598 441
rect 590 392 593 418
rect 606 392 609 418
rect 574 368 582 371
rect 574 352 577 368
rect 590 352 593 378
rect 622 372 625 418
rect 474 348 478 351
rect 554 348 558 351
rect 442 328 446 331
rect 454 292 457 318
rect 430 262 433 268
rect 454 262 457 268
rect 422 212 425 248
rect 462 202 465 248
rect 390 162 393 168
rect 350 152 353 158
rect 370 148 374 151
rect 422 151 425 158
rect 326 142 329 148
rect 342 142 345 148
rect 358 92 361 148
rect 406 142 409 148
rect 406 82 409 138
rect 470 111 473 328
rect 486 302 489 348
rect 566 342 569 348
rect 542 312 545 338
rect 502 282 505 288
rect 490 278 494 281
rect 478 272 481 278
rect 482 258 486 261
rect 494 252 497 278
rect 502 262 505 278
rect 496 203 498 207
rect 502 203 505 207
rect 509 203 512 207
rect 510 152 513 168
rect 526 142 529 278
rect 542 272 545 278
rect 542 222 545 268
rect 558 262 561 318
rect 566 312 569 328
rect 550 252 553 258
rect 558 242 561 258
rect 534 202 537 218
rect 562 178 566 181
rect 574 172 577 348
rect 590 332 593 348
rect 598 322 601 358
rect 582 282 585 288
rect 590 272 593 278
rect 602 258 606 261
rect 614 252 617 328
rect 622 272 625 278
rect 638 272 641 378
rect 646 342 649 348
rect 662 322 665 458
rect 670 442 673 468
rect 678 462 681 540
rect 686 452 689 538
rect 710 492 713 528
rect 718 492 721 548
rect 730 478 734 481
rect 746 468 750 471
rect 766 471 769 718
rect 782 572 785 718
rect 782 552 785 558
rect 790 551 793 698
rect 806 662 809 678
rect 830 662 833 688
rect 926 672 929 728
rect 958 692 961 788
rect 1158 772 1161 938
rect 1166 932 1169 938
rect 1230 931 1233 938
rect 1226 928 1233 931
rect 1190 912 1193 918
rect 1214 892 1217 898
rect 1182 882 1185 888
rect 1238 881 1241 948
rect 1250 928 1254 931
rect 1262 892 1265 948
rect 1270 892 1273 918
rect 1278 902 1281 958
rect 1286 922 1289 928
rect 1250 888 1254 891
rect 1238 878 1249 881
rect 1166 872 1169 878
rect 1206 872 1209 878
rect 1246 872 1249 878
rect 1286 872 1289 878
rect 1294 872 1297 938
rect 1302 872 1305 1028
rect 1318 961 1321 1058
rect 1326 1052 1329 1078
rect 1366 1071 1369 1188
rect 1374 1172 1377 1218
rect 1382 1142 1385 1318
rect 1398 1312 1401 1318
rect 1414 1292 1417 1298
rect 1406 1272 1409 1278
rect 1422 1272 1425 1298
rect 1398 1262 1401 1268
rect 1394 1248 1398 1251
rect 1430 1192 1433 1348
rect 1462 1342 1465 1418
rect 1520 1403 1522 1407
rect 1526 1403 1529 1407
rect 1533 1403 1536 1407
rect 1446 1312 1449 1338
rect 1454 1272 1457 1298
rect 1462 1272 1465 1328
rect 1438 1182 1441 1248
rect 1450 1238 1454 1241
rect 1462 1232 1465 1268
rect 1470 1252 1473 1368
rect 1494 1362 1497 1368
rect 1486 1358 1494 1361
rect 1486 1292 1489 1358
rect 1542 1352 1545 1358
rect 1506 1348 1510 1351
rect 1494 1342 1497 1348
rect 1550 1342 1553 1368
rect 1486 1282 1489 1288
rect 1486 1252 1489 1258
rect 1470 1162 1473 1248
rect 1478 1232 1481 1248
rect 1502 1212 1505 1338
rect 1518 1322 1521 1338
rect 1510 1252 1513 1258
rect 1534 1251 1537 1258
rect 1542 1252 1545 1338
rect 1534 1248 1542 1251
rect 1522 1238 1526 1241
rect 1478 1162 1481 1168
rect 1494 1162 1497 1198
rect 1502 1162 1505 1208
rect 1398 1152 1401 1158
rect 1402 1148 1406 1151
rect 1386 1138 1390 1141
rect 1414 1132 1417 1138
rect 1382 1082 1385 1118
rect 1422 1102 1425 1148
rect 1430 1142 1433 1148
rect 1438 1132 1441 1158
rect 1454 1152 1457 1158
rect 1494 1142 1497 1158
rect 1510 1141 1513 1218
rect 1520 1203 1522 1207
rect 1526 1203 1529 1207
rect 1533 1203 1536 1207
rect 1542 1142 1545 1158
rect 1550 1152 1553 1338
rect 1558 1332 1561 1458
rect 1566 1452 1569 1458
rect 1578 1438 1582 1441
rect 1590 1382 1593 1458
rect 1598 1422 1601 1468
rect 1630 1462 1633 1518
rect 1626 1448 1630 1451
rect 1638 1432 1641 1548
rect 1670 1542 1673 1568
rect 1686 1551 1689 1658
rect 1718 1642 1721 1668
rect 1750 1662 1753 1668
rect 1782 1662 1785 1718
rect 1790 1682 1793 1728
rect 1894 1722 1897 1738
rect 1950 1732 1953 1758
rect 1974 1742 1977 1868
rect 1982 1862 1985 1888
rect 2066 1878 2070 1881
rect 1994 1858 1998 1861
rect 2018 1858 2022 1861
rect 2054 1752 2057 1878
rect 2078 1872 2081 1888
rect 2182 1882 2185 1908
rect 2198 1892 2201 1978
rect 2214 1942 2217 1998
rect 2230 1952 2233 2098
rect 2246 2082 2249 2138
rect 2278 2072 2281 2128
rect 2326 2122 2329 2128
rect 2294 2082 2297 2088
rect 2342 2082 2345 2128
rect 2298 2068 2302 2071
rect 2330 2068 2334 2071
rect 2278 2062 2281 2068
rect 2254 2031 2257 2038
rect 2250 2028 2257 2031
rect 2274 2028 2278 2031
rect 2286 1962 2289 1998
rect 2290 1948 2294 1951
rect 2302 1951 2305 2068
rect 2350 2062 2353 2088
rect 2366 2082 2369 2128
rect 2318 2052 2321 2058
rect 2310 1982 2313 2018
rect 2302 1948 2313 1951
rect 2278 1932 2281 1938
rect 2302 1882 2305 1938
rect 2310 1932 2313 1948
rect 2318 1942 2321 2048
rect 2326 2032 2329 2048
rect 2350 1992 2353 2028
rect 2342 1952 2345 1978
rect 2310 1892 2313 1928
rect 2338 1878 2342 1881
rect 2102 1872 2105 1878
rect 2062 1852 2065 1868
rect 2122 1858 2126 1861
rect 1970 1738 1974 1741
rect 2006 1732 2009 1748
rect 2070 1742 2073 1758
rect 2078 1752 2081 1858
rect 2134 1812 2137 1878
rect 2182 1872 2185 1878
rect 2206 1872 2209 1878
rect 2142 1862 2145 1868
rect 2230 1862 2233 1868
rect 2214 1852 2217 1858
rect 2186 1848 2190 1851
rect 2166 1842 2169 1848
rect 2174 1842 2177 1848
rect 2230 1842 2233 1848
rect 2238 1812 2241 1868
rect 2254 1852 2257 1858
rect 2294 1852 2297 1858
rect 2302 1852 2305 1878
rect 2350 1862 2353 1978
rect 2382 1962 2385 2118
rect 2446 2092 2449 2118
rect 2462 2092 2465 2138
rect 2478 2132 2482 2135
rect 2734 2132 2737 2158
rect 2390 2082 2393 2088
rect 2478 2072 2481 2118
rect 2534 2112 2537 2118
rect 2490 2088 2494 2091
rect 2418 2068 2422 2071
rect 2466 2068 2470 2071
rect 2486 2068 2510 2071
rect 2522 2068 2526 2071
rect 2418 2058 2422 2061
rect 2442 2058 2446 2061
rect 2406 2052 2409 2058
rect 2462 2052 2465 2068
rect 2486 2062 2489 2068
rect 2522 2058 2526 2061
rect 2478 2052 2481 2058
rect 2490 2048 2494 2051
rect 2438 2032 2441 2038
rect 2450 1958 2454 1961
rect 2382 1952 2385 1958
rect 2470 1952 2473 1958
rect 2390 1948 2398 1951
rect 2374 1941 2377 1948
rect 2390 1941 2393 1948
rect 2422 1942 2425 1948
rect 2374 1938 2393 1941
rect 2398 1932 2401 1938
rect 2426 1928 2430 1931
rect 2398 1882 2401 1908
rect 2410 1878 2414 1881
rect 2422 1872 2425 1918
rect 2454 1912 2457 1938
rect 2462 1922 2465 1928
rect 2470 1912 2473 1928
rect 2478 1882 2481 1988
rect 2494 1942 2497 1948
rect 2494 1882 2497 1908
rect 2502 1892 2505 2058
rect 2526 1992 2529 2048
rect 2534 1992 2537 2108
rect 2742 2102 2745 2158
rect 2582 2092 2585 2098
rect 2590 2072 2593 2078
rect 2598 2072 2601 2078
rect 2606 2072 2609 2078
rect 2678 2072 2681 2088
rect 2734 2082 2737 2088
rect 2698 2078 2702 2081
rect 2750 2072 2753 2228
rect 2758 2192 2761 2208
rect 2838 2162 2841 2228
rect 2910 2222 2913 2468
rect 2918 2402 2921 2648
rect 2934 2642 2937 2668
rect 2950 2662 2953 2668
rect 2974 2661 2977 2758
rect 2990 2732 2993 2738
rect 2982 2692 2985 2728
rect 2990 2692 2993 2708
rect 2974 2658 2982 2661
rect 2954 2648 2958 2651
rect 2982 2648 2990 2651
rect 2950 2572 2953 2628
rect 2926 2562 2929 2568
rect 2930 2538 2934 2541
rect 2926 2502 2929 2518
rect 2934 2512 2937 2538
rect 2958 2532 2961 2598
rect 2982 2592 2985 2648
rect 2998 2641 3001 2838
rect 3006 2782 3009 2818
rect 3030 2772 3033 2818
rect 3006 2762 3009 2768
rect 3006 2662 3009 2758
rect 3014 2742 3017 2748
rect 3006 2652 3009 2658
rect 2998 2638 3009 2641
rect 3006 2592 3009 2638
rect 2966 2542 2969 2548
rect 2974 2532 2977 2538
rect 2958 2522 2961 2528
rect 2926 2482 2929 2488
rect 2934 2482 2937 2498
rect 2934 2412 2937 2468
rect 2942 2452 2945 2518
rect 2958 2462 2961 2508
rect 2982 2482 2985 2578
rect 3022 2572 3025 2718
rect 3038 2692 3041 2938
rect 3070 2932 3073 2938
rect 3048 2903 3050 2907
rect 3054 2903 3057 2907
rect 3061 2903 3064 2907
rect 3078 2902 3081 2918
rect 3070 2882 3073 2898
rect 3078 2878 3086 2881
rect 3050 2858 3054 2861
rect 3046 2752 3049 2858
rect 3078 2792 3081 2878
rect 3094 2862 3097 2938
rect 3094 2852 3097 2858
rect 3062 2752 3065 2758
rect 3078 2752 3081 2768
rect 3048 2703 3050 2707
rect 3054 2703 3057 2707
rect 3061 2703 3064 2707
rect 3030 2672 3033 2678
rect 3078 2662 3081 2748
rect 3094 2702 3097 2818
rect 3102 2762 3105 2918
rect 3118 2862 3121 2918
rect 3126 2892 3129 2938
rect 3158 2932 3161 2938
rect 3150 2911 3153 2918
rect 3150 2908 3161 2911
rect 3150 2882 3153 2898
rect 3142 2762 3145 2858
rect 3158 2772 3161 2908
rect 3174 2862 3177 2938
rect 3190 2932 3193 2938
rect 3182 2851 3185 2918
rect 3190 2912 3193 2928
rect 3190 2862 3193 2868
rect 3182 2848 3190 2851
rect 3130 2748 3134 2751
rect 3102 2722 3105 2728
rect 3098 2688 3102 2691
rect 3094 2662 3097 2678
rect 3026 2568 3033 2571
rect 3006 2552 3009 2568
rect 2994 2538 2998 2541
rect 2998 2482 3001 2498
rect 3022 2492 3025 2558
rect 2970 2468 2974 2471
rect 2982 2462 2985 2468
rect 2970 2458 2974 2461
rect 2918 2362 2921 2368
rect 2926 2352 2929 2358
rect 2950 2352 2953 2398
rect 2958 2352 2961 2358
rect 2974 2352 2977 2358
rect 2986 2348 2990 2351
rect 2918 2332 2921 2338
rect 2950 2322 2953 2338
rect 2982 2322 2985 2338
rect 2998 2331 3001 2378
rect 3006 2342 3009 2468
rect 3030 2452 3033 2568
rect 3038 2492 3041 2648
rect 3078 2552 3081 2558
rect 3110 2551 3113 2718
rect 3150 2712 3153 2728
rect 3158 2712 3161 2728
rect 3174 2712 3177 2818
rect 3198 2762 3201 2898
rect 3206 2832 3209 2918
rect 3214 2902 3217 2958
rect 3230 2952 3233 2958
rect 3222 2872 3225 2908
rect 3222 2762 3225 2868
rect 3230 2852 3233 2948
rect 3294 2942 3297 3058
rect 3314 3048 3318 3051
rect 3290 2938 3294 2941
rect 3238 2932 3241 2938
rect 3246 2912 3249 2938
rect 3302 2931 3305 3018
rect 3334 2972 3337 3118
rect 3350 3041 3353 3088
rect 3382 3063 3385 3068
rect 3350 3038 3361 3041
rect 3342 2952 3345 3018
rect 3358 2962 3361 3038
rect 3390 3032 3393 3278
rect 3398 3252 3401 3318
rect 3406 3282 3409 3318
rect 3422 3282 3425 3338
rect 3410 3258 3414 3261
rect 3430 3261 3433 3338
rect 3438 3282 3441 3298
rect 3426 3258 3433 3261
rect 3446 3232 3449 3468
rect 3454 3352 3457 3658
rect 3568 3603 3570 3607
rect 3574 3603 3577 3607
rect 3581 3603 3584 3607
rect 3590 3602 3593 3718
rect 3614 3672 3617 3818
rect 3630 3752 3633 3918
rect 3710 3912 3713 3958
rect 3722 3948 3726 3951
rect 3738 3938 3742 3941
rect 3750 3892 3753 3988
rect 3758 3892 3761 3968
rect 3774 3942 3777 4048
rect 3830 4032 3833 4048
rect 3798 3952 3801 3978
rect 3806 3962 3809 3998
rect 3782 3942 3785 3948
rect 3774 3932 3777 3938
rect 3798 3902 3801 3948
rect 3806 3942 3809 3958
rect 3814 3952 3817 4018
rect 3830 3952 3833 4028
rect 3838 3982 3841 4048
rect 3854 3961 3857 4018
rect 3850 3958 3857 3961
rect 3854 3942 3857 3948
rect 3862 3942 3865 4018
rect 3878 3962 3881 4058
rect 3894 4052 3897 4058
rect 3906 4038 3910 4041
rect 3918 4032 3921 4058
rect 3934 4052 3937 4058
rect 3942 4042 3945 4138
rect 3990 4102 3993 4148
rect 3982 4062 3985 4088
rect 4006 4072 4009 4138
rect 4022 4131 4025 4248
rect 4038 4182 4041 4258
rect 4070 4252 4073 4318
rect 4080 4303 4082 4307
rect 4086 4303 4089 4307
rect 4093 4303 4096 4307
rect 4102 4302 4105 4318
rect 4134 4312 4137 4318
rect 4122 4288 4126 4291
rect 4094 4272 4097 4288
rect 4102 4262 4105 4278
rect 4126 4262 4129 4268
rect 4134 4262 4137 4298
rect 4090 4258 4094 4261
rect 4114 4258 4118 4261
rect 4078 4192 4081 4228
rect 4038 4152 4041 4158
rect 4062 4152 4065 4158
rect 4022 4128 4038 4131
rect 4054 4122 4057 4148
rect 3994 4068 3998 4071
rect 4030 4062 4033 4118
rect 3970 4058 3974 4061
rect 3938 4038 3942 4041
rect 3950 4032 3953 4058
rect 4030 4052 4033 4058
rect 4018 4048 4022 4051
rect 3958 4042 3961 4048
rect 3966 4022 3969 4048
rect 3922 4018 3926 4021
rect 3926 3952 3929 3958
rect 3874 3948 3878 3951
rect 3890 3948 3894 3951
rect 3902 3942 3905 3948
rect 3814 3938 3822 3941
rect 3678 3872 3681 3878
rect 3702 3872 3705 3878
rect 3670 3782 3673 3868
rect 3738 3866 3742 3869
rect 3698 3858 3702 3861
rect 3678 3852 3681 3858
rect 3718 3772 3721 3858
rect 3758 3852 3761 3878
rect 3774 3862 3777 3898
rect 3798 3892 3801 3898
rect 3814 3892 3817 3938
rect 3838 3932 3841 3938
rect 3878 3932 3881 3938
rect 3918 3932 3921 3948
rect 3898 3928 3902 3931
rect 3822 3922 3825 3928
rect 3830 3922 3833 3928
rect 3910 3912 3913 3918
rect 3926 3892 3929 3938
rect 3878 3882 3881 3888
rect 3934 3882 3937 3938
rect 3942 3882 3945 3968
rect 3950 3942 3953 3948
rect 3958 3942 3961 4008
rect 3966 3952 3969 3978
rect 3982 3962 3985 3968
rect 3990 3952 3993 4018
rect 4030 4002 4033 4048
rect 4006 3952 4009 3988
rect 4022 3962 4025 3968
rect 3974 3932 3977 3938
rect 3954 3928 3958 3931
rect 3786 3878 3790 3881
rect 3846 3872 3849 3878
rect 3918 3872 3921 3878
rect 3930 3868 3934 3871
rect 3738 3748 3742 3751
rect 3662 3672 3665 3718
rect 3710 3712 3713 3738
rect 3734 3722 3737 3738
rect 3758 3712 3761 3848
rect 3766 3792 3769 3828
rect 3774 3732 3777 3858
rect 3782 3732 3785 3868
rect 3826 3858 3830 3861
rect 3806 3832 3809 3858
rect 3814 3761 3817 3848
rect 3810 3758 3817 3761
rect 3806 3752 3809 3758
rect 3830 3752 3833 3858
rect 3838 3832 3841 3868
rect 3974 3862 3977 3898
rect 3982 3872 3985 3948
rect 3990 3942 3993 3948
rect 4038 3932 4041 4108
rect 4046 4081 4049 4118
rect 4046 4078 4054 4081
rect 4050 4068 4054 4071
rect 4062 3992 4065 4148
rect 4080 4103 4082 4107
rect 4086 4103 4089 4107
rect 4093 4103 4096 4107
rect 4102 4102 4105 4258
rect 4110 4152 4113 4158
rect 4118 4142 4121 4188
rect 4078 4062 4081 4068
rect 4070 4002 4073 4058
rect 4086 3962 4089 4068
rect 4094 4052 4097 4058
rect 4110 4052 4113 4078
rect 4118 4022 4121 4138
rect 4126 4122 4129 4258
rect 4142 4192 4145 4268
rect 4150 4262 4153 4298
rect 4166 4272 4169 4318
rect 4158 4252 4161 4258
rect 4170 4248 4174 4251
rect 4190 4242 4193 4338
rect 4230 4332 4233 4378
rect 4278 4362 4281 4368
rect 4242 4348 4246 4351
rect 4282 4348 4286 4351
rect 4198 4272 4201 4318
rect 4238 4302 4241 4338
rect 4246 4302 4249 4318
rect 4238 4282 4241 4288
rect 4262 4282 4265 4348
rect 4274 4338 4278 4341
rect 4270 4272 4273 4318
rect 4294 4272 4297 4348
rect 4302 4342 4305 4348
rect 4318 4332 4321 4398
rect 4326 4352 4329 4358
rect 4342 4352 4345 4358
rect 4350 4351 4353 4398
rect 4382 4392 4385 4428
rect 4430 4402 4433 4428
rect 4362 4358 4366 4361
rect 4414 4352 4417 4368
rect 4442 4358 4446 4361
rect 4350 4348 4358 4351
rect 4386 4348 4390 4351
rect 4446 4348 4454 4351
rect 4474 4348 4478 4351
rect 4490 4348 4494 4351
rect 4330 4338 4334 4341
rect 4354 4338 4358 4341
rect 4306 4288 4310 4291
rect 4370 4288 4374 4291
rect 4358 4281 4361 4288
rect 4358 4278 4369 4281
rect 4254 4262 4257 4268
rect 4134 4162 4137 4168
rect 4146 4158 4150 4161
rect 4158 4151 4161 4158
rect 4154 4148 4161 4151
rect 4174 4152 4177 4178
rect 4182 4142 4185 4168
rect 4198 4162 4201 4258
rect 4206 4252 4209 4258
rect 4230 4182 4233 4258
rect 4238 4162 4241 4248
rect 4262 4212 4265 4258
rect 4270 4252 4273 4268
rect 4290 4258 4294 4261
rect 4278 4202 4281 4258
rect 4298 4248 4302 4251
rect 4302 4232 4305 4238
rect 4198 4152 4201 4158
rect 4206 4142 4209 4158
rect 4218 4148 4222 4151
rect 4186 4138 4193 4141
rect 4134 4112 4137 4138
rect 4174 4131 4177 4138
rect 4174 4128 4185 4131
rect 4126 4082 4129 4088
rect 4126 4062 4129 4078
rect 4134 4062 4137 4068
rect 4142 4062 4145 4068
rect 4150 4062 4153 4098
rect 4166 4072 4169 4078
rect 4174 4072 4177 4118
rect 4182 4112 4185 4128
rect 4190 4082 4193 4138
rect 4206 4092 4209 4108
rect 4214 4081 4217 4098
rect 4206 4078 4217 4081
rect 4198 4072 4201 4078
rect 4170 4058 4182 4061
rect 4150 3992 4153 4008
rect 4058 3948 4062 3951
rect 4038 3922 4041 3928
rect 3998 3882 4001 3918
rect 3890 3858 3894 3861
rect 3914 3858 3918 3861
rect 3938 3858 3942 3861
rect 3986 3858 3990 3861
rect 3838 3762 3841 3828
rect 3846 3752 3849 3858
rect 4006 3852 4009 3898
rect 4046 3882 4049 3938
rect 4102 3912 4105 3948
rect 4126 3942 4129 3948
rect 4080 3903 4082 3907
rect 4086 3903 4089 3907
rect 4093 3903 4096 3907
rect 4058 3888 4062 3891
rect 4038 3872 4041 3878
rect 4018 3868 4022 3871
rect 3866 3848 3870 3851
rect 3890 3848 3894 3851
rect 4030 3842 4033 3858
rect 3862 3792 3865 3838
rect 3978 3828 3982 3831
rect 3926 3792 3929 3808
rect 3854 3762 3857 3768
rect 3926 3752 3929 3758
rect 3934 3752 3937 3768
rect 3966 3752 3969 3788
rect 3974 3752 3977 3778
rect 4006 3752 4009 3788
rect 4046 3752 4049 3878
rect 4058 3868 4062 3871
rect 4062 3862 4065 3868
rect 4078 3862 4081 3878
rect 4102 3872 4105 3888
rect 4078 3852 4081 3858
rect 4066 3848 4070 3851
rect 4122 3848 4126 3851
rect 4134 3832 4137 3948
rect 4142 3872 4145 3958
rect 4158 3872 4161 4018
rect 4166 3952 4169 3978
rect 4206 3952 4209 4078
rect 4214 4062 4217 4068
rect 4222 4062 4225 4108
rect 4230 4072 4233 4138
rect 4238 4102 4241 4158
rect 4234 4068 4238 4071
rect 4246 4061 4249 4198
rect 4254 4162 4257 4168
rect 4286 4162 4289 4168
rect 4266 4158 4270 4161
rect 4294 4152 4297 4198
rect 4302 4152 4305 4208
rect 4254 4142 4257 4148
rect 4262 4132 4265 4138
rect 4262 4072 4265 4128
rect 4270 4062 4273 4138
rect 4294 4132 4297 4138
rect 4302 4112 4305 4148
rect 4310 4142 4313 4158
rect 4318 4142 4321 4258
rect 4326 4232 4329 4268
rect 4334 4252 4337 4258
rect 4350 4252 4353 4258
rect 4358 4242 4361 4268
rect 4366 4252 4369 4278
rect 4382 4252 4385 4348
rect 4398 4342 4401 4348
rect 4418 4338 4422 4341
rect 4390 4332 4393 4338
rect 4406 4332 4409 4338
rect 4430 4332 4433 4348
rect 4390 4272 4393 4318
rect 4406 4272 4409 4288
rect 4422 4282 4425 4298
rect 4438 4282 4441 4318
rect 4446 4302 4449 4348
rect 4458 4338 4462 4341
rect 4478 4312 4481 4318
rect 4486 4312 4489 4328
rect 4502 4282 4505 4378
rect 4566 4362 4569 4368
rect 4514 4348 4518 4351
rect 4538 4348 4542 4351
rect 4582 4342 4585 4348
rect 4462 4262 4465 4278
rect 4502 4272 4505 4278
rect 4470 4262 4473 4268
rect 4390 4202 4393 4258
rect 4398 4212 4401 4258
rect 4334 4152 4337 4178
rect 4406 4172 4409 4228
rect 4430 4182 4433 4258
rect 4478 4252 4481 4258
rect 4458 4248 4462 4251
rect 4486 4232 4489 4268
rect 4494 4262 4497 4268
rect 4510 4242 4513 4328
rect 4518 4292 4521 4338
rect 4526 4282 4529 4318
rect 4534 4312 4537 4328
rect 4550 4272 4553 4318
rect 4522 4268 4526 4271
rect 4362 4158 4366 4161
rect 4394 4158 4398 4161
rect 4362 4148 4366 4151
rect 4382 4142 4385 4158
rect 4406 4142 4409 4168
rect 4438 4162 4441 4208
rect 4446 4162 4449 4168
rect 4438 4152 4441 4158
rect 4454 4152 4457 4218
rect 4518 4212 4521 4248
rect 4502 4152 4505 4188
rect 4514 4158 4518 4161
rect 4534 4152 4537 4258
rect 4542 4212 4545 4258
rect 4550 4192 4553 4268
rect 4558 4181 4561 4268
rect 4566 4262 4569 4268
rect 4550 4178 4561 4181
rect 4466 4148 4470 4151
rect 4482 4148 4486 4151
rect 4522 4148 4526 4151
rect 4430 4142 4433 4148
rect 4418 4138 4422 4141
rect 4326 4132 4329 4138
rect 4366 4132 4369 4138
rect 4318 4092 4321 4098
rect 4290 4068 4294 4071
rect 4322 4068 4326 4071
rect 4242 4058 4249 4061
rect 4258 4058 4262 4061
rect 4298 4058 4302 4061
rect 4322 4058 4326 4061
rect 4222 4032 4225 4058
rect 4246 3972 4249 4058
rect 4258 4048 4262 4051
rect 4334 4051 4337 4128
rect 4438 4112 4441 4138
rect 4362 4068 4366 4071
rect 4326 4048 4337 4051
rect 4270 4042 4273 4048
rect 4286 4042 4289 4048
rect 4318 4042 4321 4048
rect 4246 3952 4249 3958
rect 4318 3952 4321 4038
rect 4326 3992 4329 4048
rect 4334 3962 4337 4018
rect 4350 3982 4353 4038
rect 4358 3952 4361 3968
rect 4374 3952 4377 4108
rect 4446 4092 4449 4148
rect 4454 4142 4457 4148
rect 4478 4122 4481 4138
rect 4486 4122 4489 4128
rect 4510 4102 4513 4138
rect 4534 4092 4537 4148
rect 4542 4102 4545 4138
rect 4390 4072 4393 4088
rect 4398 4062 4401 4078
rect 4422 4072 4425 4088
rect 4430 4062 4433 4078
rect 4470 4062 4473 4088
rect 4514 4078 4518 4081
rect 4478 4072 4481 4078
rect 4506 4068 4510 4071
rect 4506 4058 4510 4061
rect 4390 4002 4393 4058
rect 4422 4052 4425 4058
rect 4454 4052 4457 4058
rect 4526 4052 4529 4078
rect 4542 4072 4545 4078
rect 4550 4072 4553 4178
rect 4562 4148 4566 4151
rect 4574 4142 4577 4228
rect 4582 4152 4585 4248
rect 4590 4222 4593 4338
rect 4598 4152 4601 4158
rect 4558 4122 4561 4128
rect 4590 4112 4593 4138
rect 4558 4072 4561 4108
rect 4570 4068 4574 4071
rect 4410 4048 4414 4051
rect 4490 4048 4494 4051
rect 4446 4042 4449 4048
rect 4470 4042 4473 4048
rect 4194 3948 4198 3951
rect 4234 3948 4238 3951
rect 4274 3948 4278 3951
rect 4366 3942 4369 3948
rect 4178 3938 4182 3941
rect 4218 3938 4222 3941
rect 4250 3938 4254 3941
rect 4306 3938 4310 3941
rect 4190 3932 4193 3938
rect 4162 3858 4166 3861
rect 4174 3842 4177 3908
rect 4054 3752 4057 3788
rect 4134 3772 4137 3828
rect 4142 3762 4145 3818
rect 4106 3758 4110 3761
rect 4174 3752 4177 3838
rect 4190 3832 4193 3918
rect 4214 3872 4217 3908
rect 4222 3902 4225 3918
rect 4230 3872 4233 3938
rect 4238 3932 4241 3938
rect 4294 3932 4297 3938
rect 4350 3932 4353 3938
rect 4298 3918 4302 3921
rect 4210 3868 4214 3871
rect 4222 3862 4225 3868
rect 4198 3812 4201 3858
rect 4206 3792 4209 3858
rect 4230 3852 4233 3868
rect 4238 3862 4241 3918
rect 4270 3882 4273 3918
rect 4334 3881 4337 3928
rect 4334 3878 4345 3881
rect 4266 3868 4270 3871
rect 4274 3858 4286 3861
rect 4290 3858 4294 3861
rect 4262 3851 4265 3858
rect 4262 3848 4278 3851
rect 4214 3792 4217 3848
rect 4246 3832 4249 3848
rect 4194 3788 4198 3791
rect 4230 3752 4233 3808
rect 3882 3748 3889 3751
rect 3798 3732 3801 3748
rect 3826 3738 3830 3741
rect 3806 3732 3809 3738
rect 3838 3732 3841 3748
rect 3874 3728 3878 3731
rect 3782 3722 3785 3728
rect 3814 3712 3817 3718
rect 3774 3682 3777 3698
rect 3782 3692 3785 3708
rect 3630 3663 3633 3668
rect 3726 3662 3729 3668
rect 3694 3612 3697 3618
rect 3462 3562 3465 3598
rect 3510 3562 3513 3588
rect 3610 3578 3614 3581
rect 3542 3551 3545 3558
rect 3494 3542 3497 3548
rect 3574 3542 3577 3548
rect 3462 3512 3465 3518
rect 3470 3512 3473 3528
rect 3494 3472 3497 3538
rect 3510 3532 3513 3538
rect 3654 3532 3657 3547
rect 3686 3542 3689 3548
rect 3518 3482 3521 3498
rect 3550 3482 3553 3498
rect 3514 3478 3518 3481
rect 3622 3472 3625 3478
rect 3466 3468 3470 3471
rect 3514 3468 3518 3471
rect 3574 3462 3577 3468
rect 3654 3463 3657 3468
rect 3482 3458 3486 3461
rect 3602 3458 3606 3461
rect 3462 3452 3465 3458
rect 3462 3392 3465 3448
rect 3598 3442 3601 3448
rect 3606 3442 3609 3448
rect 3522 3438 3526 3441
rect 3534 3412 3537 3438
rect 3568 3403 3570 3407
rect 3574 3403 3577 3407
rect 3581 3403 3584 3407
rect 3614 3382 3617 3418
rect 3474 3378 3489 3381
rect 3486 3372 3489 3378
rect 3502 3372 3505 3378
rect 3478 3362 3481 3368
rect 3638 3362 3641 3378
rect 3462 3352 3465 3358
rect 3526 3352 3529 3358
rect 3550 3352 3553 3358
rect 3454 3332 3457 3348
rect 3622 3342 3625 3348
rect 3646 3342 3649 3348
rect 3482 3338 3486 3341
rect 3506 3338 3510 3341
rect 3530 3338 3534 3341
rect 3554 3338 3558 3341
rect 3578 3338 3582 3341
rect 3454 3221 3457 3228
rect 3450 3218 3457 3221
rect 3430 3142 3433 3147
rect 3494 3142 3497 3318
rect 3502 3252 3505 3258
rect 3510 3151 3513 3328
rect 3518 3312 3521 3318
rect 3526 3272 3529 3278
rect 3542 3252 3545 3318
rect 3558 3242 3561 3318
rect 3598 3302 3601 3328
rect 3598 3282 3601 3298
rect 3566 3222 3569 3258
rect 3606 3242 3609 3248
rect 3518 3192 3521 3218
rect 3506 3148 3513 3151
rect 3558 3152 3561 3218
rect 3568 3203 3570 3207
rect 3574 3203 3577 3207
rect 3581 3203 3584 3207
rect 3574 3151 3577 3158
rect 3398 3112 3401 3128
rect 3414 3062 3417 3138
rect 3498 3118 3502 3121
rect 3454 3082 3457 3098
rect 3458 3068 3462 3071
rect 3414 2952 3417 3058
rect 3470 3052 3473 3108
rect 3510 3082 3513 3148
rect 3518 3072 3521 3118
rect 3566 3082 3569 3098
rect 3582 3072 3585 3138
rect 3606 3102 3609 3238
rect 3638 3132 3641 3318
rect 3646 3172 3649 3298
rect 3662 3282 3665 3468
rect 3686 3462 3689 3538
rect 3674 3358 3678 3361
rect 3690 3348 3694 3351
rect 3670 3332 3673 3348
rect 3690 3338 3694 3341
rect 3702 3332 3705 3658
rect 3734 3652 3737 3678
rect 3814 3662 3817 3668
rect 3746 3658 3750 3661
rect 3722 3588 3726 3591
rect 3738 3568 3742 3571
rect 3726 3562 3729 3568
rect 3742 3552 3745 3558
rect 3750 3552 3753 3618
rect 3798 3551 3801 3568
rect 3722 3488 3726 3491
rect 3742 3482 3745 3548
rect 3766 3512 3769 3528
rect 3750 3482 3753 3498
rect 3806 3492 3809 3538
rect 3742 3472 3745 3478
rect 3742 3462 3745 3468
rect 3770 3458 3774 3461
rect 3786 3458 3790 3461
rect 3726 3452 3729 3458
rect 3746 3448 3750 3451
rect 3786 3448 3790 3451
rect 3734 3382 3737 3388
rect 3742 3362 3745 3368
rect 3806 3352 3809 3418
rect 3726 3342 3729 3348
rect 3774 3342 3777 3347
rect 3718 3312 3721 3328
rect 3702 3282 3705 3288
rect 3742 3282 3745 3298
rect 3662 3272 3665 3278
rect 3670 3263 3673 3278
rect 3702 3252 3705 3258
rect 3662 3152 3665 3218
rect 3670 3162 3673 3238
rect 3718 3222 3721 3258
rect 3750 3252 3753 3318
rect 3806 3272 3809 3348
rect 3822 3301 3825 3728
rect 3886 3722 3889 3748
rect 4018 3748 4022 3751
rect 4082 3748 4086 3751
rect 3894 3732 3897 3738
rect 3910 3732 3913 3748
rect 3910 3662 3913 3728
rect 3926 3672 3929 3748
rect 3946 3738 3950 3741
rect 4018 3738 4022 3741
rect 4082 3738 4086 3741
rect 3958 3732 3961 3738
rect 3958 3692 3961 3718
rect 3830 3352 3833 3658
rect 3902 3592 3905 3659
rect 3874 3568 3878 3571
rect 3886 3542 3889 3558
rect 3950 3552 3953 3638
rect 3982 3562 3985 3738
rect 3998 3732 4001 3738
rect 4038 3732 4041 3738
rect 3998 3682 4001 3718
rect 4026 3668 4030 3671
rect 3990 3632 3993 3668
rect 4038 3662 4041 3718
rect 4070 3671 4073 3718
rect 4126 3712 4129 3748
rect 4080 3703 4082 3707
rect 4086 3703 4089 3707
rect 4093 3703 4096 3707
rect 4070 3668 4081 3671
rect 4026 3658 4030 3661
rect 4070 3652 4073 3658
rect 4078 3652 4081 3668
rect 4110 3662 4113 3708
rect 4134 3682 4137 3738
rect 4158 3712 4161 3748
rect 4202 3738 4206 3741
rect 4166 3682 4169 3738
rect 4118 3672 4121 3678
rect 4142 3672 4145 3681
rect 4146 3668 4150 3671
rect 4178 3668 4182 3671
rect 4218 3668 4222 3671
rect 4114 3658 4118 3661
rect 4094 3652 4097 3658
rect 4126 3652 4129 3668
rect 4146 3658 4150 3661
rect 4178 3658 4182 3661
rect 4210 3658 4214 3661
rect 4018 3648 4022 3651
rect 4050 3648 4054 3651
rect 4154 3648 4158 3651
rect 4186 3648 4190 3651
rect 4030 3642 4033 3648
rect 3922 3547 3926 3550
rect 4014 3551 4017 3578
rect 3950 3542 3953 3548
rect 3998 3542 4001 3548
rect 3862 3522 3865 3528
rect 3862 3472 3865 3478
rect 3842 3368 3846 3371
rect 3862 3352 3865 3458
rect 3870 3452 3873 3518
rect 3886 3462 3889 3538
rect 3910 3482 3913 3498
rect 3950 3472 3953 3538
rect 3986 3518 3993 3521
rect 3946 3459 3950 3462
rect 3886 3442 3889 3448
rect 3990 3432 3993 3518
rect 4006 3472 4009 3488
rect 3886 3362 3889 3378
rect 4022 3352 4025 3618
rect 4038 3482 4041 3538
rect 4038 3452 4041 3459
rect 3886 3342 3889 3348
rect 3918 3342 3921 3347
rect 4070 3342 4073 3648
rect 4110 3542 4113 3548
rect 4098 3518 4105 3521
rect 4080 3503 4082 3507
rect 4086 3503 4089 3507
rect 4093 3503 4096 3507
rect 4102 3452 4105 3518
rect 4126 3492 4129 3547
rect 4214 3542 4217 3628
rect 4230 3622 4233 3748
rect 4242 3738 4246 3741
rect 4254 3692 4257 3768
rect 4294 3762 4297 3768
rect 4262 3752 4265 3758
rect 4274 3748 4278 3751
rect 4302 3742 4305 3868
rect 4310 3852 4313 3878
rect 4310 3752 4313 3758
rect 4266 3738 4270 3741
rect 4254 3662 4257 3688
rect 4262 3672 4265 3678
rect 4286 3672 4289 3728
rect 4310 3662 4313 3718
rect 4318 3672 4321 3878
rect 4330 3868 4334 3871
rect 4334 3762 4337 3858
rect 4342 3812 4345 3878
rect 4350 3862 4353 3898
rect 4374 3882 4377 3948
rect 4390 3942 4393 3998
rect 4430 3962 4433 3988
rect 4446 3952 4449 3958
rect 4462 3952 4465 3968
rect 4474 3958 4478 3961
rect 4410 3948 4414 3951
rect 4438 3942 4441 3948
rect 4470 3942 4473 3948
rect 4382 3932 4385 3938
rect 4390 3892 4393 3928
rect 4398 3922 4401 3928
rect 4378 3858 4382 3861
rect 4366 3852 4369 3858
rect 4326 3752 4329 3758
rect 4334 3752 4337 3758
rect 4358 3742 4361 3758
rect 4366 3752 4369 3758
rect 4374 3742 4377 3848
rect 4406 3842 4409 3858
rect 4398 3752 4401 3758
rect 4406 3752 4409 3838
rect 4330 3738 4334 3741
rect 4386 3738 4390 3741
rect 4398 3732 4401 3738
rect 4398 3692 4401 3718
rect 4382 3662 4385 3688
rect 4414 3662 4417 3938
rect 4486 3932 4489 3948
rect 4450 3918 4454 3921
rect 4434 3888 4438 3891
rect 4446 3882 4449 3888
rect 4474 3868 4478 3871
rect 4430 3862 4433 3868
rect 4450 3858 4454 3861
rect 4454 3852 4457 3858
rect 4462 3842 4465 3868
rect 4486 3862 4489 3888
rect 4494 3862 4497 3978
rect 4502 3932 4505 3938
rect 4510 3892 4513 4048
rect 4534 4042 4537 4058
rect 4542 4032 4545 4038
rect 4518 3982 4521 3988
rect 4542 3972 4545 3978
rect 4526 3952 4529 3968
rect 4534 3942 4537 3958
rect 4546 3948 4550 3951
rect 4518 3912 4521 3938
rect 4558 3932 4561 4068
rect 4578 4058 4582 4061
rect 4566 4052 4569 4058
rect 4598 4042 4601 4048
rect 4582 3962 4585 3968
rect 4566 3952 4569 3958
rect 4582 3942 4585 3948
rect 4534 3872 4537 3878
rect 4554 3868 4558 3871
rect 4438 3792 4441 3828
rect 4462 3802 4465 3818
rect 4422 3742 4425 3748
rect 4430 3692 4433 3738
rect 4438 3731 4441 3768
rect 4478 3762 4481 3798
rect 4486 3752 4489 3808
rect 4450 3738 4454 3741
rect 4454 3732 4457 3738
rect 4438 3728 4446 3731
rect 4462 3722 4465 3748
rect 4502 3742 4505 3868
rect 4526 3852 4529 3858
rect 4514 3768 4529 3771
rect 4526 3762 4529 3768
rect 4518 3752 4521 3758
rect 4534 3752 4537 3868
rect 4590 3862 4593 3958
rect 4598 3932 4601 4028
rect 4542 3802 4545 3818
rect 4582 3762 4585 3798
rect 4510 3742 4513 3748
rect 4478 3662 4481 3698
rect 4486 3672 4489 3738
rect 4510 3672 4513 3738
rect 4506 3668 4510 3671
rect 4518 3662 4521 3748
rect 4550 3732 4553 3738
rect 4534 3662 4537 3718
rect 4542 3672 4545 3728
rect 4566 3722 4569 3748
rect 4570 3668 4574 3671
rect 4282 3658 4286 3661
rect 4410 3658 4414 3661
rect 4310 3652 4313 3658
rect 4326 3642 4329 3658
rect 4374 3642 4377 3658
rect 4446 3622 4449 3658
rect 4542 3652 4545 3658
rect 4518 3642 4521 3648
rect 4502 3632 4505 3638
rect 4238 3552 4241 3558
rect 4270 3551 4273 3598
rect 4326 3582 4329 3618
rect 4218 3538 4222 3541
rect 4182 3492 4185 3508
rect 4110 3472 4113 3478
rect 4206 3472 4209 3538
rect 4254 3512 4257 3538
rect 4102 3392 4105 3418
rect 3814 3298 3825 3301
rect 3766 3222 3769 3268
rect 3798 3252 3801 3259
rect 3686 3162 3689 3168
rect 3758 3162 3761 3218
rect 3770 3188 3774 3191
rect 3682 3148 3686 3151
rect 3738 3148 3742 3151
rect 3754 3148 3758 3151
rect 3662 3142 3665 3148
rect 3638 3112 3641 3118
rect 3654 3101 3657 3118
rect 3710 3112 3713 3128
rect 3718 3112 3721 3128
rect 3654 3098 3665 3101
rect 3490 3068 3494 3071
rect 3518 3062 3521 3068
rect 3542 3062 3545 3068
rect 3498 3058 3502 3061
rect 3530 3058 3534 3061
rect 3630 3062 3633 3068
rect 3614 3052 3617 3059
rect 3506 3048 3510 3051
rect 3450 3038 3454 3041
rect 3458 2988 3462 2991
rect 3342 2942 3345 2948
rect 3358 2942 3361 2948
rect 3418 2948 3422 2951
rect 3390 2942 3393 2947
rect 3314 2938 3318 2941
rect 3302 2928 3313 2931
rect 3274 2918 3278 2921
rect 3238 2892 3241 2898
rect 3254 2872 3257 2888
rect 3262 2872 3265 2918
rect 3278 2892 3281 2898
rect 3246 2822 3249 2868
rect 3246 2812 3249 2818
rect 3254 2772 3257 2868
rect 3294 2852 3297 2858
rect 3302 2852 3305 2918
rect 3310 2912 3313 2928
rect 3318 2912 3321 2928
rect 3326 2892 3329 2928
rect 3342 2902 3345 2938
rect 3338 2888 3342 2891
rect 3318 2872 3321 2878
rect 3334 2862 3337 2878
rect 3266 2848 3270 2851
rect 3246 2762 3249 2768
rect 3222 2752 3225 2758
rect 3186 2748 3190 2751
rect 3242 2748 3246 2751
rect 3278 2742 3281 2747
rect 3198 2702 3201 2718
rect 3206 2712 3209 2728
rect 3278 2682 3281 2728
rect 3182 2672 3185 2678
rect 3154 2658 3158 2661
rect 3150 2592 3153 2628
rect 3150 2552 3153 2568
rect 3146 2538 3153 2541
rect 3048 2503 3050 2507
rect 3054 2503 3057 2507
rect 3061 2503 3064 2507
rect 3078 2502 3081 2528
rect 3106 2478 3110 2481
rect 3126 2472 3129 2538
rect 3058 2468 3062 2471
rect 3058 2358 3062 2361
rect 3014 2342 3017 2358
rect 3038 2342 3041 2348
rect 2998 2328 3006 2331
rect 2990 2282 2993 2298
rect 3030 2282 3033 2338
rect 3046 2331 3049 2338
rect 3038 2328 3049 2331
rect 3038 2292 3041 2328
rect 3048 2303 3050 2307
rect 3054 2303 3057 2307
rect 3061 2303 3064 2307
rect 2998 2272 3001 2278
rect 3062 2272 3065 2278
rect 3070 2272 3073 2338
rect 3010 2268 3014 2271
rect 2918 2262 2921 2268
rect 2930 2258 2934 2261
rect 2954 2258 2958 2261
rect 2978 2258 2982 2261
rect 3022 2252 3025 2258
rect 3046 2252 3049 2258
rect 2942 2242 2945 2248
rect 2962 2238 2966 2241
rect 2906 2188 2910 2191
rect 2918 2182 2921 2188
rect 3006 2162 3009 2178
rect 2758 2122 2761 2148
rect 2782 2142 2785 2158
rect 2798 2142 2801 2148
rect 2766 2122 2769 2138
rect 2806 2132 2809 2158
rect 2842 2148 2846 2151
rect 2822 2132 2825 2138
rect 2778 2128 2782 2131
rect 2758 2102 2761 2118
rect 2782 2092 2785 2118
rect 2758 2072 2761 2078
rect 2626 2068 2630 2071
rect 2722 2068 2726 2071
rect 2574 2052 2577 2068
rect 2598 2022 2601 2068
rect 2606 2012 2609 2068
rect 2686 2062 2689 2068
rect 2710 2062 2713 2068
rect 2650 2058 2654 2061
rect 2630 2052 2633 2058
rect 2678 2052 2681 2058
rect 2646 2012 2649 2048
rect 2710 2032 2713 2048
rect 2750 2032 2753 2068
rect 2762 2058 2766 2061
rect 2774 2052 2777 2068
rect 2790 2061 2793 2078
rect 2798 2072 2801 2128
rect 2814 2062 2817 2118
rect 2838 2082 2841 2128
rect 2862 2092 2865 2118
rect 2870 2082 2873 2138
rect 2910 2132 2913 2138
rect 2926 2132 2929 2158
rect 3006 2152 3009 2158
rect 3038 2152 3041 2198
rect 3026 2148 3030 2151
rect 3038 2142 3041 2148
rect 3062 2142 3065 2178
rect 3078 2172 3081 2468
rect 3122 2458 3126 2461
rect 3150 2421 3153 2538
rect 3166 2492 3169 2558
rect 3182 2542 3185 2668
rect 3198 2662 3201 2668
rect 3202 2648 3206 2651
rect 3214 2572 3217 2658
rect 3198 2551 3201 2558
rect 3198 2492 3201 2518
rect 3182 2472 3185 2478
rect 3170 2448 3174 2451
rect 3182 2432 3185 2468
rect 3142 2418 3153 2421
rect 3142 2392 3145 2418
rect 3190 2392 3193 2468
rect 3206 2452 3209 2568
rect 3222 2492 3225 2618
rect 3222 2482 3225 2488
rect 3230 2462 3233 2678
rect 3278 2672 3281 2678
rect 3270 2652 3273 2659
rect 3278 2592 3281 2628
rect 3266 2538 3270 2541
rect 3262 2512 3265 2518
rect 3238 2482 3241 2488
rect 3254 2482 3257 2498
rect 3286 2472 3289 2558
rect 3294 2542 3297 2768
rect 3310 2732 3313 2748
rect 3334 2671 3337 2798
rect 3350 2762 3353 2868
rect 3394 2858 3398 2861
rect 3390 2822 3393 2858
rect 3358 2721 3361 2808
rect 3398 2762 3401 2828
rect 3366 2752 3369 2758
rect 3414 2752 3417 2758
rect 3402 2738 3406 2741
rect 3422 2732 3425 2868
rect 3454 2862 3457 2898
rect 3470 2871 3473 3008
rect 3486 2951 3489 3018
rect 3568 3003 3570 3007
rect 3574 3003 3577 3007
rect 3581 3003 3584 3007
rect 3630 2992 3633 3058
rect 3630 2952 3633 2988
rect 3662 2982 3665 3098
rect 3686 3062 3689 3078
rect 3706 3068 3710 3071
rect 3726 3062 3729 3068
rect 3750 3062 3753 3128
rect 3814 3092 3817 3298
rect 3822 3152 3825 3158
rect 3682 3018 3686 3021
rect 3646 2962 3649 2968
rect 3702 2952 3705 3018
rect 3710 2962 3713 3008
rect 3514 2948 3518 2951
rect 3666 2948 3670 2951
rect 3722 2948 3726 2951
rect 3570 2938 3574 2941
rect 3714 2938 3718 2941
rect 3478 2882 3481 2898
rect 3502 2872 3505 2898
rect 3470 2868 3481 2871
rect 3438 2852 3441 2858
rect 3478 2852 3481 2868
rect 3510 2852 3513 2918
rect 3518 2862 3521 2868
rect 3526 2862 3529 2898
rect 3502 2842 3505 2848
rect 3454 2752 3457 2818
rect 3470 2751 3473 2758
rect 3502 2732 3505 2748
rect 3358 2718 3369 2721
rect 3342 2692 3345 2718
rect 3334 2668 3342 2671
rect 3318 2592 3321 2638
rect 3334 2572 3337 2618
rect 3350 2602 3353 2718
rect 3358 2692 3361 2708
rect 3366 2672 3369 2718
rect 3390 2712 3393 2728
rect 3430 2692 3433 2718
rect 3438 2712 3441 2728
rect 3518 2692 3521 2728
rect 3534 2672 3537 2938
rect 3554 2918 3558 2921
rect 3550 2882 3553 2898
rect 3646 2872 3649 2918
rect 3686 2912 3689 2928
rect 3694 2912 3697 2928
rect 3568 2803 3570 2807
rect 3574 2803 3577 2807
rect 3581 2803 3584 2807
rect 3582 2742 3585 2747
rect 3598 2742 3601 2868
rect 3606 2862 3609 2868
rect 3670 2852 3673 2858
rect 3666 2828 3670 2831
rect 3646 2762 3649 2768
rect 3678 2751 3681 2908
rect 3702 2871 3705 2918
rect 3710 2882 3713 2898
rect 3702 2868 3710 2871
rect 3726 2862 3729 2948
rect 3698 2858 3702 2861
rect 3686 2752 3689 2818
rect 3726 2772 3729 2838
rect 3662 2742 3665 2748
rect 3566 2732 3569 2738
rect 3374 2668 3382 2671
rect 3410 2668 3414 2671
rect 3442 2668 3446 2671
rect 3466 2668 3470 2671
rect 3362 2648 3366 2651
rect 3374 2642 3377 2668
rect 3386 2658 3390 2661
rect 3462 2652 3465 2658
rect 3402 2648 3406 2651
rect 3426 2648 3430 2651
rect 3450 2648 3454 2651
rect 3306 2558 3310 2561
rect 3330 2558 3334 2561
rect 3314 2548 3318 2551
rect 3334 2542 3337 2548
rect 3350 2542 3353 2588
rect 3366 2551 3369 2598
rect 3318 2532 3321 2538
rect 3382 2492 3385 2648
rect 3394 2638 3398 2641
rect 3454 2562 3457 2648
rect 3534 2612 3537 2668
rect 3462 2562 3465 2568
rect 3470 2551 3473 2558
rect 3466 2548 3473 2551
rect 3486 2552 3489 2568
rect 3494 2562 3497 2578
rect 3538 2558 3542 2561
rect 3550 2552 3553 2718
rect 3598 2672 3601 2738
rect 3662 2682 3665 2688
rect 3710 2682 3713 2698
rect 3694 2672 3697 2678
rect 3690 2668 3694 2671
rect 3622 2642 3625 2648
rect 3646 2612 3649 2668
rect 3726 2661 3729 2688
rect 3734 2672 3737 2858
rect 3742 2852 3745 2978
rect 3782 2942 3785 2947
rect 3790 2942 3793 3038
rect 3750 2912 3753 2928
rect 3806 2902 3809 3018
rect 3758 2842 3761 2868
rect 3774 2863 3777 2868
rect 3746 2778 3750 2781
rect 3742 2758 3750 2761
rect 3742 2712 3745 2758
rect 3742 2672 3745 2678
rect 3726 2658 3734 2661
rect 3742 2652 3745 2668
rect 3766 2662 3769 2678
rect 3774 2672 3777 2738
rect 3786 2728 3790 2731
rect 3798 2722 3801 2758
rect 3786 2688 3790 2691
rect 3798 2682 3801 2688
rect 3806 2682 3809 2798
rect 3818 2738 3822 2741
rect 3830 2702 3833 3338
rect 3846 3312 3849 3328
rect 3862 3282 3865 3288
rect 3902 3272 3905 3338
rect 3934 3332 3937 3338
rect 4030 3332 4033 3338
rect 3982 3302 3985 3318
rect 4014 3282 4017 3288
rect 4030 3272 4033 3328
rect 3986 3268 3990 3271
rect 3894 3263 3897 3268
rect 3894 3258 3897 3259
rect 4018 3258 4022 3261
rect 3890 3147 3894 3150
rect 3918 3142 3921 3148
rect 3942 3072 3945 3238
rect 4006 3182 4009 3248
rect 4070 3202 4073 3338
rect 4080 3303 4082 3307
rect 4086 3303 4089 3307
rect 4093 3303 4096 3307
rect 4110 3272 4113 3468
rect 4222 3463 4225 3468
rect 4222 3458 4225 3459
rect 4190 3392 4193 3438
rect 4126 3351 4129 3368
rect 4222 3351 4225 3428
rect 4230 3342 4233 3508
rect 4126 3322 4129 3328
rect 4126 3272 4129 3318
rect 4206 3292 4209 3338
rect 4214 3272 4217 3278
rect 4070 3172 4073 3178
rect 3950 3162 3953 3168
rect 3966 3142 3969 3148
rect 4074 3148 4078 3151
rect 3982 3122 3985 3147
rect 3998 3072 4001 3078
rect 4014 3072 4017 3148
rect 4046 3142 4049 3148
rect 4102 3142 4105 3268
rect 4142 3192 4145 3259
rect 4218 3258 4222 3261
rect 4190 3192 4193 3238
rect 4198 3151 4201 3158
rect 4078 3122 4081 3138
rect 4080 3103 4082 3107
rect 4086 3103 4089 3107
rect 4093 3103 4096 3107
rect 3850 2968 3854 2971
rect 3854 2952 3857 2958
rect 3846 2862 3849 2868
rect 3854 2851 3857 2918
rect 3862 2892 3865 3058
rect 3878 2992 3881 3058
rect 3934 2992 3937 3059
rect 3998 2951 4001 2968
rect 3870 2862 3873 2938
rect 3886 2882 3889 2898
rect 3894 2882 3897 2898
rect 3918 2882 3921 2948
rect 4014 2942 4017 3068
rect 4030 3042 4033 3059
rect 4062 3052 4065 3058
rect 4094 2992 4097 3058
rect 4102 2942 4105 3138
rect 4110 3082 4113 3088
rect 4118 3072 4121 3128
rect 4150 3072 4153 3088
rect 4122 3058 4126 3061
rect 4150 3052 4153 3068
rect 4158 3052 4161 3118
rect 4174 3072 4177 3108
rect 4206 3082 4209 3188
rect 4170 3058 4174 3061
rect 4030 2892 4033 2928
rect 4080 2903 4082 2907
rect 4086 2903 4089 2907
rect 4093 2903 4096 2907
rect 4142 2882 4145 2888
rect 4158 2872 4161 3048
rect 4206 3022 4209 3059
rect 4166 2942 4169 2948
rect 4182 2942 4185 2948
rect 4198 2922 4201 2947
rect 3866 2858 3870 2861
rect 3914 2858 3918 2861
rect 3850 2848 3857 2851
rect 3930 2848 3934 2851
rect 3950 2842 3953 2868
rect 3966 2863 3969 2868
rect 4110 2862 4113 2868
rect 4158 2862 4161 2868
rect 3838 2802 3841 2818
rect 3854 2742 3857 2838
rect 3918 2752 3921 2818
rect 3982 2762 3985 2808
rect 3874 2747 3878 2750
rect 3838 2722 3841 2728
rect 3790 2672 3793 2678
rect 3854 2672 3857 2738
rect 3942 2732 3945 2758
rect 3982 2742 3985 2758
rect 3998 2742 4001 2758
rect 4014 2742 4017 2838
rect 4030 2772 4033 2818
rect 4078 2812 4081 2859
rect 4174 2792 4177 2859
rect 4098 2788 4102 2791
rect 4078 2752 4081 2768
rect 4034 2747 4038 2750
rect 4142 2742 4145 2748
rect 4122 2738 4126 2741
rect 3930 2718 3934 2721
rect 3966 2702 3969 2718
rect 3906 2668 3910 2671
rect 3750 2652 3753 2658
rect 3774 2652 3777 2668
rect 3838 2652 3841 2659
rect 3714 2648 3718 2651
rect 3670 2632 3673 2648
rect 3568 2603 3570 2607
rect 3574 2603 3577 2607
rect 3581 2603 3584 2607
rect 3578 2568 3582 2571
rect 3566 2552 3569 2558
rect 3414 2501 3417 2548
rect 3434 2538 3438 2541
rect 3562 2538 3566 2541
rect 3486 2532 3489 2538
rect 3430 2522 3433 2528
rect 3406 2498 3417 2501
rect 3294 2472 3297 2488
rect 3406 2482 3409 2498
rect 3342 2472 3345 2478
rect 3314 2468 3318 2471
rect 3218 2438 3222 2441
rect 3230 2412 3233 2418
rect 3246 2402 3249 2418
rect 3134 2352 3137 2358
rect 3090 2348 3094 2351
rect 3158 2342 3161 2348
rect 3106 2338 3110 2341
rect 3094 2332 3097 2338
rect 3118 2332 3121 2338
rect 3174 2332 3177 2378
rect 3214 2362 3217 2388
rect 3262 2372 3265 2458
rect 3286 2452 3289 2468
rect 3430 2462 3433 2488
rect 3478 2482 3481 2488
rect 3486 2482 3489 2488
rect 3438 2472 3441 2478
rect 3462 2462 3465 2478
rect 3474 2468 3478 2471
rect 3510 2462 3513 2478
rect 3518 2472 3521 2538
rect 3598 2532 3601 2578
rect 3538 2528 3542 2531
rect 3598 2492 3601 2498
rect 3558 2482 3561 2488
rect 3570 2478 3574 2481
rect 3522 2468 3526 2471
rect 3546 2468 3550 2471
rect 3586 2468 3590 2471
rect 3606 2462 3609 2548
rect 3622 2482 3625 2578
rect 3630 2552 3633 2608
rect 3638 2562 3641 2568
rect 3650 2558 3654 2561
rect 3630 2542 3633 2548
rect 3674 2538 3678 2541
rect 3694 2532 3697 2598
rect 3834 2568 3838 2571
rect 3742 2558 3750 2561
rect 3762 2558 3766 2561
rect 3734 2542 3737 2558
rect 3742 2552 3745 2558
rect 3798 2552 3801 2558
rect 3822 2542 3825 2558
rect 3858 2548 3878 2551
rect 3886 2542 3889 2618
rect 3894 2542 3897 2668
rect 3902 2602 3905 2618
rect 3910 2572 3913 2658
rect 3918 2622 3921 2628
rect 3926 2611 3929 2658
rect 3934 2652 3937 2698
rect 3982 2692 3985 2738
rect 3942 2672 3945 2678
rect 3982 2672 3985 2688
rect 3962 2658 3966 2661
rect 3990 2661 3993 2718
rect 3998 2682 4001 2738
rect 4158 2732 4161 2747
rect 4206 2742 4209 3018
rect 4222 2792 4225 3208
rect 4230 3152 4233 3338
rect 4246 3272 4249 3498
rect 4294 3472 4297 3498
rect 4318 3492 4321 3548
rect 4342 3542 4345 3558
rect 4350 3542 4353 3548
rect 4334 3522 4337 3528
rect 4358 3472 4361 3618
rect 4366 3552 4369 3618
rect 4462 3592 4465 3618
rect 4422 3551 4425 3568
rect 4534 3562 4537 3578
rect 4514 3558 4518 3561
rect 4566 3552 4569 3578
rect 4574 3552 4577 3618
rect 4514 3538 4518 3541
rect 4382 3482 4385 3518
rect 4406 3512 4409 3538
rect 4494 3532 4497 3538
rect 4366 3472 4369 3478
rect 4282 3468 4286 3471
rect 4326 3462 4329 3468
rect 4350 3462 4353 3468
rect 4298 3458 4302 3461
rect 4254 3262 4257 3458
rect 4314 3448 4318 3451
rect 4318 3382 4321 3448
rect 4310 3352 4313 3358
rect 4326 3352 4329 3458
rect 4354 3448 4358 3451
rect 4370 3448 4374 3451
rect 4382 3442 4385 3468
rect 4390 3442 4393 3458
rect 4334 3362 4337 3368
rect 4242 3248 4246 3251
rect 4254 3242 4257 3248
rect 4262 3181 4265 3268
rect 4270 3252 4273 3328
rect 4278 3272 4281 3348
rect 4294 3342 4297 3348
rect 4306 3338 4310 3341
rect 4318 3312 4321 3338
rect 4342 3262 4345 3288
rect 4262 3178 4273 3181
rect 4262 3162 4265 3168
rect 4270 3142 4273 3178
rect 4278 3152 4281 3258
rect 4302 3241 4305 3248
rect 4302 3238 4313 3241
rect 4290 3158 4294 3161
rect 4270 3112 4273 3138
rect 4278 3102 4281 3148
rect 4294 3142 4297 3148
rect 4274 3078 4278 3081
rect 4294 3072 4297 3108
rect 4278 3062 4281 3068
rect 4302 3062 4305 3098
rect 4282 3048 4286 3051
rect 4278 2992 4281 3028
rect 4310 2992 4313 3238
rect 4326 3152 4329 3218
rect 4350 3142 4353 3348
rect 4358 3342 4361 3348
rect 4366 3282 4369 3308
rect 4366 3262 4369 3268
rect 4358 3258 4366 3261
rect 4358 3152 4361 3258
rect 4390 3232 4393 3347
rect 4406 3342 4409 3508
rect 4486 3472 4489 3518
rect 4430 3462 4433 3468
rect 4454 3462 4457 3468
rect 4502 3462 4505 3468
rect 4430 3452 4433 3458
rect 4510 3452 4513 3518
rect 4518 3462 4521 3468
rect 4542 3452 4545 3458
rect 4350 3072 4353 3128
rect 4390 3102 4393 3118
rect 4390 3072 4393 3078
rect 4350 3052 4353 3058
rect 4318 3042 4321 3048
rect 4318 2981 4321 3038
rect 4310 2978 4321 2981
rect 4290 2948 4294 2951
rect 4270 2942 4273 2948
rect 4290 2938 4294 2941
rect 4254 2922 4257 2938
rect 4238 2892 4241 2908
rect 4254 2872 4257 2918
rect 4310 2912 4313 2978
rect 4326 2961 4329 3038
rect 4358 2992 4361 3058
rect 4378 3048 4382 3051
rect 4398 3051 4401 3338
rect 4414 3272 4417 3338
rect 4414 3262 4417 3268
rect 4430 3242 4433 3259
rect 4406 3182 4409 3188
rect 4414 3152 4417 3158
rect 4422 3142 4425 3158
rect 4430 3152 4433 3178
rect 4438 3172 4441 3448
rect 4502 3442 4505 3448
rect 4550 3442 4553 3448
rect 4526 3432 4529 3438
rect 4454 3352 4457 3358
rect 4478 3332 4481 3348
rect 4486 3342 4489 3378
rect 4506 3358 4510 3361
rect 4546 3358 4550 3361
rect 4522 3348 4526 3351
rect 4534 3332 4537 3338
rect 4542 3331 4545 3358
rect 4558 3352 4561 3468
rect 4566 3462 4569 3538
rect 4590 3522 4593 3558
rect 4566 3392 4569 3458
rect 4590 3362 4593 3518
rect 4542 3328 4553 3331
rect 4494 3312 4497 3318
rect 4438 3152 4441 3168
rect 4478 3162 4481 3308
rect 4494 3292 4497 3298
rect 4510 3292 4513 3308
rect 4530 3278 4534 3281
rect 4526 3262 4529 3268
rect 4542 3252 4545 3318
rect 4550 3262 4553 3328
rect 4558 3302 4561 3338
rect 4566 3292 4569 3318
rect 4534 3152 4537 3168
rect 4550 3162 4553 3258
rect 4570 3248 4574 3251
rect 4562 3158 4566 3161
rect 4506 3148 4510 3151
rect 4462 3142 4465 3148
rect 4486 3142 4489 3148
rect 4562 3138 4566 3141
rect 4406 3092 4409 3138
rect 4446 3092 4449 3108
rect 4438 3072 4441 3088
rect 4454 3081 4457 3138
rect 4446 3078 4457 3081
rect 4486 3082 4489 3098
rect 4398 3048 4406 3051
rect 4406 2962 4409 3048
rect 4446 3032 4449 3078
rect 4510 3072 4513 3138
rect 4538 3068 4542 3071
rect 4454 3052 4457 3068
rect 4462 3042 4465 3068
rect 4478 3052 4481 3068
rect 4510 3062 4513 3068
rect 4538 3058 4542 3061
rect 4470 3042 4473 3048
rect 4326 2958 4337 2961
rect 4318 2952 4321 2958
rect 4334 2952 4337 2958
rect 4350 2952 4353 2958
rect 4326 2942 4329 2948
rect 4318 2872 4321 2938
rect 4326 2862 4329 2938
rect 4334 2892 4337 2938
rect 4366 2921 4369 2928
rect 4382 2922 4385 2938
rect 4398 2932 4401 2947
rect 4366 2918 4377 2921
rect 4358 2892 4361 2898
rect 4342 2872 4345 2878
rect 4270 2832 4273 2859
rect 4358 2852 4361 2868
rect 4374 2852 4377 2918
rect 4382 2862 4385 2908
rect 4406 2892 4409 2948
rect 4398 2872 4401 2878
rect 4422 2872 4425 2958
rect 4486 2952 4489 3058
rect 4558 3052 4561 3118
rect 4566 3072 4569 3078
rect 4522 3048 4526 3051
rect 4526 2992 4529 3038
rect 4574 3032 4577 3118
rect 4582 3052 4585 3058
rect 4558 2982 4561 3028
rect 4558 2972 4561 2978
rect 4574 2972 4577 3018
rect 4510 2962 4513 2968
rect 4550 2952 4553 2958
rect 4462 2932 4465 2938
rect 4454 2882 4457 2918
rect 4470 2882 4473 2928
rect 4486 2892 4489 2948
rect 4522 2938 4534 2941
rect 4546 2938 4550 2941
rect 4518 2932 4521 2938
rect 4558 2902 4561 2958
rect 4566 2942 4569 2948
rect 4394 2858 4398 2861
rect 4238 2762 4241 2798
rect 4414 2792 4417 2848
rect 4306 2758 4310 2761
rect 4238 2752 4241 2758
rect 4262 2752 4265 2758
rect 4234 2738 4238 2741
rect 4038 2692 4041 2728
rect 4080 2703 4082 2707
rect 4086 2703 4089 2707
rect 4093 2703 4096 2707
rect 4126 2702 4129 2718
rect 4038 2682 4041 2688
rect 4026 2678 4030 2681
rect 4018 2668 4022 2671
rect 4050 2668 4054 2671
rect 4090 2668 4094 2671
rect 3990 2658 3998 2661
rect 4054 2652 4057 2658
rect 3962 2648 3966 2651
rect 4066 2648 4070 2651
rect 3918 2608 3929 2611
rect 3918 2592 3921 2608
rect 3926 2562 3929 2568
rect 3942 2562 3945 2648
rect 4062 2622 4065 2638
rect 3958 2562 3961 2618
rect 3974 2562 3977 2618
rect 3942 2552 3945 2558
rect 3910 2542 3913 2548
rect 3850 2538 3854 2541
rect 3930 2538 3934 2541
rect 3962 2538 3966 2541
rect 3978 2538 3982 2541
rect 3646 2522 3649 2528
rect 3694 2491 3697 2528
rect 3702 2522 3705 2528
rect 3690 2488 3697 2491
rect 3634 2478 3638 2481
rect 3686 2472 3689 2478
rect 3642 2468 3646 2471
rect 3662 2462 3665 2468
rect 3694 2462 3697 2468
rect 3702 2462 3705 2498
rect 3718 2492 3721 2518
rect 3742 2492 3745 2528
rect 3750 2512 3753 2518
rect 3782 2502 3785 2538
rect 3822 2532 3825 2538
rect 3894 2532 3897 2538
rect 3966 2522 3969 2528
rect 3814 2492 3817 2518
rect 3750 2472 3753 2478
rect 3782 2472 3785 2478
rect 3814 2472 3817 2488
rect 3834 2478 3838 2481
rect 3862 2472 3865 2518
rect 3902 2482 3905 2518
rect 3890 2478 3894 2481
rect 3938 2478 3942 2481
rect 3834 2468 3838 2471
rect 3522 2458 3526 2461
rect 3334 2452 3337 2458
rect 3358 2452 3361 2458
rect 3306 2448 3310 2451
rect 3330 2448 3334 2451
rect 3346 2448 3350 2451
rect 3322 2438 3326 2441
rect 3302 2432 3305 2438
rect 3358 2392 3361 2398
rect 3346 2388 3350 2391
rect 3302 2362 3305 2388
rect 3366 2372 3369 2458
rect 3646 2452 3649 2458
rect 3670 2452 3673 2458
rect 3442 2448 3446 2451
rect 3658 2448 3662 2451
rect 3714 2448 3718 2451
rect 3726 2451 3729 2468
rect 3766 2462 3769 2468
rect 3790 2462 3793 2468
rect 3942 2462 3945 2468
rect 3810 2458 3814 2461
rect 3722 2448 3729 2451
rect 3746 2448 3750 2451
rect 3778 2448 3782 2451
rect 3850 2448 3854 2451
rect 3414 2442 3417 2448
rect 3494 2432 3497 2448
rect 3398 2412 3401 2418
rect 3202 2358 3206 2361
rect 3234 2358 3238 2361
rect 3258 2348 3262 2351
rect 3302 2342 3305 2348
rect 3310 2342 3313 2358
rect 3350 2352 3353 2358
rect 3374 2352 3377 2368
rect 3470 2362 3473 2388
rect 3406 2352 3409 2358
rect 3486 2352 3489 2368
rect 3510 2352 3513 2378
rect 3526 2362 3529 2438
rect 3546 2378 3550 2381
rect 3558 2362 3561 2428
rect 3568 2403 3570 2407
rect 3574 2403 3577 2407
rect 3581 2403 3584 2407
rect 3742 2392 3745 2448
rect 3798 2442 3801 2448
rect 3854 2442 3857 2448
rect 3634 2378 3638 2381
rect 3670 2362 3673 2378
rect 3634 2358 3638 2361
rect 3714 2358 3718 2361
rect 3522 2348 3526 2351
rect 3546 2348 3550 2351
rect 3234 2338 3238 2341
rect 3266 2338 3270 2341
rect 3350 2342 3353 2348
rect 3454 2342 3457 2348
rect 3206 2332 3209 2338
rect 3318 2332 3321 2340
rect 3434 2338 3438 2341
rect 3366 2332 3369 2338
rect 3274 2328 3278 2331
rect 3102 2272 3105 2328
rect 3098 2268 3102 2271
rect 3122 2258 3126 2261
rect 3102 2252 3105 2258
rect 3134 2252 3137 2318
rect 3150 2312 3153 2328
rect 3174 2302 3177 2328
rect 3214 2291 3217 2318
rect 3206 2288 3217 2291
rect 3206 2282 3209 2288
rect 3238 2282 3241 2318
rect 3246 2292 3249 2298
rect 3254 2282 3257 2318
rect 3302 2292 3305 2308
rect 3218 2278 3222 2281
rect 3274 2278 3278 2281
rect 3298 2278 3305 2281
rect 3150 2272 3153 2278
rect 3170 2268 3174 2271
rect 3194 2268 3198 2271
rect 3290 2268 3294 2271
rect 3142 2262 3145 2268
rect 3186 2258 3190 2261
rect 3158 2252 3161 2258
rect 3182 2252 3185 2258
rect 3114 2248 3118 2251
rect 3170 2248 3174 2251
rect 3230 2242 3233 2258
rect 3266 2248 3270 2251
rect 3182 2192 3185 2218
rect 3230 2192 3233 2198
rect 3134 2182 3137 2188
rect 3118 2172 3121 2178
rect 2994 2138 2998 2141
rect 3026 2138 3030 2141
rect 2946 2128 2950 2131
rect 2894 2112 2897 2128
rect 2878 2082 2881 2108
rect 2894 2072 2897 2108
rect 2934 2102 2937 2128
rect 2958 2102 2961 2128
rect 2966 2092 2969 2138
rect 2982 2122 2985 2128
rect 2938 2078 2942 2081
rect 2950 2072 2953 2088
rect 2854 2062 2857 2068
rect 2878 2062 2881 2068
rect 2950 2062 2953 2068
rect 2790 2058 2801 2061
rect 2544 2003 2546 2007
rect 2550 2003 2553 2007
rect 2557 2003 2560 2007
rect 2630 1982 2633 1988
rect 2514 1958 2518 1961
rect 2630 1958 2638 1961
rect 2518 1942 2521 1958
rect 2530 1948 2534 1951
rect 2510 1881 2513 1918
rect 2510 1878 2521 1881
rect 2370 1868 2374 1871
rect 2422 1862 2425 1868
rect 2478 1862 2481 1878
rect 2486 1862 2489 1878
rect 2518 1872 2521 1878
rect 2450 1858 2454 1861
rect 2270 1848 2278 1851
rect 2318 1851 2321 1858
rect 2486 1852 2489 1858
rect 2510 1852 2513 1868
rect 2318 1848 2329 1851
rect 2246 1832 2249 1848
rect 2262 1842 2265 1848
rect 2254 1822 2257 1828
rect 2094 1792 2097 1808
rect 2138 1768 2142 1771
rect 2030 1732 2033 1738
rect 2118 1732 2121 1738
rect 2126 1732 2129 1768
rect 2134 1731 2137 1748
rect 2150 1732 2153 1808
rect 2158 1742 2161 1788
rect 2174 1762 2177 1768
rect 2198 1762 2201 1798
rect 2270 1792 2273 1848
rect 2290 1838 2294 1841
rect 2230 1762 2233 1768
rect 2174 1742 2177 1748
rect 2182 1742 2185 1758
rect 2198 1742 2201 1758
rect 2214 1752 2217 1758
rect 2234 1748 2238 1751
rect 2246 1742 2249 1758
rect 2318 1752 2321 1758
rect 2274 1748 2278 1751
rect 2190 1732 2193 1738
rect 2254 1732 2257 1738
rect 2262 1732 2265 1748
rect 2314 1738 2318 1741
rect 2326 1732 2329 1848
rect 2434 1848 2438 1851
rect 2382 1762 2385 1768
rect 2390 1762 2393 1818
rect 2342 1752 2345 1758
rect 2406 1742 2409 1788
rect 2414 1742 2417 1818
rect 2422 1752 2425 1848
rect 2430 1761 2433 1818
rect 2446 1762 2449 1768
rect 2470 1762 2473 1818
rect 2430 1758 2438 1761
rect 2486 1752 2489 1838
rect 2358 1732 2361 1738
rect 2366 1732 2369 1738
rect 2130 1728 2137 1731
rect 2146 1728 2150 1731
rect 2242 1728 2246 1731
rect 2298 1728 2302 1731
rect 2330 1728 2334 1731
rect 2078 1722 2081 1728
rect 1866 1718 1870 1721
rect 1986 1718 1990 1721
rect 2330 1718 2334 1721
rect 1846 1691 1849 1718
rect 2286 1712 2289 1718
rect 2024 1703 2026 1707
rect 2030 1703 2033 1707
rect 2037 1703 2040 1707
rect 1846 1688 1857 1691
rect 1890 1688 1894 1691
rect 1726 1652 1729 1658
rect 1734 1642 1737 1648
rect 1694 1592 1697 1638
rect 1702 1592 1705 1618
rect 1742 1612 1745 1658
rect 1790 1652 1793 1678
rect 1798 1672 1801 1678
rect 1814 1672 1817 1688
rect 1846 1672 1849 1678
rect 1854 1672 1857 1688
rect 1982 1682 1985 1698
rect 2042 1688 2046 1691
rect 2170 1688 2174 1691
rect 1970 1678 1974 1681
rect 2114 1678 2118 1681
rect 1902 1672 1905 1678
rect 1930 1668 1934 1671
rect 1986 1668 1990 1671
rect 1830 1652 1833 1668
rect 1854 1652 1857 1668
rect 1878 1652 1881 1668
rect 1910 1652 1913 1658
rect 1766 1642 1769 1648
rect 1774 1642 1777 1648
rect 1830 1642 1833 1648
rect 1886 1642 1889 1648
rect 1682 1548 1689 1551
rect 1654 1532 1657 1538
rect 1678 1522 1681 1548
rect 1694 1522 1697 1528
rect 1710 1512 1713 1548
rect 1718 1542 1721 1588
rect 1718 1532 1721 1538
rect 1698 1488 1702 1491
rect 1646 1462 1649 1488
rect 1654 1472 1657 1478
rect 1662 1472 1665 1478
rect 1698 1468 1702 1471
rect 1726 1462 1729 1578
rect 1758 1552 1761 1638
rect 1766 1552 1769 1558
rect 1750 1542 1753 1548
rect 1742 1492 1745 1518
rect 1746 1478 1750 1481
rect 1706 1458 1710 1461
rect 1646 1432 1649 1438
rect 1646 1392 1649 1418
rect 1678 1382 1681 1448
rect 1590 1352 1593 1358
rect 1598 1342 1601 1368
rect 1678 1352 1681 1378
rect 1630 1332 1633 1338
rect 1662 1332 1665 1348
rect 1670 1342 1673 1348
rect 1586 1328 1590 1331
rect 1558 1282 1561 1318
rect 1582 1302 1585 1328
rect 1606 1322 1609 1328
rect 1630 1282 1633 1328
rect 1650 1288 1654 1291
rect 1574 1272 1577 1278
rect 1614 1272 1617 1278
rect 1618 1258 1622 1261
rect 1566 1162 1569 1218
rect 1574 1192 1577 1258
rect 1606 1252 1609 1258
rect 1630 1252 1633 1268
rect 1638 1262 1641 1268
rect 1666 1258 1670 1261
rect 1586 1248 1590 1251
rect 1650 1248 1654 1251
rect 1594 1238 1598 1241
rect 1598 1152 1601 1188
rect 1606 1182 1609 1248
rect 1614 1232 1617 1248
rect 1606 1142 1609 1168
rect 1510 1138 1518 1141
rect 1446 1132 1449 1138
rect 1482 1118 1486 1121
rect 1358 1068 1369 1071
rect 1406 1072 1409 1078
rect 1342 1042 1345 1068
rect 1350 1062 1353 1068
rect 1358 952 1361 1068
rect 1386 1058 1390 1061
rect 1390 1032 1393 1038
rect 1414 1022 1417 1028
rect 1422 992 1425 1058
rect 1430 1052 1433 1088
rect 1446 1072 1449 1078
rect 1470 1072 1473 1118
rect 1478 1072 1481 1098
rect 1490 1088 1494 1091
rect 1502 1071 1505 1118
rect 1526 1082 1529 1138
rect 1550 1112 1553 1118
rect 1614 1102 1617 1228
rect 1482 1068 1489 1071
rect 1442 1058 1446 1061
rect 1474 1058 1478 1061
rect 1458 1038 1462 1041
rect 1366 952 1369 958
rect 1374 942 1377 978
rect 1430 952 1433 958
rect 1438 952 1441 958
rect 1446 942 1449 978
rect 1470 962 1473 1058
rect 1486 982 1489 1068
rect 1494 1068 1505 1071
rect 1542 1072 1545 1098
rect 1554 1078 1558 1081
rect 1614 1072 1617 1098
rect 1494 1052 1497 1068
rect 1478 952 1481 958
rect 1502 952 1505 1058
rect 1510 992 1513 1058
rect 1520 1003 1522 1007
rect 1526 1003 1529 1007
rect 1533 1003 1536 1007
rect 1542 962 1545 1068
rect 1558 1012 1561 1068
rect 1582 1062 1585 1068
rect 1566 962 1569 968
rect 1490 948 1494 951
rect 1346 938 1350 941
rect 1398 938 1406 941
rect 1314 928 1334 931
rect 1398 922 1401 938
rect 1410 928 1414 931
rect 1462 922 1465 928
rect 1382 892 1385 918
rect 1318 872 1321 878
rect 1194 868 1198 871
rect 1170 858 1174 861
rect 1222 852 1225 868
rect 1186 848 1190 851
rect 1158 751 1161 768
rect 1214 758 1222 761
rect 1206 752 1209 758
rect 1158 748 1169 751
rect 1094 742 1097 748
rect 1166 742 1169 748
rect 1174 742 1177 748
rect 1066 738 1070 741
rect 1154 738 1158 741
rect 1214 741 1217 758
rect 1230 752 1233 858
rect 1238 792 1241 868
rect 1278 862 1281 868
rect 1294 862 1297 868
rect 1326 862 1329 868
rect 1266 848 1270 851
rect 1314 848 1318 851
rect 1206 738 1217 741
rect 1246 742 1249 748
rect 1254 742 1257 748
rect 1270 742 1273 768
rect 1326 742 1329 818
rect 1334 741 1337 888
rect 1350 872 1353 878
rect 1398 872 1401 898
rect 1430 872 1433 878
rect 1454 871 1457 918
rect 1470 912 1473 948
rect 1478 942 1481 948
rect 1494 922 1497 938
rect 1510 912 1513 958
rect 1550 942 1553 948
rect 1518 912 1521 918
rect 1574 902 1577 918
rect 1566 892 1569 898
rect 1582 891 1585 1058
rect 1598 1052 1601 1058
rect 1590 952 1593 1028
rect 1574 888 1585 891
rect 1594 888 1598 891
rect 1470 882 1473 888
rect 1454 868 1462 871
rect 1474 868 1478 871
rect 1350 852 1353 858
rect 1402 848 1406 851
rect 1342 822 1345 848
rect 1422 842 1425 858
rect 1438 852 1441 868
rect 1458 858 1462 861
rect 1366 772 1369 818
rect 1342 762 1345 768
rect 1350 762 1353 768
rect 1370 758 1374 761
rect 1422 752 1425 818
rect 1454 762 1457 818
rect 1446 758 1454 761
rect 1374 742 1377 748
rect 1430 742 1433 758
rect 1446 742 1449 758
rect 1462 751 1465 838
rect 1470 762 1473 768
rect 1462 748 1470 751
rect 1334 738 1342 741
rect 1086 732 1089 738
rect 990 692 993 718
rect 1000 703 1002 707
rect 1006 703 1009 707
rect 1013 703 1016 707
rect 966 672 969 678
rect 894 663 897 668
rect 902 602 905 648
rect 850 568 854 571
rect 798 562 801 568
rect 834 558 838 561
rect 790 548 798 551
rect 774 542 777 548
rect 778 488 782 491
rect 766 468 777 471
rect 698 458 702 461
rect 702 442 705 448
rect 682 438 686 441
rect 694 432 697 438
rect 710 432 713 448
rect 686 342 689 358
rect 702 332 705 428
rect 726 392 729 468
rect 734 382 737 468
rect 766 452 769 458
rect 774 452 777 468
rect 790 462 793 548
rect 802 538 806 541
rect 814 502 817 548
rect 742 362 745 378
rect 790 362 793 378
rect 750 352 753 358
rect 702 312 705 328
rect 726 322 729 348
rect 742 342 745 348
rect 762 338 766 341
rect 786 328 790 331
rect 646 272 649 298
rect 634 268 638 271
rect 654 268 662 271
rect 626 248 630 251
rect 582 162 585 168
rect 462 108 473 111
rect 530 138 534 141
rect 486 122 489 138
rect 550 132 553 158
rect 558 142 561 148
rect 574 142 577 148
rect 598 122 601 138
rect 606 132 609 148
rect 614 142 617 198
rect 638 162 641 268
rect 646 252 649 258
rect 654 192 657 268
rect 678 262 681 298
rect 702 272 705 298
rect 754 288 758 291
rect 698 258 702 261
rect 726 252 729 268
rect 662 212 665 248
rect 718 202 721 248
rect 774 232 777 268
rect 798 262 801 458
rect 814 421 817 458
rect 806 418 817 421
rect 806 392 809 418
rect 806 362 809 388
rect 838 302 841 558
rect 862 552 865 568
rect 874 558 878 561
rect 846 463 849 518
rect 862 402 865 518
rect 878 482 881 558
rect 894 552 897 598
rect 902 572 905 598
rect 902 552 905 558
rect 894 472 897 548
rect 918 542 921 658
rect 986 618 990 621
rect 942 542 945 548
rect 902 472 905 538
rect 890 458 894 461
rect 878 452 881 458
rect 894 442 897 448
rect 862 342 865 398
rect 902 372 905 468
rect 926 442 929 458
rect 934 452 937 478
rect 950 442 953 598
rect 998 562 1001 568
rect 1014 552 1017 688
rect 1022 672 1025 718
rect 1030 712 1033 732
rect 1122 718 1126 721
rect 1038 662 1041 718
rect 1046 672 1049 688
rect 1054 672 1057 678
rect 1062 672 1065 678
rect 1070 672 1073 688
rect 1126 672 1129 708
rect 1142 702 1145 738
rect 1158 712 1161 718
rect 1174 672 1177 708
rect 1182 692 1185 738
rect 1198 732 1201 738
rect 1206 712 1209 738
rect 1246 732 1249 738
rect 1226 728 1230 731
rect 1290 718 1294 721
rect 1194 678 1198 681
rect 1214 672 1217 718
rect 1222 692 1225 708
rect 1238 682 1241 698
rect 1118 662 1121 668
rect 1126 662 1129 668
rect 1198 662 1201 668
rect 1238 662 1241 678
rect 1262 672 1265 718
rect 1302 702 1305 735
rect 1338 728 1342 731
rect 1398 712 1401 718
rect 1290 688 1294 691
rect 1278 675 1282 678
rect 1310 672 1313 688
rect 1318 662 1321 668
rect 1202 658 1209 661
rect 1326 661 1329 698
rect 1398 692 1401 698
rect 1362 678 1366 681
rect 1378 678 1382 681
rect 1422 681 1425 738
rect 1414 678 1425 681
rect 1334 672 1337 678
rect 1342 672 1345 678
rect 1362 668 1366 671
rect 1414 662 1417 678
rect 1422 662 1425 668
rect 1430 662 1433 678
rect 1438 672 1441 698
rect 1462 678 1465 748
rect 1478 742 1481 858
rect 1534 842 1537 868
rect 1558 862 1561 878
rect 1574 872 1577 888
rect 1582 878 1590 881
rect 1594 878 1598 881
rect 1574 862 1577 868
rect 1582 862 1585 878
rect 1606 871 1609 1058
rect 1622 1052 1625 1158
rect 1630 1092 1633 1238
rect 1646 1162 1649 1178
rect 1662 1142 1665 1218
rect 1678 1192 1681 1208
rect 1686 1192 1689 1458
rect 1702 1352 1705 1438
rect 1718 1362 1721 1388
rect 1742 1362 1745 1378
rect 1758 1362 1761 1548
rect 1766 1462 1769 1468
rect 1774 1451 1777 1518
rect 1782 1512 1785 1638
rect 1798 1592 1801 1618
rect 1862 1582 1865 1618
rect 1886 1592 1889 1598
rect 1814 1562 1817 1568
rect 1830 1552 1833 1568
rect 1870 1561 1873 1578
rect 1866 1558 1873 1561
rect 1790 1542 1793 1548
rect 1790 1482 1793 1498
rect 1774 1448 1782 1451
rect 1798 1442 1801 1518
rect 1814 1462 1817 1548
rect 1838 1542 1841 1558
rect 1854 1472 1857 1548
rect 1878 1541 1881 1558
rect 1886 1552 1889 1578
rect 1894 1542 1897 1568
rect 1910 1542 1913 1598
rect 1926 1552 1929 1668
rect 1950 1662 1953 1668
rect 1994 1648 1998 1651
rect 1986 1638 1990 1641
rect 2006 1622 2009 1668
rect 2054 1622 2057 1668
rect 2094 1662 2097 1668
rect 2142 1662 2145 1688
rect 2150 1682 2153 1688
rect 2170 1678 2174 1681
rect 2182 1672 2185 1678
rect 2222 1670 2225 1678
rect 2246 1672 2249 1678
rect 2262 1672 2265 1688
rect 2266 1668 2273 1671
rect 2106 1658 2110 1661
rect 2070 1652 2073 1658
rect 2126 1652 2129 1658
rect 2206 1652 2209 1658
rect 2242 1648 2246 1651
rect 2078 1642 2081 1648
rect 2094 1642 2097 1648
rect 1950 1582 1953 1618
rect 1962 1568 1966 1571
rect 1946 1558 1950 1561
rect 2006 1552 2009 1578
rect 2022 1552 2025 1558
rect 1962 1548 1966 1551
rect 1878 1538 1889 1541
rect 1862 1472 1865 1538
rect 1870 1532 1873 1538
rect 1886 1492 1889 1538
rect 1910 1532 1913 1538
rect 1918 1492 1921 1518
rect 1926 1492 1929 1538
rect 1862 1452 1865 1468
rect 1902 1462 1905 1468
rect 1918 1462 1921 1468
rect 1878 1452 1881 1458
rect 1834 1448 1838 1451
rect 1926 1451 1929 1488
rect 1934 1482 1937 1548
rect 1962 1538 1966 1541
rect 1974 1532 1977 1548
rect 1982 1512 1985 1518
rect 1990 1492 1993 1538
rect 2030 1532 2033 1538
rect 1970 1478 1974 1481
rect 1934 1462 1937 1478
rect 2006 1472 2009 1528
rect 2024 1503 2026 1507
rect 2030 1503 2033 1507
rect 2037 1503 2040 1507
rect 2046 1492 2049 1558
rect 2078 1552 2081 1568
rect 2126 1552 2129 1618
rect 2150 1602 2153 1618
rect 2134 1562 2137 1568
rect 2198 1552 2201 1618
rect 2238 1592 2241 1618
rect 2246 1592 2249 1648
rect 2238 1552 2241 1588
rect 2162 1548 2166 1551
rect 2218 1548 2222 1551
rect 2142 1542 2145 1548
rect 2074 1538 2078 1541
rect 2114 1538 2118 1541
rect 2194 1538 2198 1541
rect 2226 1538 2230 1541
rect 2246 1541 2249 1558
rect 2242 1538 2249 1541
rect 2262 1542 2265 1638
rect 2102 1532 2105 1538
rect 2166 1522 2169 1538
rect 2262 1532 2265 1538
rect 2054 1482 2057 1488
rect 2086 1482 2089 1518
rect 1946 1468 1950 1471
rect 1950 1462 1953 1468
rect 2014 1462 2017 1478
rect 2102 1472 2105 1478
rect 2070 1462 2073 1468
rect 2090 1466 2094 1469
rect 1962 1458 1966 1461
rect 2082 1458 2086 1461
rect 2106 1458 2110 1461
rect 1922 1448 1929 1451
rect 1978 1448 1982 1451
rect 1866 1438 1870 1441
rect 1890 1438 1894 1441
rect 1766 1402 1769 1418
rect 1766 1361 1769 1398
rect 1798 1392 1801 1418
rect 1814 1382 1817 1418
rect 1870 1392 1873 1408
rect 1898 1388 1902 1391
rect 1866 1368 1873 1371
rect 1878 1362 1881 1388
rect 1766 1358 1774 1361
rect 1794 1358 1798 1361
rect 1742 1352 1745 1358
rect 1774 1352 1777 1358
rect 1814 1352 1817 1358
rect 1846 1352 1849 1358
rect 1894 1352 1897 1368
rect 1762 1348 1766 1351
rect 1702 1342 1705 1348
rect 1694 1302 1697 1318
rect 1726 1312 1729 1338
rect 1790 1332 1793 1348
rect 1814 1342 1817 1348
rect 1822 1331 1825 1338
rect 1814 1328 1825 1331
rect 1830 1332 1833 1348
rect 1698 1258 1702 1261
rect 1710 1242 1713 1268
rect 1742 1262 1745 1318
rect 1750 1312 1753 1328
rect 1758 1271 1761 1318
rect 1774 1272 1777 1328
rect 1806 1282 1809 1318
rect 1814 1292 1817 1328
rect 1846 1322 1849 1328
rect 1862 1292 1865 1348
rect 1886 1342 1889 1348
rect 1886 1332 1889 1338
rect 1902 1292 1905 1318
rect 1826 1288 1830 1291
rect 1870 1282 1873 1288
rect 1882 1278 1886 1281
rect 1758 1268 1769 1271
rect 1766 1262 1769 1268
rect 1730 1258 1734 1261
rect 1754 1258 1758 1261
rect 1718 1202 1721 1258
rect 1746 1248 1750 1251
rect 1734 1232 1737 1248
rect 1718 1182 1721 1188
rect 1670 1152 1673 1178
rect 1734 1152 1737 1158
rect 1742 1152 1745 1208
rect 1694 1142 1697 1148
rect 1682 1138 1686 1141
rect 1642 1128 1646 1131
rect 1634 1068 1638 1071
rect 1634 1058 1638 1061
rect 1622 952 1625 1048
rect 1646 1042 1649 1118
rect 1678 1112 1681 1128
rect 1654 1082 1657 1088
rect 1654 1062 1657 1078
rect 1678 1062 1681 1108
rect 1686 1062 1689 1108
rect 1694 1102 1697 1138
rect 1686 1032 1689 1058
rect 1670 982 1673 1018
rect 1694 962 1697 1018
rect 1702 972 1705 1148
rect 1710 1052 1713 1058
rect 1726 1052 1729 1058
rect 1670 952 1673 958
rect 1710 952 1713 998
rect 1726 952 1729 958
rect 1690 948 1694 951
rect 1614 932 1617 948
rect 1710 942 1713 948
rect 1658 938 1662 941
rect 1722 938 1726 941
rect 1630 872 1633 908
rect 1638 902 1641 918
rect 1598 868 1609 871
rect 1618 868 1622 871
rect 1642 868 1646 871
rect 1506 818 1510 821
rect 1520 803 1522 807
rect 1526 803 1529 807
rect 1533 803 1536 807
rect 1478 702 1481 738
rect 1486 732 1489 768
rect 1494 672 1497 678
rect 1326 658 1334 661
rect 1158 652 1161 658
rect 1098 618 1102 621
rect 1134 592 1137 618
rect 1150 592 1153 608
rect 1070 551 1073 578
rect 966 542 969 548
rect 1102 542 1105 548
rect 1142 532 1145 538
rect 1158 531 1161 558
rect 1166 542 1169 548
rect 1158 528 1169 531
rect 1000 503 1002 507
rect 1006 503 1009 507
rect 1013 503 1016 507
rect 958 462 961 468
rect 982 442 985 448
rect 914 438 918 441
rect 902 352 905 358
rect 926 352 929 418
rect 810 268 814 271
rect 782 252 785 258
rect 830 252 833 258
rect 838 252 841 298
rect 846 272 849 288
rect 854 282 857 338
rect 874 318 881 321
rect 854 262 857 278
rect 870 252 873 288
rect 798 242 801 248
rect 818 238 822 241
rect 814 191 817 218
rect 806 188 817 191
rect 846 192 849 248
rect 878 222 881 318
rect 934 272 937 368
rect 906 268 910 271
rect 890 258 894 261
rect 922 258 926 261
rect 950 261 953 438
rect 1006 351 1009 378
rect 1014 322 1017 459
rect 1030 352 1033 468
rect 1000 303 1002 307
rect 1006 303 1009 307
rect 1013 303 1016 307
rect 942 258 953 261
rect 930 248 934 251
rect 894 242 897 248
rect 678 162 681 188
rect 622 152 625 158
rect 630 152 633 158
rect 702 152 705 188
rect 650 148 654 151
rect 718 142 721 148
rect 642 138 646 141
rect 698 138 702 141
rect 706 128 710 131
rect 450 88 454 91
rect 406 72 409 78
rect 310 58 313 59
rect 354 58 358 61
rect 394 59 398 62
rect 462 62 465 108
rect 486 62 489 118
rect 518 62 521 88
rect 6 42 9 48
rect 102 -19 105 18
rect 110 -19 114 -18
rect 102 -22 114 -19
rect 222 -19 225 18
rect 230 -19 234 -18
rect 222 -22 234 -19
rect 342 -19 345 18
rect 350 -19 354 -18
rect 342 -22 354 -19
rect 470 -19 474 -18
rect 478 -19 481 18
rect 470 -22 481 -19
rect 486 -19 489 18
rect 496 3 498 7
rect 502 3 505 7
rect 509 3 512 7
rect 518 -19 522 -18
rect 486 -22 522 -19
rect 526 -19 529 118
rect 574 72 577 78
rect 622 62 625 128
rect 734 92 737 98
rect 654 72 657 78
rect 578 58 582 61
rect 626 58 630 61
rect 674 59 678 62
rect 742 62 745 118
rect 758 62 761 178
rect 806 151 809 188
rect 858 168 862 171
rect 902 152 905 158
rect 774 112 777 148
rect 850 148 854 151
rect 910 151 913 238
rect 942 172 945 258
rect 958 251 961 298
rect 1038 282 1041 518
rect 1094 462 1097 468
rect 1110 442 1113 459
rect 1166 442 1169 528
rect 1174 492 1177 658
rect 1206 492 1209 658
rect 1382 652 1385 658
rect 1406 652 1409 658
rect 1262 551 1265 568
rect 1222 522 1225 538
rect 1246 532 1249 538
rect 1222 472 1225 518
rect 1270 492 1273 628
rect 1326 592 1329 618
rect 1350 552 1353 618
rect 1390 592 1393 638
rect 1486 592 1489 668
rect 1502 662 1505 728
rect 1470 582 1473 588
rect 1382 562 1385 568
rect 1390 552 1393 578
rect 1366 532 1369 548
rect 1330 528 1334 531
rect 1342 502 1345 518
rect 1382 512 1385 518
rect 1278 472 1281 498
rect 1326 472 1329 478
rect 1382 472 1385 478
rect 1390 472 1393 498
rect 1334 462 1337 468
rect 1398 462 1401 578
rect 1442 568 1446 571
rect 1474 568 1478 571
rect 1502 571 1505 618
rect 1494 568 1505 571
rect 1510 572 1513 718
rect 1518 652 1521 768
rect 1546 728 1550 731
rect 1558 692 1561 858
rect 1566 752 1569 758
rect 1574 742 1577 858
rect 1598 792 1601 868
rect 1670 862 1673 928
rect 1686 892 1689 938
rect 1734 922 1737 938
rect 1742 932 1745 1148
rect 1758 1101 1761 1218
rect 1782 1172 1785 1218
rect 1798 1162 1801 1258
rect 1806 1252 1809 1278
rect 1822 1252 1825 1278
rect 1902 1272 1905 1288
rect 1910 1282 1913 1448
rect 2030 1442 2033 1448
rect 1918 1362 1921 1368
rect 1922 1348 1929 1351
rect 1918 1322 1921 1328
rect 1926 1322 1929 1348
rect 1934 1332 1937 1348
rect 1866 1268 1870 1271
rect 1890 1268 1894 1271
rect 1922 1268 1926 1271
rect 1838 1262 1841 1268
rect 1858 1258 1862 1261
rect 1838 1252 1841 1258
rect 1886 1222 1889 1258
rect 1894 1232 1897 1238
rect 1766 1142 1769 1148
rect 1750 1098 1761 1101
rect 1750 1082 1753 1098
rect 1762 1088 1766 1091
rect 1774 1082 1777 1158
rect 1790 1142 1793 1148
rect 1790 1112 1793 1138
rect 1762 1048 1766 1051
rect 1750 932 1753 978
rect 1766 952 1769 1018
rect 1774 992 1777 1068
rect 1782 1062 1785 1088
rect 1790 1072 1793 1088
rect 1798 1082 1801 1158
rect 1810 1148 1814 1151
rect 1782 982 1785 1018
rect 1770 948 1774 951
rect 1698 918 1702 921
rect 1766 892 1769 938
rect 1782 932 1785 938
rect 1682 878 1686 881
rect 1758 872 1761 878
rect 1730 868 1734 871
rect 1702 862 1705 868
rect 1634 858 1638 861
rect 1738 858 1742 861
rect 1606 781 1609 858
rect 1622 852 1625 858
rect 1694 792 1697 848
rect 1718 842 1721 848
rect 1726 842 1729 848
rect 1598 778 1609 781
rect 1578 728 1582 731
rect 1520 603 1522 607
rect 1526 603 1529 607
rect 1533 603 1536 607
rect 1550 592 1553 678
rect 1562 668 1566 671
rect 1570 658 1574 661
rect 1486 552 1489 568
rect 1494 562 1497 568
rect 1510 561 1513 568
rect 1506 558 1513 561
rect 1494 552 1497 558
rect 1414 542 1417 548
rect 1518 542 1521 548
rect 1558 542 1561 568
rect 1598 562 1601 778
rect 1606 752 1609 758
rect 1654 752 1657 758
rect 1694 752 1697 778
rect 1618 738 1622 741
rect 1642 738 1646 741
rect 1682 738 1686 741
rect 1662 732 1665 738
rect 1622 722 1625 728
rect 1626 688 1630 691
rect 1646 682 1649 688
rect 1614 672 1617 678
rect 1654 672 1657 718
rect 1662 692 1665 728
rect 1670 672 1673 728
rect 1678 692 1681 728
rect 1682 678 1686 681
rect 1634 668 1638 671
rect 1694 662 1697 708
rect 1642 658 1646 661
rect 1606 632 1609 658
rect 1630 592 1633 658
rect 1654 572 1657 618
rect 1702 582 1705 818
rect 1714 758 1718 761
rect 1722 748 1726 751
rect 1734 732 1737 848
rect 1742 752 1745 858
rect 1750 852 1753 868
rect 1782 852 1785 858
rect 1790 852 1793 948
rect 1798 942 1801 958
rect 1798 842 1801 878
rect 1806 782 1809 1138
rect 1814 991 1817 1148
rect 1822 1092 1825 1178
rect 1838 1152 1841 1168
rect 1846 1142 1849 1148
rect 1834 1128 1838 1131
rect 1846 1092 1849 1138
rect 1846 1062 1849 1078
rect 1854 1062 1857 1218
rect 1870 1162 1873 1168
rect 1878 1142 1881 1148
rect 1886 1132 1889 1188
rect 1894 1162 1897 1178
rect 1894 1142 1897 1148
rect 1870 1112 1873 1118
rect 1886 1082 1889 1128
rect 1902 1092 1905 1268
rect 1934 1262 1937 1328
rect 1942 1312 1945 1348
rect 1958 1332 1961 1418
rect 1974 1392 1977 1438
rect 1990 1372 1993 1418
rect 1950 1322 1953 1328
rect 1942 1272 1945 1308
rect 1910 1152 1913 1258
rect 1918 1142 1921 1248
rect 1926 1222 1929 1228
rect 1950 1222 1953 1278
rect 1958 1252 1961 1298
rect 1966 1292 1969 1338
rect 1974 1332 1977 1348
rect 1990 1322 1993 1358
rect 2014 1352 2017 1368
rect 2002 1328 2006 1331
rect 2006 1282 2009 1318
rect 1974 1272 1977 1278
rect 1990 1252 1993 1258
rect 1926 1182 1929 1198
rect 1926 1142 1929 1178
rect 1934 1152 1937 1158
rect 1918 1132 1921 1138
rect 1918 1092 1921 1118
rect 1830 1052 1833 1058
rect 1846 1042 1849 1058
rect 1858 1048 1862 1051
rect 1814 988 1825 991
rect 1814 972 1817 978
rect 1822 952 1825 988
rect 1830 952 1833 1008
rect 1838 1002 1841 1018
rect 1870 992 1873 1078
rect 1898 1068 1902 1071
rect 1926 1062 1929 1078
rect 1934 1072 1937 1078
rect 1930 1058 1934 1061
rect 1878 1032 1881 1038
rect 1886 1032 1889 1058
rect 1886 992 1889 998
rect 1942 992 1945 1188
rect 1950 1162 1953 1218
rect 1958 1162 1961 1248
rect 1954 1148 1958 1151
rect 1966 1142 1969 1148
rect 1954 1128 1958 1131
rect 1974 1092 1977 1208
rect 1982 1192 1985 1238
rect 1998 1182 2001 1188
rect 1982 1112 1985 1128
rect 1990 1102 1993 1138
rect 1998 1082 2001 1128
rect 1986 1068 1990 1071
rect 1998 1062 2001 1078
rect 1958 1052 1961 1058
rect 1998 992 2001 1008
rect 1846 962 1849 968
rect 1854 952 1857 988
rect 1882 968 1886 971
rect 1902 962 1905 988
rect 1938 968 1942 971
rect 2006 962 2009 1218
rect 2014 1192 2017 1328
rect 2046 1322 2049 1348
rect 2024 1303 2026 1307
rect 2030 1303 2033 1307
rect 2037 1303 2040 1307
rect 2054 1272 2057 1458
rect 2126 1432 2129 1478
rect 2142 1462 2145 1478
rect 2150 1472 2153 1518
rect 2174 1512 2177 1518
rect 2190 1492 2193 1508
rect 2206 1492 2209 1518
rect 2246 1512 2249 1518
rect 2174 1472 2177 1478
rect 2154 1468 2158 1471
rect 2210 1468 2214 1471
rect 2214 1462 2217 1468
rect 2222 1462 2225 1468
rect 2146 1458 2150 1461
rect 2194 1458 2198 1461
rect 2158 1451 2161 1458
rect 2222 1452 2225 1458
rect 2154 1448 2161 1451
rect 2206 1442 2209 1448
rect 2194 1438 2198 1441
rect 2226 1438 2230 1441
rect 2070 1362 2073 1368
rect 2102 1362 2105 1398
rect 2110 1362 2113 1378
rect 2166 1372 2169 1408
rect 2178 1388 2182 1391
rect 2198 1362 2201 1368
rect 2146 1358 2150 1361
rect 2062 1332 2065 1358
rect 2138 1348 2142 1351
rect 2154 1348 2158 1351
rect 2182 1342 2185 1358
rect 2214 1352 2217 1378
rect 2238 1352 2241 1488
rect 2270 1482 2273 1668
rect 2278 1662 2281 1698
rect 2342 1692 2345 1718
rect 2302 1662 2305 1688
rect 2350 1682 2353 1718
rect 2382 1702 2385 1718
rect 2310 1662 2313 1668
rect 2350 1662 2353 1668
rect 2358 1652 2361 1698
rect 2378 1668 2382 1671
rect 2390 1662 2393 1718
rect 2422 1672 2425 1748
rect 2466 1738 2470 1741
rect 2490 1738 2494 1741
rect 2502 1732 2505 1828
rect 2526 1792 2529 1858
rect 2534 1802 2537 1928
rect 2542 1892 2545 1958
rect 2618 1940 2622 1943
rect 2562 1928 2566 1931
rect 2598 1912 2601 1928
rect 2566 1882 2569 1888
rect 2606 1882 2609 1938
rect 2602 1858 2606 1861
rect 2554 1848 2558 1851
rect 2594 1848 2598 1851
rect 2614 1842 2617 1940
rect 2622 1882 2625 1908
rect 2630 1892 2633 1958
rect 2654 1922 2657 1938
rect 2662 1932 2665 2018
rect 2674 1958 2678 1961
rect 2682 1948 2686 1951
rect 2670 1942 2673 1948
rect 2638 1912 2641 1918
rect 2630 1882 2633 1888
rect 2630 1872 2633 1878
rect 2662 1872 2665 1878
rect 2686 1862 2689 1928
rect 2694 1882 2697 1948
rect 2702 1942 2705 2018
rect 2710 1942 2713 1948
rect 2726 1944 2729 2008
rect 2750 1982 2753 1988
rect 2766 1952 2769 2028
rect 2798 1992 2801 2058
rect 2814 2052 2817 2058
rect 2894 2052 2897 2058
rect 2918 2052 2921 2058
rect 2858 2048 2862 2051
rect 2870 2032 2873 2048
rect 2926 2041 2929 2048
rect 2914 2038 2929 2041
rect 2934 2042 2937 2058
rect 2946 2048 2950 2051
rect 2974 2032 2977 2078
rect 3006 2072 3009 2118
rect 3038 2092 3041 2118
rect 3048 2103 3050 2107
rect 3054 2103 3057 2107
rect 3061 2103 3064 2107
rect 3070 2092 3073 2148
rect 3078 2142 3081 2148
rect 3102 2122 3105 2158
rect 3110 2132 3113 2148
rect 3122 2128 3126 2131
rect 3094 2102 3097 2118
rect 3118 2092 3121 2118
rect 3134 2112 3137 2148
rect 3134 2092 3137 2108
rect 3046 2082 3049 2088
rect 3102 2082 3105 2088
rect 3134 2082 3137 2088
rect 2986 2068 2990 2071
rect 3078 2062 3081 2078
rect 3094 2068 3102 2071
rect 3094 2062 3097 2068
rect 3106 2058 3110 2061
rect 3014 2052 3017 2058
rect 2810 2028 2814 2031
rect 3022 2022 3025 2058
rect 2838 1952 2841 1958
rect 2862 1952 2865 1978
rect 2878 1952 2881 2008
rect 2886 1992 2889 2018
rect 2722 1940 2726 1943
rect 2742 1941 2745 1948
rect 2766 1942 2769 1948
rect 2726 1938 2729 1940
rect 2742 1938 2753 1941
rect 2750 1932 2753 1938
rect 2798 1932 2801 1948
rect 2854 1932 2857 1938
rect 2878 1932 2881 1948
rect 2886 1942 2889 1948
rect 2738 1928 2742 1931
rect 2842 1928 2846 1931
rect 2886 1922 2889 1928
rect 2650 1838 2654 1841
rect 2674 1838 2678 1841
rect 2544 1803 2546 1807
rect 2550 1803 2553 1807
rect 2557 1803 2560 1807
rect 2534 1762 2537 1798
rect 2514 1728 2518 1731
rect 2450 1718 2454 1721
rect 2430 1682 2433 1688
rect 2398 1662 2401 1668
rect 2286 1602 2289 1618
rect 2278 1562 2281 1568
rect 2294 1562 2297 1578
rect 2286 1551 2289 1558
rect 2318 1552 2321 1558
rect 2282 1548 2289 1551
rect 2294 1542 2297 1548
rect 2278 1532 2281 1538
rect 2310 1532 2313 1538
rect 2318 1521 2321 1538
rect 2310 1518 2321 1521
rect 2246 1422 2249 1478
rect 2258 1468 2262 1471
rect 2278 1462 2281 1518
rect 2286 1512 2289 1518
rect 2290 1478 2294 1481
rect 2302 1472 2305 1508
rect 2266 1458 2270 1461
rect 2310 1452 2313 1518
rect 2326 1512 2329 1618
rect 2390 1592 2393 1638
rect 2366 1552 2369 1578
rect 2382 1552 2385 1558
rect 2390 1552 2393 1588
rect 2398 1562 2401 1618
rect 2414 1552 2417 1558
rect 2342 1542 2345 1548
rect 2350 1542 2353 1548
rect 2394 1538 2398 1541
rect 2358 1532 2361 1538
rect 2338 1518 2342 1521
rect 2350 1472 2353 1498
rect 2318 1462 2321 1468
rect 2342 1462 2345 1468
rect 2362 1458 2366 1461
rect 2326 1452 2329 1458
rect 2314 1448 2318 1451
rect 2354 1448 2358 1451
rect 2342 1442 2345 1448
rect 2382 1441 2385 1518
rect 2390 1462 2393 1508
rect 2414 1492 2417 1548
rect 2422 1442 2425 1638
rect 2430 1622 2433 1658
rect 2438 1592 2441 1718
rect 2470 1682 2473 1718
rect 2494 1682 2497 1728
rect 2502 1691 2505 1728
rect 2502 1688 2513 1691
rect 2450 1678 2454 1681
rect 2438 1531 2441 1558
rect 2430 1528 2441 1531
rect 2430 1522 2433 1528
rect 2438 1492 2441 1518
rect 2446 1472 2449 1678
rect 2454 1652 2457 1668
rect 2502 1662 2505 1678
rect 2510 1672 2513 1688
rect 2518 1672 2521 1688
rect 2534 1672 2537 1728
rect 2566 1682 2569 1818
rect 2574 1732 2577 1808
rect 2614 1772 2617 1818
rect 2646 1772 2649 1798
rect 2666 1768 2670 1771
rect 2582 1702 2585 1748
rect 2590 1742 2593 1758
rect 2646 1752 2649 1768
rect 2686 1762 2689 1818
rect 2694 1802 2697 1858
rect 2702 1852 2705 1918
rect 2734 1892 2737 1908
rect 2866 1888 2870 1891
rect 2710 1862 2713 1888
rect 2742 1872 2745 1878
rect 2766 1872 2769 1878
rect 2774 1862 2777 1878
rect 2798 1872 2801 1888
rect 2878 1872 2881 1878
rect 2894 1871 2897 1998
rect 3086 1992 3089 2018
rect 3142 2002 3145 2178
rect 3150 2152 3153 2168
rect 3246 2162 3249 2168
rect 3202 2158 3209 2161
rect 3182 2142 3185 2148
rect 3158 2138 3166 2141
rect 3158 2132 3161 2138
rect 3170 2128 3174 2131
rect 3158 2102 3161 2118
rect 3198 2092 3201 2158
rect 3206 2132 3209 2158
rect 3226 2148 3230 2151
rect 3254 2151 3257 2248
rect 3262 2192 3265 2218
rect 3270 2162 3273 2168
rect 3246 2148 3257 2151
rect 3218 2138 3222 2141
rect 3214 2102 3217 2118
rect 3206 2082 3209 2098
rect 3214 2082 3217 2088
rect 3238 2082 3241 2098
rect 3246 2092 3249 2148
rect 3254 2132 3257 2138
rect 3270 2132 3273 2138
rect 3278 2132 3281 2138
rect 3294 2092 3297 2238
rect 3302 2222 3305 2278
rect 3310 2272 3313 2278
rect 3334 2272 3337 2318
rect 3374 2292 3377 2328
rect 3382 2302 3385 2338
rect 3398 2332 3401 2338
rect 3434 2328 3438 2331
rect 3390 2281 3393 2318
rect 3406 2282 3409 2298
rect 3454 2292 3457 2328
rect 3478 2292 3481 2348
rect 3502 2332 3505 2338
rect 3390 2278 3401 2281
rect 3434 2278 3438 2281
rect 3362 2268 3366 2271
rect 3310 2258 3318 2261
rect 3330 2258 3334 2261
rect 3302 2152 3305 2178
rect 3310 2092 3313 2258
rect 3318 2251 3321 2258
rect 3318 2248 3326 2251
rect 3334 2231 3337 2258
rect 3342 2242 3345 2248
rect 3358 2242 3361 2248
rect 3334 2228 3345 2231
rect 3334 2171 3337 2218
rect 3326 2168 3337 2171
rect 3318 2142 3321 2148
rect 3326 2142 3329 2168
rect 3334 2132 3337 2148
rect 3318 2122 3321 2128
rect 3278 2082 3281 2088
rect 3246 2068 3254 2071
rect 3150 2052 3153 2068
rect 3174 2052 3177 2068
rect 3182 2062 3185 2068
rect 3190 2062 3193 2068
rect 3218 2058 3222 2061
rect 3230 2052 3233 2058
rect 3246 2032 3249 2068
rect 3258 2058 3262 2061
rect 3286 2052 3289 2058
rect 3182 1992 3185 2028
rect 3010 1988 3014 1991
rect 2914 1958 2918 1961
rect 2902 1942 2905 1948
rect 2938 1938 2942 1941
rect 2938 1928 2942 1931
rect 2906 1878 2918 1881
rect 2938 1878 2942 1881
rect 2890 1868 2897 1871
rect 2786 1858 2790 1861
rect 2718 1842 2721 1848
rect 2710 1812 2713 1818
rect 2606 1742 2609 1748
rect 2614 1742 2617 1748
rect 2618 1738 2625 1741
rect 2622 1732 2625 1738
rect 2630 1732 2633 1738
rect 2594 1728 2598 1731
rect 2638 1702 2641 1738
rect 2654 1732 2657 1748
rect 2662 1742 2665 1758
rect 2694 1752 2697 1798
rect 2718 1752 2721 1838
rect 2750 1832 2753 1848
rect 2790 1842 2793 1848
rect 2678 1742 2681 1748
rect 2686 1712 2689 1748
rect 2726 1742 2729 1748
rect 2734 1742 2737 1748
rect 2702 1732 2705 1738
rect 2750 1732 2753 1828
rect 2766 1792 2769 1798
rect 2770 1748 2774 1751
rect 2622 1682 2625 1688
rect 2678 1682 2681 1688
rect 2590 1662 2593 1668
rect 2614 1662 2617 1678
rect 2634 1668 2638 1671
rect 2622 1662 2625 1668
rect 2654 1662 2657 1678
rect 2694 1662 2697 1678
rect 2474 1658 2478 1661
rect 2534 1652 2537 1658
rect 2702 1652 2705 1728
rect 2718 1712 2721 1728
rect 2734 1718 2742 1721
rect 2714 1668 2718 1671
rect 2718 1652 2721 1668
rect 2554 1648 2558 1651
rect 2586 1618 2590 1621
rect 2642 1618 2646 1621
rect 2462 1602 2465 1618
rect 2544 1603 2546 1607
rect 2550 1603 2553 1607
rect 2557 1603 2560 1607
rect 2478 1552 2481 1558
rect 2494 1552 2497 1588
rect 2526 1562 2529 1568
rect 2454 1542 2457 1548
rect 2470 1532 2473 1548
rect 2486 1542 2489 1548
rect 2522 1538 2526 1541
rect 2466 1468 2470 1471
rect 2502 1462 2505 1538
rect 2510 1462 2513 1518
rect 2378 1438 2385 1441
rect 2406 1432 2409 1438
rect 2278 1412 2281 1418
rect 2366 1412 2369 1418
rect 2262 1352 2265 1358
rect 2278 1352 2281 1358
rect 2130 1338 2142 1341
rect 2202 1338 2206 1341
rect 2026 1268 2030 1271
rect 2022 1152 2025 1248
rect 2030 1172 2033 1268
rect 2038 1172 2041 1218
rect 2062 1152 2065 1318
rect 2070 1282 2073 1328
rect 2102 1292 2105 1318
rect 2110 1282 2113 1318
rect 2150 1292 2153 1318
rect 2118 1272 2121 1278
rect 2126 1272 2129 1288
rect 2106 1268 2110 1271
rect 2098 1258 2102 1261
rect 2074 1248 2078 1251
rect 2094 1242 2097 1248
rect 2118 1192 2121 1258
rect 2134 1212 2137 1218
rect 2050 1148 2054 1151
rect 2086 1142 2089 1148
rect 2118 1142 2121 1148
rect 2106 1138 2110 1141
rect 2022 1132 2025 1138
rect 2058 1128 2062 1131
rect 2106 1128 2110 1131
rect 2024 1103 2026 1107
rect 2030 1103 2033 1107
rect 2037 1103 2040 1107
rect 2134 1092 2137 1158
rect 2142 1142 2145 1288
rect 2190 1282 2193 1318
rect 2218 1278 2222 1281
rect 2154 1268 2158 1271
rect 2166 1262 2169 1278
rect 2230 1272 2233 1318
rect 2246 1302 2249 1338
rect 2262 1332 2265 1338
rect 2262 1302 2265 1318
rect 2262 1292 2265 1298
rect 2254 1272 2257 1278
rect 2190 1262 2193 1268
rect 2202 1258 2206 1261
rect 2166 1162 2169 1258
rect 2190 1202 2193 1248
rect 2198 1242 2201 1248
rect 2214 1242 2217 1268
rect 2242 1266 2246 1269
rect 2230 1252 2233 1258
rect 2278 1252 2281 1348
rect 2294 1332 2297 1378
rect 2338 1358 2342 1361
rect 2294 1281 2297 1328
rect 2290 1278 2297 1281
rect 2302 1262 2305 1358
rect 2318 1332 2321 1338
rect 2326 1322 2329 1348
rect 2350 1342 2353 1378
rect 2358 1332 2361 1348
rect 2266 1248 2270 1251
rect 2162 1158 2166 1161
rect 2170 1148 2174 1151
rect 2158 1142 2161 1148
rect 2182 1142 2185 1188
rect 2214 1162 2217 1188
rect 2222 1162 2225 1228
rect 2238 1152 2241 1208
rect 2286 1192 2289 1258
rect 2310 1212 2313 1318
rect 2318 1252 2321 1258
rect 2334 1252 2337 1318
rect 2346 1288 2350 1291
rect 2358 1281 2361 1328
rect 2366 1312 2369 1338
rect 2382 1332 2385 1418
rect 2422 1362 2425 1438
rect 2430 1392 2433 1458
rect 2446 1412 2449 1418
rect 2454 1402 2457 1458
rect 2462 1452 2465 1458
rect 2478 1452 2481 1458
rect 2486 1392 2489 1398
rect 2462 1362 2465 1368
rect 2434 1358 2438 1361
rect 2390 1352 2393 1358
rect 2402 1348 2406 1351
rect 2418 1348 2422 1351
rect 2466 1348 2470 1351
rect 2410 1338 2414 1341
rect 2390 1332 2393 1338
rect 2406 1282 2409 1328
rect 2438 1312 2441 1348
rect 2446 1332 2449 1338
rect 2470 1332 2473 1338
rect 2478 1292 2481 1358
rect 2486 1332 2489 1388
rect 2494 1362 2497 1368
rect 2498 1348 2502 1351
rect 2446 1282 2449 1288
rect 2494 1282 2497 1348
rect 2510 1332 2513 1418
rect 2526 1392 2529 1458
rect 2534 1452 2537 1558
rect 2542 1542 2545 1578
rect 2570 1548 2574 1551
rect 2574 1492 2577 1538
rect 2554 1468 2558 1471
rect 2518 1332 2521 1378
rect 2526 1352 2529 1358
rect 2510 1312 2513 1318
rect 2526 1292 2529 1328
rect 2358 1278 2369 1281
rect 2342 1252 2345 1278
rect 2258 1158 2262 1161
rect 2270 1152 2273 1158
rect 2154 1118 2158 1121
rect 2190 1112 2193 1148
rect 2214 1142 2217 1148
rect 2050 1078 2054 1081
rect 2018 1068 2022 1071
rect 2090 1068 2094 1071
rect 2082 1058 2086 1061
rect 1890 958 1894 961
rect 1830 942 1833 948
rect 1818 928 1822 931
rect 1814 862 1817 878
rect 1838 862 1841 908
rect 1846 862 1849 948
rect 1886 932 1889 948
rect 1918 942 1921 948
rect 1942 932 1945 948
rect 1910 922 1913 928
rect 1870 902 1873 918
rect 1870 892 1873 898
rect 1930 878 1934 881
rect 1854 872 1857 878
rect 1890 868 1894 871
rect 1814 792 1817 848
rect 1886 842 1889 858
rect 1902 832 1905 878
rect 1950 871 1953 958
rect 1982 952 1985 958
rect 1986 928 1990 931
rect 1966 922 1969 928
rect 1958 882 1961 898
rect 1966 892 1969 908
rect 1950 868 1961 871
rect 1910 842 1913 868
rect 1934 862 1937 868
rect 1946 858 1950 861
rect 1950 842 1953 848
rect 1794 758 1798 761
rect 1750 752 1753 758
rect 1774 752 1777 758
rect 1814 752 1817 758
rect 1822 752 1825 818
rect 1886 772 1889 798
rect 1894 792 1897 798
rect 1830 752 1833 768
rect 1762 748 1766 751
rect 1790 742 1793 748
rect 1770 738 1777 741
rect 1730 728 1734 731
rect 1746 728 1750 731
rect 1734 722 1737 728
rect 1726 702 1729 718
rect 1718 662 1721 688
rect 1726 672 1729 698
rect 1734 672 1737 708
rect 1750 681 1753 718
rect 1766 692 1769 728
rect 1774 692 1777 738
rect 1782 682 1785 738
rect 1822 702 1825 738
rect 1830 732 1833 738
rect 1846 732 1849 748
rect 1854 732 1857 738
rect 1746 678 1753 681
rect 1742 662 1745 678
rect 1750 662 1753 668
rect 1758 652 1761 678
rect 1798 672 1801 698
rect 1806 662 1809 688
rect 1846 681 1849 728
rect 1870 692 1873 758
rect 1902 752 1905 758
rect 1958 752 1961 868
rect 1974 812 1977 868
rect 1966 752 1969 758
rect 1922 748 1926 751
rect 1878 742 1881 748
rect 1902 712 1905 748
rect 1934 742 1937 748
rect 1846 678 1857 681
rect 1854 672 1857 678
rect 1890 668 1894 671
rect 1778 658 1782 661
rect 1822 652 1825 668
rect 1846 662 1849 668
rect 1718 642 1721 648
rect 1770 638 1774 641
rect 1790 622 1793 648
rect 1702 562 1705 568
rect 1658 558 1662 561
rect 1582 552 1585 558
rect 1410 528 1414 531
rect 1430 492 1433 498
rect 1206 452 1209 459
rect 1414 452 1417 478
rect 1442 468 1457 471
rect 1074 438 1078 441
rect 1102 351 1105 388
rect 1134 342 1137 348
rect 1074 318 1078 321
rect 1158 301 1161 438
rect 1166 392 1169 428
rect 1202 348 1206 351
rect 1294 351 1297 438
rect 1354 418 1358 421
rect 1302 412 1305 418
rect 1230 342 1233 348
rect 1310 342 1313 348
rect 1266 318 1270 321
rect 1158 298 1169 301
rect 1166 292 1169 298
rect 1058 288 1062 291
rect 1166 282 1169 288
rect 1262 282 1265 288
rect 970 268 974 271
rect 1066 268 1070 271
rect 978 258 982 261
rect 1010 258 1014 261
rect 1042 258 1046 261
rect 958 248 966 251
rect 950 242 953 248
rect 1030 242 1033 258
rect 1042 248 1046 251
rect 958 231 961 238
rect 950 228 961 231
rect 950 192 953 228
rect 958 182 961 218
rect 930 158 934 161
rect 950 152 953 158
rect 910 148 918 151
rect 774 82 777 108
rect 790 92 793 118
rect 838 102 841 148
rect 782 62 785 88
rect 806 72 809 78
rect 846 72 849 108
rect 870 82 873 148
rect 878 132 881 138
rect 894 112 897 128
rect 826 58 830 61
rect 866 59 870 62
rect 894 62 897 108
rect 958 92 961 148
rect 974 112 977 118
rect 930 88 934 91
rect 934 62 937 78
rect 958 62 961 68
rect 982 62 985 218
rect 998 162 1001 238
rect 1054 222 1057 248
rect 1038 182 1041 218
rect 1070 182 1073 268
rect 1086 262 1089 268
rect 1102 262 1105 278
rect 1310 272 1313 338
rect 1134 262 1137 268
rect 1166 263 1169 268
rect 1114 258 1118 261
rect 1274 258 1278 261
rect 1078 192 1081 258
rect 1030 152 1033 178
rect 1086 172 1089 238
rect 1082 168 1086 171
rect 1094 152 1097 258
rect 1106 248 1110 251
rect 1230 242 1233 258
rect 1122 238 1126 241
rect 1230 232 1233 238
rect 1102 162 1105 168
rect 1090 148 1094 151
rect 1014 122 1017 148
rect 1106 138 1110 141
rect 1158 132 1161 138
rect 1000 103 1002 107
rect 1006 103 1009 107
rect 1013 103 1016 107
rect 1046 82 1049 128
rect 1110 92 1113 128
rect 1110 82 1113 88
rect 1134 62 1137 118
rect 1166 63 1169 208
rect 1174 152 1177 178
rect 1238 162 1241 188
rect 1218 158 1222 161
rect 1182 152 1185 158
rect 1174 142 1177 148
rect 1198 112 1201 158
rect 1294 152 1297 268
rect 1318 202 1321 418
rect 1398 402 1401 418
rect 1366 342 1369 398
rect 1414 342 1417 358
rect 1422 352 1425 468
rect 1454 462 1457 468
rect 1462 462 1465 538
rect 1570 528 1574 531
rect 1470 472 1473 508
rect 1478 472 1481 528
rect 1486 482 1489 528
rect 1502 492 1505 518
rect 1442 458 1446 461
rect 1442 448 1446 451
rect 1462 432 1465 458
rect 1478 451 1481 468
rect 1486 462 1489 478
rect 1510 472 1513 518
rect 1510 462 1513 468
rect 1518 462 1521 468
rect 1526 462 1529 478
rect 1478 448 1489 451
rect 1446 352 1449 378
rect 1438 342 1441 348
rect 1454 342 1457 398
rect 1486 392 1489 448
rect 1502 392 1505 448
rect 1542 422 1545 528
rect 1550 472 1553 508
rect 1598 472 1601 548
rect 1646 542 1649 548
rect 1618 538 1622 541
rect 1642 528 1646 531
rect 1614 512 1617 518
rect 1654 492 1657 498
rect 1626 488 1630 491
rect 1662 482 1665 558
rect 1734 552 1737 558
rect 1758 552 1761 618
rect 1830 602 1833 648
rect 1870 642 1873 648
rect 1878 632 1881 658
rect 1910 652 1913 658
rect 1862 592 1865 618
rect 1886 592 1889 648
rect 1894 572 1897 648
rect 1790 562 1793 568
rect 1822 562 1825 568
rect 1814 552 1817 558
rect 1878 552 1881 558
rect 1902 552 1905 598
rect 1910 562 1913 568
rect 1690 548 1694 551
rect 1722 548 1726 551
rect 1786 548 1790 551
rect 1670 502 1673 518
rect 1614 472 1617 478
rect 1634 468 1638 471
rect 1598 432 1601 468
rect 1646 462 1649 478
rect 1686 472 1689 538
rect 1658 468 1662 471
rect 1670 462 1673 468
rect 1694 462 1697 478
rect 1682 458 1686 461
rect 1606 452 1609 458
rect 1646 452 1649 458
rect 1520 403 1522 407
rect 1526 403 1529 407
rect 1533 403 1536 407
rect 1530 388 1534 391
rect 1470 332 1473 338
rect 1362 318 1369 321
rect 1326 282 1329 288
rect 1358 263 1361 278
rect 1210 138 1214 141
rect 1270 132 1273 147
rect 1294 72 1297 148
rect 1318 111 1321 198
rect 1330 168 1334 171
rect 1342 152 1345 258
rect 1366 152 1369 318
rect 1310 108 1321 111
rect 790 52 793 58
rect 1046 52 1049 59
rect 1198 62 1201 68
rect 1294 62 1297 68
rect 1310 62 1313 108
rect 1166 58 1169 59
rect 534 -19 538 -18
rect 526 -22 538 -19
rect 630 -19 634 -18
rect 638 -19 641 18
rect 630 -22 641 -19
rect 742 -19 745 18
rect 766 -18 769 18
rect 790 -18 793 8
rect 750 -19 754 -18
rect 742 -22 754 -19
rect 766 -22 770 -18
rect 790 -22 794 -18
rect 814 -19 817 18
rect 822 -19 826 -18
rect 814 -22 826 -19
rect 942 -19 946 -18
rect 950 -19 953 18
rect 942 -22 953 -19
rect 966 -19 970 -18
rect 974 -19 977 18
rect 966 -22 977 -19
rect 990 -19 994 -18
rect 998 -19 1001 18
rect 990 -22 1001 -19
rect 1030 -18 1033 8
rect 1030 -22 1034 -18
rect 1118 -19 1121 18
rect 1126 -19 1130 -18
rect 1118 -22 1130 -19
rect 1246 -19 1250 -18
rect 1254 -19 1257 18
rect 1246 -22 1257 -19
rect 1350 -19 1354 -18
rect 1358 -19 1361 118
rect 1374 61 1377 318
rect 1390 312 1393 318
rect 1422 292 1425 308
rect 1462 291 1465 318
rect 1454 288 1465 291
rect 1478 292 1481 358
rect 1494 342 1497 378
rect 1502 332 1505 348
rect 1510 292 1513 338
rect 1526 322 1529 328
rect 1542 312 1545 418
rect 1694 382 1697 418
rect 1666 378 1670 381
rect 1606 362 1609 368
rect 1702 352 1705 548
rect 1722 538 1726 541
rect 1710 452 1713 518
rect 1734 482 1737 548
rect 1718 472 1721 478
rect 1738 458 1742 461
rect 1710 362 1713 368
rect 1718 362 1721 458
rect 1750 442 1753 518
rect 1766 462 1769 468
rect 1774 462 1777 548
rect 1790 538 1798 541
rect 1790 492 1793 538
rect 1830 532 1833 548
rect 1862 542 1865 548
rect 1918 542 1921 638
rect 1926 622 1929 738
rect 1934 692 1937 738
rect 1934 652 1937 658
rect 1942 652 1945 678
rect 1950 662 1953 688
rect 1974 682 1977 748
rect 1982 732 1985 918
rect 2006 892 2009 918
rect 2014 892 2017 1058
rect 2102 1052 2105 1058
rect 2038 1012 2041 1048
rect 2042 1008 2049 1011
rect 2026 938 2030 941
rect 2024 903 2026 907
rect 2030 903 2033 907
rect 2037 903 2040 907
rect 1998 882 2001 888
rect 2046 882 2049 1008
rect 2054 1002 2057 1048
rect 2062 992 2065 1048
rect 2094 1042 2097 1048
rect 2054 972 2057 978
rect 2078 962 2081 1018
rect 2102 992 2105 1038
rect 2110 981 2113 1068
rect 2126 1062 2129 1068
rect 2142 1062 2145 1088
rect 2178 1078 2182 1081
rect 2158 1072 2161 1078
rect 2186 1068 2190 1071
rect 2150 1052 2153 1058
rect 2182 1052 2185 1058
rect 2174 1012 2177 1018
rect 2166 992 2169 998
rect 2102 978 2113 981
rect 2094 962 2097 968
rect 2062 932 2065 948
rect 1990 832 1993 858
rect 1990 752 1993 758
rect 1982 692 1985 708
rect 1990 662 1993 748
rect 1998 692 2001 868
rect 2006 842 2009 878
rect 2026 868 2030 871
rect 2046 852 2049 868
rect 2058 866 2062 869
rect 2018 848 2022 851
rect 2006 772 2009 838
rect 2014 762 2017 768
rect 2006 682 2009 738
rect 2030 732 2033 738
rect 2014 692 2017 718
rect 2046 711 2049 848
rect 2070 842 2073 958
rect 2102 952 2105 978
rect 2078 892 2081 928
rect 2094 892 2097 948
rect 2070 782 2073 818
rect 2086 792 2089 868
rect 2102 862 2105 948
rect 2110 932 2113 948
rect 2126 942 2129 948
rect 2110 922 2113 928
rect 2134 922 2137 958
rect 2174 952 2177 1008
rect 2154 948 2158 951
rect 2182 942 2185 1038
rect 2198 1032 2201 1138
rect 2210 1128 2214 1131
rect 2250 1128 2254 1131
rect 2230 1092 2233 1118
rect 2206 1072 2209 1078
rect 2214 1072 2217 1078
rect 2230 1068 2238 1071
rect 2250 1068 2254 1071
rect 2222 1062 2225 1068
rect 2210 1058 2214 1061
rect 2222 1052 2225 1058
rect 2206 992 2209 1048
rect 2230 1002 2233 1068
rect 2258 1058 2262 1061
rect 2246 1052 2249 1058
rect 2278 1052 2281 1188
rect 2302 1152 2305 1208
rect 2286 1142 2289 1148
rect 2310 1142 2313 1198
rect 2318 1192 2321 1218
rect 2334 1202 2337 1248
rect 2318 1141 2321 1178
rect 2326 1172 2329 1178
rect 2334 1152 2337 1178
rect 2318 1138 2326 1141
rect 2302 1102 2305 1138
rect 2310 1132 2313 1138
rect 2334 1102 2337 1148
rect 2342 1142 2345 1158
rect 2350 1152 2353 1158
rect 2358 1112 2361 1268
rect 2366 1262 2369 1278
rect 2370 1258 2374 1261
rect 2382 1252 2385 1278
rect 2390 1262 2393 1278
rect 2370 1248 2374 1251
rect 2390 1232 2393 1258
rect 2422 1252 2425 1278
rect 2482 1268 2486 1271
rect 2458 1258 2462 1261
rect 2366 1162 2369 1168
rect 2438 1162 2441 1198
rect 2446 1192 2449 1228
rect 2454 1222 2457 1258
rect 2466 1188 2470 1191
rect 2486 1172 2489 1258
rect 2494 1192 2497 1268
rect 2458 1158 2462 1161
rect 2386 1148 2390 1151
rect 2366 1102 2369 1118
rect 2350 1072 2353 1098
rect 2374 1082 2377 1138
rect 2398 1122 2401 1158
rect 2434 1148 2438 1151
rect 2406 1142 2409 1148
rect 2414 1132 2417 1138
rect 2454 1122 2457 1138
rect 2470 1132 2473 1168
rect 2482 1148 2486 1151
rect 2494 1142 2497 1148
rect 2510 1142 2513 1248
rect 2518 1222 2521 1268
rect 2534 1262 2537 1448
rect 2544 1403 2546 1407
rect 2550 1403 2553 1407
rect 2557 1403 2560 1407
rect 2574 1392 2577 1448
rect 2582 1381 2585 1558
rect 2590 1542 2593 1558
rect 2622 1552 2625 1608
rect 2654 1602 2657 1618
rect 2670 1562 2673 1648
rect 2694 1642 2697 1648
rect 2650 1558 2654 1561
rect 2634 1548 2638 1551
rect 2666 1548 2670 1551
rect 2590 1512 2593 1518
rect 2598 1472 2601 1548
rect 2606 1542 2609 1548
rect 2606 1482 2609 1538
rect 2622 1492 2625 1548
rect 2634 1538 2638 1541
rect 2654 1482 2657 1488
rect 2670 1482 2673 1508
rect 2602 1468 2606 1471
rect 2594 1388 2598 1391
rect 2574 1378 2585 1381
rect 2606 1382 2609 1468
rect 2630 1432 2633 1468
rect 2670 1462 2673 1478
rect 2642 1438 2646 1441
rect 2654 1432 2657 1458
rect 2686 1452 2689 1518
rect 2666 1448 2670 1451
rect 2674 1438 2678 1441
rect 2694 1441 2697 1538
rect 2710 1492 2713 1518
rect 2706 1458 2710 1461
rect 2694 1438 2702 1441
rect 2694 1422 2697 1438
rect 2646 1392 2649 1408
rect 2542 1332 2545 1378
rect 2566 1332 2569 1358
rect 2574 1292 2577 1378
rect 2586 1368 2590 1371
rect 2610 1368 2614 1371
rect 2638 1362 2641 1368
rect 2546 1268 2550 1271
rect 2558 1242 2561 1268
rect 2574 1242 2577 1248
rect 2518 1192 2521 1218
rect 2526 1142 2529 1238
rect 2582 1231 2585 1348
rect 2614 1342 2617 1348
rect 2598 1332 2601 1338
rect 2622 1292 2625 1358
rect 2662 1352 2665 1358
rect 2670 1352 2673 1398
rect 2702 1352 2705 1428
rect 2710 1352 2713 1458
rect 2718 1452 2721 1638
rect 2734 1631 2737 1718
rect 2742 1672 2745 1708
rect 2750 1662 2753 1718
rect 2758 1712 2761 1728
rect 2782 1682 2785 1718
rect 2790 1692 2793 1738
rect 2798 1732 2801 1868
rect 2830 1862 2833 1868
rect 2886 1862 2889 1868
rect 2902 1862 2905 1868
rect 2934 1862 2937 1868
rect 2818 1858 2822 1861
rect 2914 1858 2918 1861
rect 2954 1858 2958 1861
rect 2862 1852 2865 1858
rect 2826 1848 2838 1851
rect 2806 1792 2809 1848
rect 2814 1782 2817 1818
rect 2822 1752 2825 1758
rect 2814 1742 2817 1748
rect 2830 1741 2833 1808
rect 2846 1762 2849 1818
rect 2854 1802 2857 1848
rect 2902 1832 2905 1858
rect 2966 1852 2969 1978
rect 3166 1962 3169 1968
rect 3050 1958 3054 1961
rect 2974 1932 2977 1938
rect 2982 1892 2985 1948
rect 2998 1882 3001 1928
rect 2974 1872 2977 1878
rect 2998 1862 3001 1878
rect 3014 1872 3017 1948
rect 3030 1932 3033 1958
rect 3038 1932 3041 1938
rect 3038 1902 3041 1918
rect 3048 1903 3050 1907
rect 3054 1903 3057 1907
rect 3061 1903 3064 1907
rect 3078 1892 3081 1948
rect 3110 1932 3113 1948
rect 3150 1942 3153 1948
rect 3138 1938 3142 1941
rect 3174 1932 3177 1988
rect 3222 1962 3225 1968
rect 3254 1952 3257 1958
rect 3202 1948 3206 1951
rect 3218 1948 3222 1951
rect 3234 1948 3238 1951
rect 3182 1938 3190 1941
rect 3250 1938 3254 1941
rect 3162 1928 3166 1931
rect 3118 1892 3121 1908
rect 3026 1888 3030 1891
rect 3086 1882 3089 1888
rect 3042 1878 3046 1881
rect 3166 1872 3169 1878
rect 3070 1852 3073 1858
rect 2946 1838 2950 1841
rect 2910 1812 2913 1818
rect 2862 1752 2865 1758
rect 2826 1738 2833 1741
rect 2854 1722 2857 1748
rect 2878 1732 2881 1798
rect 2918 1792 2921 1838
rect 2942 1822 2945 1828
rect 3102 1792 3105 1858
rect 3170 1848 3174 1851
rect 3182 1832 3185 1938
rect 3198 1872 3201 1878
rect 3190 1862 3193 1868
rect 3206 1852 3209 1858
rect 3158 1802 3161 1818
rect 3190 1792 3193 1818
rect 3138 1788 3142 1791
rect 3130 1768 3134 1771
rect 2938 1758 2942 1761
rect 2942 1742 2945 1758
rect 3006 1752 3009 1768
rect 3162 1758 3166 1761
rect 2994 1748 2998 1751
rect 3038 1748 3046 1751
rect 3130 1748 3134 1751
rect 2930 1738 2934 1741
rect 2974 1741 2977 1748
rect 2910 1732 2913 1738
rect 2866 1728 2870 1731
rect 2902 1722 2905 1728
rect 2798 1682 2801 1718
rect 2766 1662 2769 1678
rect 2806 1672 2809 1698
rect 2834 1688 2838 1691
rect 2790 1662 2793 1668
rect 2838 1662 2841 1678
rect 2806 1658 2814 1661
rect 2806 1652 2809 1658
rect 2734 1628 2745 1631
rect 2726 1552 2729 1618
rect 2734 1572 2737 1618
rect 2730 1548 2734 1551
rect 2742 1542 2745 1628
rect 2750 1562 2753 1618
rect 2774 1582 2777 1618
rect 2814 1592 2817 1648
rect 2838 1592 2841 1628
rect 2846 1582 2849 1718
rect 2870 1692 2873 1708
rect 2854 1682 2857 1688
rect 2894 1672 2897 1698
rect 2918 1672 2921 1678
rect 2926 1672 2929 1678
rect 2934 1672 2937 1678
rect 2942 1672 2945 1718
rect 2950 1662 2953 1668
rect 2886 1652 2889 1658
rect 2958 1652 2961 1740
rect 2974 1738 2982 1741
rect 3002 1718 3006 1721
rect 2974 1702 2977 1718
rect 3014 1712 3017 1738
rect 3022 1722 3025 1728
rect 3030 1712 3033 1718
rect 2966 1692 2969 1698
rect 3006 1692 3009 1698
rect 2978 1678 2982 1681
rect 2978 1658 2982 1661
rect 2870 1632 2873 1648
rect 2990 1622 2993 1668
rect 3006 1652 3009 1668
rect 3014 1652 3017 1658
rect 3022 1632 3025 1658
rect 3038 1632 3041 1748
rect 3094 1742 3097 1748
rect 3066 1728 3070 1731
rect 3048 1703 3050 1707
rect 3054 1703 3057 1707
rect 3061 1703 3064 1707
rect 3094 1682 3097 1738
rect 3114 1728 3118 1731
rect 3026 1618 3030 1621
rect 2810 1548 2814 1551
rect 2734 1538 2742 1541
rect 2734 1531 2737 1538
rect 2730 1528 2737 1531
rect 2750 1522 2753 1528
rect 2742 1472 2745 1518
rect 2750 1472 2753 1478
rect 2634 1348 2638 1351
rect 2650 1328 2654 1331
rect 2674 1328 2678 1331
rect 2634 1288 2638 1291
rect 2614 1272 2617 1278
rect 2622 1272 2625 1278
rect 2614 1252 2617 1268
rect 2610 1238 2614 1241
rect 2574 1228 2585 1231
rect 2638 1232 2641 1268
rect 2646 1262 2649 1308
rect 2658 1258 2662 1261
rect 2544 1203 2546 1207
rect 2550 1203 2553 1207
rect 2557 1203 2560 1207
rect 2498 1128 2502 1131
rect 2518 1128 2526 1131
rect 2446 1118 2454 1121
rect 2438 1112 2441 1118
rect 2406 1082 2409 1088
rect 2266 1048 2270 1051
rect 2278 1032 2281 1048
rect 2206 962 2209 988
rect 2198 952 2201 958
rect 2190 942 2193 948
rect 2170 938 2174 941
rect 2118 912 2121 918
rect 2150 892 2153 938
rect 2214 932 2217 988
rect 2238 972 2241 998
rect 2250 968 2254 971
rect 2162 928 2166 931
rect 2222 922 2225 958
rect 2234 948 2238 951
rect 2230 932 2233 938
rect 2174 882 2177 888
rect 2138 878 2142 881
rect 2110 872 2113 878
rect 2194 868 2198 871
rect 2162 858 2166 861
rect 2106 848 2110 851
rect 2130 848 2134 851
rect 2102 792 2105 838
rect 2118 802 2121 818
rect 2134 792 2137 828
rect 2174 812 2177 868
rect 2206 862 2209 898
rect 2222 882 2225 918
rect 2230 882 2233 908
rect 2194 858 2198 861
rect 2182 852 2185 858
rect 2214 852 2217 868
rect 2230 862 2233 868
rect 2238 862 2241 948
rect 2246 942 2249 948
rect 2262 932 2265 1028
rect 2286 1012 2289 1068
rect 2322 1058 2326 1061
rect 2358 1061 2361 1078
rect 2414 1072 2417 1108
rect 2390 1062 2393 1068
rect 2354 1058 2361 1061
rect 2278 962 2281 978
rect 2294 972 2297 1058
rect 2314 1048 2318 1051
rect 2290 958 2294 961
rect 2278 952 2281 958
rect 2274 938 2278 941
rect 2246 861 2249 878
rect 2254 872 2257 918
rect 2262 882 2265 928
rect 2270 872 2273 938
rect 2294 912 2297 948
rect 2310 942 2313 1008
rect 2318 952 2321 968
rect 2302 932 2305 938
rect 2326 922 2329 1058
rect 2342 1052 2345 1058
rect 2350 1002 2353 1058
rect 2382 1052 2385 1058
rect 2406 1052 2409 1068
rect 2422 1052 2425 1058
rect 2446 1052 2449 1118
rect 2486 1072 2489 1098
rect 2498 1078 2502 1081
rect 2510 1072 2513 1128
rect 2518 1092 2521 1128
rect 2550 1122 2553 1148
rect 2574 1141 2577 1228
rect 2626 1158 2630 1161
rect 2582 1152 2585 1158
rect 2646 1152 2649 1258
rect 2606 1142 2609 1148
rect 2574 1138 2585 1141
rect 2558 1092 2561 1138
rect 2570 1128 2577 1131
rect 2566 1081 2569 1118
rect 2558 1078 2569 1081
rect 2534 1072 2537 1078
rect 2482 1058 2486 1061
rect 2558 1052 2561 1078
rect 2510 1032 2513 1048
rect 2334 942 2337 948
rect 2278 882 2281 898
rect 2246 858 2254 861
rect 2278 861 2281 868
rect 2258 858 2281 861
rect 2230 842 2233 848
rect 2070 762 2073 778
rect 2106 748 2110 751
rect 2098 738 2102 741
rect 2054 722 2057 738
rect 2046 708 2057 711
rect 2024 703 2026 707
rect 2030 703 2033 707
rect 2037 703 2040 707
rect 2034 688 2046 691
rect 2010 678 2014 681
rect 2010 658 2014 661
rect 1950 652 1953 658
rect 1950 632 1953 638
rect 1958 602 1961 638
rect 1974 592 1977 598
rect 1982 561 1985 618
rect 1982 558 1990 561
rect 2002 558 2009 561
rect 1994 548 1998 551
rect 1846 532 1849 538
rect 1854 532 1857 538
rect 1938 528 1942 531
rect 1782 482 1785 488
rect 1838 481 1841 518
rect 1854 492 1857 508
rect 1910 492 1913 528
rect 1918 482 1921 508
rect 1838 478 1846 481
rect 1826 468 1830 471
rect 1726 372 1729 418
rect 1758 392 1761 418
rect 1790 392 1793 468
rect 1810 458 1814 461
rect 1866 458 1870 461
rect 1822 451 1825 458
rect 1818 448 1825 451
rect 1798 422 1801 448
rect 1822 392 1825 398
rect 1846 392 1849 458
rect 1870 392 1873 428
rect 1770 368 1774 371
rect 1806 362 1809 368
rect 1746 358 1750 361
rect 1866 358 1870 361
rect 1566 342 1569 348
rect 1554 338 1558 341
rect 1582 332 1585 348
rect 1590 342 1593 348
rect 1646 342 1649 348
rect 1702 342 1705 348
rect 1638 332 1641 338
rect 1662 332 1666 335
rect 1574 322 1577 328
rect 1694 322 1697 338
rect 1718 331 1721 358
rect 1790 352 1793 358
rect 1730 348 1734 351
rect 1850 348 1854 351
rect 1730 338 1734 341
rect 1802 338 1806 341
rect 1718 328 1729 331
rect 1646 298 1654 301
rect 1454 278 1457 288
rect 1478 272 1481 288
rect 1494 272 1497 278
rect 1550 272 1553 298
rect 1582 272 1585 278
rect 1390 262 1393 268
rect 1430 152 1433 218
rect 1454 192 1457 218
rect 1520 203 1522 207
rect 1526 203 1529 207
rect 1533 203 1536 207
rect 1526 151 1529 188
rect 1558 142 1561 148
rect 1598 142 1601 298
rect 1610 258 1614 261
rect 1646 192 1649 298
rect 1662 292 1665 318
rect 1690 288 1694 291
rect 1670 272 1673 278
rect 1718 272 1721 278
rect 1726 262 1729 328
rect 1734 292 1737 308
rect 1750 302 1753 318
rect 1758 312 1761 328
rect 1762 288 1766 291
rect 1742 282 1745 288
rect 1782 275 1786 278
rect 1746 268 1750 271
rect 1758 192 1761 258
rect 1782 252 1785 258
rect 1394 118 1398 121
rect 1382 71 1385 118
rect 1382 68 1393 71
rect 1374 58 1382 61
rect 1350 -22 1361 -19
rect 1366 -19 1370 -18
rect 1374 -19 1377 18
rect 1366 -22 1377 -19
rect 1382 -19 1386 -18
rect 1390 -19 1393 68
rect 1406 62 1409 118
rect 1454 82 1457 128
rect 1590 112 1593 118
rect 1462 62 1465 108
rect 1526 62 1529 88
rect 1566 62 1569 108
rect 1630 72 1633 138
rect 1646 82 1649 188
rect 1662 142 1665 148
rect 1678 142 1681 148
rect 1694 142 1697 147
rect 1710 82 1713 138
rect 1774 132 1777 138
rect 1614 63 1617 68
rect 1718 62 1721 88
rect 1790 62 1793 158
rect 1814 152 1817 348
rect 1822 342 1825 348
rect 1878 342 1881 468
rect 1886 352 1889 468
rect 1894 462 1897 478
rect 1942 472 1945 518
rect 1966 492 1969 538
rect 1974 532 1977 548
rect 1934 462 1937 468
rect 1842 338 1846 341
rect 1882 338 1886 341
rect 1822 292 1825 338
rect 1822 278 1830 281
rect 1822 272 1825 278
rect 1846 272 1849 328
rect 1870 312 1873 328
rect 1878 292 1881 328
rect 1834 268 1838 271
rect 1826 258 1830 261
rect 1798 122 1801 148
rect 1814 81 1817 148
rect 1814 78 1825 81
rect 1814 62 1817 68
rect 1822 62 1825 78
rect 1838 81 1841 268
rect 1846 258 1854 261
rect 1846 162 1849 258
rect 1862 251 1865 258
rect 1854 248 1865 251
rect 1854 222 1857 248
rect 1854 192 1857 218
rect 1886 212 1889 268
rect 1894 262 1897 448
rect 1934 362 1937 368
rect 1910 332 1913 358
rect 1942 352 1945 468
rect 1966 462 1969 488
rect 1990 472 1993 528
rect 2006 522 2009 558
rect 2014 552 2017 628
rect 2054 592 2057 708
rect 2062 652 2065 718
rect 2078 662 2081 728
rect 2118 712 2121 758
rect 2138 748 2142 751
rect 2130 738 2134 741
rect 2118 692 2121 698
rect 2134 692 2137 708
rect 2086 672 2089 678
rect 2090 668 2094 671
rect 2074 658 2078 661
rect 2106 658 2110 661
rect 2094 632 2097 658
rect 2110 648 2118 651
rect 1998 482 2001 488
rect 2014 462 2017 548
rect 2022 542 2025 558
rect 2062 552 2065 618
rect 2110 592 2113 648
rect 2126 612 2129 678
rect 2142 662 2145 668
rect 2150 662 2153 738
rect 2158 732 2161 778
rect 2174 752 2177 808
rect 2198 792 2201 838
rect 2190 752 2193 768
rect 2174 742 2177 748
rect 2182 742 2185 748
rect 2214 742 2217 758
rect 2222 752 2225 758
rect 2238 742 2241 848
rect 2286 842 2289 848
rect 2278 832 2281 838
rect 2246 792 2249 808
rect 2254 752 2257 758
rect 2262 752 2265 768
rect 2282 748 2286 751
rect 2294 742 2297 878
rect 2318 872 2321 918
rect 2302 862 2305 868
rect 2310 862 2313 868
rect 2342 861 2345 938
rect 2350 902 2353 948
rect 2358 942 2361 968
rect 2374 962 2377 968
rect 2378 948 2382 951
rect 2374 892 2377 948
rect 2386 938 2390 941
rect 2398 872 2401 988
rect 2422 962 2425 1018
rect 2454 1012 2457 1018
rect 2406 952 2409 958
rect 2406 932 2409 938
rect 2354 868 2358 871
rect 2386 868 2390 871
rect 2374 862 2377 868
rect 2342 858 2353 861
rect 2342 842 2345 848
rect 2310 792 2313 838
rect 2310 772 2313 788
rect 2318 762 2321 798
rect 2326 752 2329 818
rect 2350 792 2353 858
rect 2358 852 2361 858
rect 2370 848 2374 851
rect 2234 738 2238 741
rect 2158 682 2161 718
rect 2166 661 2169 728
rect 2174 722 2177 738
rect 2190 732 2193 738
rect 2242 728 2246 731
rect 2214 692 2217 728
rect 2254 692 2257 738
rect 2286 732 2289 738
rect 2302 682 2305 688
rect 2178 668 2182 671
rect 2194 668 2198 671
rect 2214 662 2217 668
rect 2166 658 2174 661
rect 2150 622 2153 658
rect 2178 648 2182 651
rect 2126 592 2129 598
rect 2074 558 2078 561
rect 2054 532 2057 538
rect 2046 522 2049 528
rect 2024 503 2026 507
rect 2030 503 2033 507
rect 2037 503 2040 507
rect 2062 492 2065 548
rect 2074 528 2078 531
rect 2078 492 2081 508
rect 2022 472 2025 478
rect 1950 452 1953 458
rect 1974 452 1977 458
rect 2002 448 2006 451
rect 1922 348 1926 351
rect 1942 342 1945 348
rect 1922 338 1926 341
rect 1954 338 1958 341
rect 1914 328 1918 331
rect 1910 292 1913 318
rect 1950 292 1953 308
rect 1966 292 1969 358
rect 1974 352 1977 358
rect 1982 342 1985 378
rect 1998 362 2001 368
rect 2006 352 2009 428
rect 2014 412 2017 458
rect 2030 392 2033 488
rect 2062 482 2065 488
rect 2070 472 2073 488
rect 2046 452 2049 468
rect 1998 342 2001 348
rect 2014 342 2017 358
rect 2046 352 2049 448
rect 2070 372 2073 448
rect 2078 392 2081 398
rect 2058 358 2062 361
rect 2086 351 2089 578
rect 2134 572 2137 578
rect 2118 552 2121 558
rect 2098 538 2102 541
rect 2094 482 2097 498
rect 2110 492 2113 538
rect 2114 478 2118 481
rect 2098 468 2102 471
rect 2122 468 2126 471
rect 2122 458 2126 461
rect 2094 392 2097 408
rect 2118 362 2121 418
rect 2134 392 2137 548
rect 2150 441 2153 558
rect 2158 552 2161 638
rect 2158 492 2161 548
rect 2174 532 2177 618
rect 2190 552 2193 568
rect 2198 552 2201 658
rect 2230 652 2233 658
rect 2238 622 2241 668
rect 2158 462 2161 468
rect 2166 451 2169 488
rect 2174 482 2177 518
rect 2190 502 2193 548
rect 2182 482 2185 488
rect 2162 448 2169 451
rect 2174 452 2177 468
rect 2198 452 2201 548
rect 2206 492 2209 548
rect 2214 512 2217 538
rect 2230 532 2233 538
rect 2222 522 2225 528
rect 2238 521 2241 558
rect 2230 518 2241 521
rect 2230 492 2233 518
rect 2222 472 2225 488
rect 2214 452 2217 468
rect 2230 462 2233 468
rect 2150 438 2161 441
rect 2158 392 2161 438
rect 2190 392 2193 428
rect 2170 368 2174 371
rect 2122 358 2134 361
rect 2154 358 2158 361
rect 2086 348 2094 351
rect 2014 292 2017 338
rect 2046 312 2049 348
rect 2078 342 2081 348
rect 2024 303 2026 307
rect 2030 303 2033 307
rect 2037 303 2040 307
rect 2054 302 2057 338
rect 2086 302 2089 338
rect 2002 288 2006 291
rect 2054 282 2057 298
rect 1910 272 1913 278
rect 1958 272 1961 278
rect 1990 272 1993 278
rect 2070 272 2073 278
rect 1922 268 1926 271
rect 2026 268 2030 271
rect 1942 262 1945 268
rect 1858 158 1862 161
rect 1910 151 1913 168
rect 1878 142 1881 148
rect 1894 132 1897 138
rect 1918 131 1921 188
rect 1910 128 1921 131
rect 1834 78 1841 81
rect 1830 72 1833 78
rect 1850 58 1854 61
rect 1798 52 1801 58
rect 1862 51 1865 118
rect 1878 92 1881 118
rect 1910 92 1913 128
rect 1926 92 1929 208
rect 1934 202 1937 258
rect 1942 252 1945 258
rect 1990 252 1993 268
rect 2094 262 2097 348
rect 2102 292 2105 308
rect 2110 292 2113 328
rect 2134 322 2137 348
rect 2146 338 2153 341
rect 2126 292 2129 318
rect 2150 292 2153 338
rect 2158 312 2161 348
rect 2182 332 2185 348
rect 2190 342 2193 378
rect 2214 352 2217 358
rect 2238 352 2241 488
rect 2246 362 2249 668
rect 2270 662 2273 668
rect 2278 662 2281 668
rect 2294 652 2297 668
rect 2254 592 2257 608
rect 2294 592 2297 628
rect 2262 552 2265 568
rect 2282 558 2286 561
rect 2270 552 2273 558
rect 2310 542 2313 748
rect 2330 738 2334 741
rect 2338 738 2345 741
rect 2354 738 2358 741
rect 2326 662 2329 728
rect 2342 682 2345 738
rect 2366 692 2369 738
rect 2374 692 2377 838
rect 2382 802 2385 848
rect 2382 782 2385 788
rect 2406 752 2409 918
rect 2414 842 2417 948
rect 2422 942 2425 948
rect 2454 942 2457 958
rect 2430 932 2433 938
rect 2450 928 2454 931
rect 2430 881 2433 928
rect 2438 922 2441 928
rect 2462 922 2465 948
rect 2478 942 2481 1028
rect 2518 972 2521 1048
rect 2550 1042 2553 1048
rect 2558 1021 2561 1048
rect 2566 1032 2569 1068
rect 2558 1018 2569 1021
rect 2544 1003 2546 1007
rect 2550 1003 2553 1007
rect 2557 1003 2560 1007
rect 2514 968 2518 971
rect 2522 958 2526 961
rect 2566 952 2569 1018
rect 2574 992 2577 1128
rect 2582 1092 2585 1138
rect 2622 1132 2625 1138
rect 2646 1132 2649 1138
rect 2654 1132 2657 1138
rect 2602 1128 2606 1131
rect 2634 1118 2638 1121
rect 2614 1102 2617 1118
rect 2662 1112 2665 1118
rect 2670 1101 2673 1288
rect 2678 1282 2681 1318
rect 2686 1292 2689 1318
rect 2682 1278 2686 1281
rect 2678 1172 2681 1258
rect 2686 1242 2689 1268
rect 2694 1212 2697 1338
rect 2702 1312 2705 1348
rect 2718 1342 2721 1448
rect 2726 1442 2729 1448
rect 2746 1438 2750 1441
rect 2734 1382 2737 1418
rect 2758 1371 2761 1518
rect 2766 1512 2769 1548
rect 2766 1472 2769 1498
rect 2774 1462 2777 1508
rect 2774 1432 2777 1458
rect 2782 1442 2785 1448
rect 2774 1392 2777 1418
rect 2790 1412 2793 1538
rect 2822 1522 2825 1568
rect 2830 1562 2833 1578
rect 2854 1572 2857 1618
rect 2902 1602 2905 1618
rect 3046 1612 3049 1658
rect 3022 1592 3025 1608
rect 3046 1592 3049 1598
rect 2842 1568 2846 1571
rect 2866 1558 2870 1561
rect 2858 1548 2862 1551
rect 2890 1548 2894 1551
rect 2914 1538 2918 1541
rect 2874 1528 2878 1531
rect 2910 1522 2913 1528
rect 2882 1488 2886 1491
rect 2842 1478 2846 1481
rect 2806 1472 2809 1478
rect 2862 1472 2865 1478
rect 2802 1458 2806 1461
rect 2810 1448 2814 1451
rect 2822 1441 2825 1458
rect 2814 1438 2825 1441
rect 2814 1422 2817 1438
rect 2830 1432 2833 1438
rect 2758 1368 2766 1371
rect 2766 1362 2769 1368
rect 2790 1362 2793 1378
rect 2738 1358 2742 1361
rect 2782 1352 2785 1358
rect 2742 1348 2750 1351
rect 2710 1292 2713 1338
rect 2726 1322 2729 1328
rect 2718 1282 2721 1318
rect 2726 1262 2729 1268
rect 2734 1262 2737 1318
rect 2742 1272 2745 1348
rect 2750 1342 2753 1348
rect 2774 1332 2777 1348
rect 2798 1312 2801 1418
rect 2806 1392 2809 1408
rect 2822 1382 2825 1418
rect 2838 1362 2841 1448
rect 2846 1432 2849 1438
rect 2862 1372 2865 1458
rect 2814 1322 2817 1338
rect 2822 1332 2825 1338
rect 2846 1332 2849 1358
rect 2862 1352 2865 1368
rect 2854 1332 2857 1338
rect 2762 1288 2766 1291
rect 2742 1262 2745 1268
rect 2706 1258 2710 1261
rect 2750 1252 2753 1268
rect 2706 1248 2710 1251
rect 2766 1222 2769 1278
rect 2774 1272 2777 1278
rect 2786 1268 2790 1271
rect 2798 1262 2801 1288
rect 2810 1268 2817 1271
rect 2782 1252 2785 1258
rect 2806 1222 2809 1258
rect 2814 1252 2817 1268
rect 2678 1152 2681 1168
rect 2702 1142 2705 1218
rect 2726 1162 2729 1198
rect 2662 1098 2673 1101
rect 2694 1132 2697 1138
rect 2662 1092 2665 1098
rect 2694 1092 2697 1128
rect 2702 1092 2705 1108
rect 2670 1082 2673 1088
rect 2710 1082 2713 1148
rect 2750 1142 2753 1158
rect 2774 1132 2777 1148
rect 2782 1142 2785 1168
rect 2790 1152 2793 1198
rect 2822 1172 2825 1328
rect 2830 1311 2833 1318
rect 2830 1308 2838 1311
rect 2862 1282 2865 1308
rect 2870 1302 2873 1458
rect 2878 1452 2881 1458
rect 2894 1452 2897 1468
rect 2902 1462 2905 1468
rect 2910 1462 2913 1518
rect 2926 1462 2929 1568
rect 2946 1558 2950 1561
rect 2942 1532 2945 1558
rect 2950 1548 2958 1551
rect 2950 1482 2953 1548
rect 2966 1492 2969 1548
rect 2974 1542 2977 1548
rect 2998 1532 3001 1538
rect 2990 1492 2993 1528
rect 2938 1478 2942 1481
rect 2890 1388 2894 1391
rect 2926 1382 2929 1458
rect 2950 1442 2953 1468
rect 2946 1348 2950 1351
rect 2886 1312 2889 1338
rect 2910 1332 2913 1348
rect 2874 1298 2881 1301
rect 2870 1272 2873 1288
rect 2842 1258 2846 1261
rect 2854 1251 2857 1258
rect 2834 1248 2857 1251
rect 2862 1242 2865 1248
rect 2830 1192 2833 1238
rect 2814 1152 2817 1168
rect 2730 1128 2758 1131
rect 2738 1118 2742 1121
rect 2782 1102 2785 1118
rect 2798 1092 2801 1108
rect 2838 1092 2841 1168
rect 2846 1152 2849 1238
rect 2878 1171 2881 1298
rect 2886 1292 2889 1308
rect 2918 1302 2921 1338
rect 2930 1328 2934 1331
rect 2942 1292 2945 1348
rect 2958 1341 2961 1458
rect 2954 1338 2961 1341
rect 2950 1332 2953 1338
rect 2966 1332 2969 1478
rect 2982 1472 2985 1488
rect 2990 1462 2993 1468
rect 3006 1452 3009 1548
rect 3030 1532 3033 1558
rect 3038 1548 3046 1551
rect 3022 1461 3025 1518
rect 3038 1492 3041 1548
rect 3058 1538 3062 1541
rect 3048 1503 3050 1507
rect 3054 1503 3057 1507
rect 3061 1503 3064 1507
rect 3054 1472 3057 1488
rect 3070 1482 3073 1678
rect 3082 1668 3086 1671
rect 3098 1658 3102 1661
rect 3106 1658 3110 1661
rect 3098 1648 3102 1651
rect 3110 1642 3113 1648
rect 3094 1592 3097 1628
rect 3078 1532 3081 1558
rect 3086 1522 3089 1578
rect 3062 1472 3065 1478
rect 3022 1458 3030 1461
rect 3018 1448 3025 1451
rect 2974 1442 2977 1448
rect 3006 1441 3009 1448
rect 3006 1438 3017 1441
rect 2990 1432 2993 1438
rect 3014 1392 3017 1438
rect 3002 1348 3006 1351
rect 2974 1342 2977 1348
rect 2950 1272 2953 1288
rect 2958 1272 2961 1318
rect 2974 1302 2977 1338
rect 3006 1292 3009 1298
rect 3022 1292 3025 1448
rect 3046 1352 3049 1468
rect 3078 1442 3081 1468
rect 3086 1462 3089 1518
rect 3094 1482 3097 1548
rect 3102 1542 3105 1558
rect 3118 1552 3121 1668
rect 3126 1651 3129 1728
rect 3142 1702 3145 1758
rect 3206 1752 3209 1848
rect 3222 1842 3225 1918
rect 3230 1822 3233 1858
rect 3238 1852 3241 1878
rect 3254 1832 3257 1858
rect 3222 1761 3225 1818
rect 3222 1758 3230 1761
rect 3194 1748 3198 1751
rect 3154 1738 3158 1741
rect 3194 1738 3198 1741
rect 3234 1738 3238 1741
rect 3182 1732 3185 1738
rect 3206 1732 3209 1738
rect 3138 1678 3142 1681
rect 3166 1662 3169 1668
rect 3154 1658 3158 1661
rect 3126 1648 3134 1651
rect 3122 1548 3126 1551
rect 3142 1551 3145 1648
rect 3150 1582 3153 1618
rect 3150 1562 3153 1568
rect 3158 1552 3161 1558
rect 3166 1552 3169 1658
rect 3182 1652 3185 1698
rect 3190 1672 3193 1678
rect 3198 1662 3201 1668
rect 3174 1572 3177 1618
rect 3190 1562 3193 1568
rect 3174 1552 3177 1558
rect 3142 1548 3153 1551
rect 3134 1542 3137 1548
rect 3110 1522 3113 1538
rect 3142 1532 3145 1538
rect 3142 1492 3145 1528
rect 3150 1492 3153 1548
rect 3166 1532 3169 1538
rect 3206 1492 3209 1728
rect 3222 1661 3225 1708
rect 3230 1702 3233 1718
rect 3246 1672 3249 1748
rect 3254 1682 3257 1768
rect 3262 1762 3265 2028
rect 3302 2022 3305 2068
rect 3334 2062 3337 2068
rect 3326 2022 3329 2058
rect 3334 2052 3337 2058
rect 3342 2042 3345 2228
rect 3350 2152 3353 2178
rect 3358 2142 3361 2148
rect 3366 2122 3369 2268
rect 3374 2152 3377 2248
rect 3382 2232 3385 2258
rect 3382 2172 3385 2228
rect 3390 2212 3393 2268
rect 3398 2252 3401 2278
rect 3446 2262 3449 2278
rect 3422 2242 3425 2258
rect 3434 2248 3438 2251
rect 3446 2192 3449 2238
rect 3462 2202 3465 2268
rect 3474 2258 3478 2261
rect 3486 2182 3489 2318
rect 3534 2312 3537 2338
rect 3494 2270 3497 2278
rect 3510 2272 3513 2288
rect 3530 2268 3534 2271
rect 3502 2261 3505 2268
rect 3502 2258 3513 2261
rect 3454 2172 3457 2178
rect 3382 2152 3385 2158
rect 3438 2152 3441 2158
rect 3458 2148 3462 2151
rect 3398 2142 3401 2148
rect 3422 2142 3425 2148
rect 3410 2138 3414 2141
rect 3366 2082 3369 2118
rect 3374 2112 3377 2128
rect 3430 2122 3433 2138
rect 3398 2092 3401 2098
rect 3438 2082 3441 2088
rect 3486 2082 3489 2158
rect 3494 2142 3497 2148
rect 3502 2132 3505 2168
rect 3510 2162 3513 2258
rect 3534 2252 3537 2258
rect 3518 2172 3521 2178
rect 3514 2158 3518 2161
rect 3494 2092 3497 2108
rect 3502 2092 3505 2118
rect 3494 2082 3497 2088
rect 3374 2062 3377 2068
rect 3390 2062 3393 2068
rect 3510 2062 3513 2128
rect 3518 2122 3521 2148
rect 3526 2092 3529 2168
rect 3542 2161 3545 2348
rect 3586 2328 3590 2331
rect 3550 2282 3553 2288
rect 3590 2282 3593 2288
rect 3578 2278 3582 2281
rect 3598 2272 3601 2358
rect 3686 2352 3689 2358
rect 3750 2352 3753 2358
rect 3618 2348 3622 2351
rect 3650 2348 3654 2351
rect 3698 2348 3702 2351
rect 3654 2342 3657 2348
rect 3766 2342 3769 2348
rect 3610 2338 3614 2341
rect 3730 2338 3734 2341
rect 3622 2292 3625 2318
rect 3638 2302 3641 2318
rect 3646 2272 3649 2278
rect 3602 2268 3606 2271
rect 3550 2262 3553 2268
rect 3662 2262 3665 2338
rect 3686 2332 3689 2338
rect 3694 2322 3697 2328
rect 3686 2292 3689 2308
rect 3702 2282 3705 2298
rect 3674 2278 3678 2281
rect 3726 2272 3729 2278
rect 3742 2272 3745 2328
rect 3774 2312 3777 2358
rect 3806 2352 3809 2358
rect 3822 2352 3825 2398
rect 3830 2352 3833 2358
rect 3818 2348 3822 2351
rect 3786 2338 3790 2341
rect 3786 2328 3790 2331
rect 3750 2272 3753 2278
rect 3758 2272 3761 2278
rect 3690 2258 3694 2261
rect 3738 2258 3742 2261
rect 3782 2261 3785 2318
rect 3798 2302 3801 2328
rect 3814 2282 3817 2338
rect 3822 2292 3825 2338
rect 3838 2311 3841 2428
rect 3910 2402 3913 2448
rect 3918 2431 3921 2458
rect 3958 2452 3961 2458
rect 3966 2452 3969 2488
rect 3974 2482 3977 2518
rect 3990 2512 3993 2548
rect 3994 2508 4001 2511
rect 3986 2468 3990 2471
rect 3926 2442 3929 2448
rect 3974 2442 3977 2458
rect 3998 2452 4001 2508
rect 4006 2462 4009 2558
rect 4038 2542 4041 2578
rect 4046 2532 4049 2568
rect 4062 2562 4065 2618
rect 4062 2542 4065 2558
rect 4078 2552 4081 2558
rect 4086 2542 4089 2658
rect 4102 2572 4105 2618
rect 4118 2592 4121 2678
rect 4126 2662 4129 2668
rect 4142 2652 4145 2698
rect 4210 2678 4214 2681
rect 4230 2672 4233 2698
rect 4246 2672 4249 2678
rect 4254 2672 4257 2718
rect 4262 2682 4265 2748
rect 4302 2742 4305 2748
rect 4310 2742 4313 2758
rect 4378 2748 4382 2751
rect 4282 2738 4286 2741
rect 4346 2738 4350 2741
rect 4278 2732 4281 2738
rect 4286 2732 4289 2738
rect 4306 2728 4310 2731
rect 4270 2682 4273 2718
rect 4274 2668 4278 2671
rect 4214 2662 4217 2668
rect 4286 2662 4289 2678
rect 4310 2672 4313 2678
rect 4318 2662 4321 2718
rect 4358 2712 4361 2718
rect 4390 2692 4393 2748
rect 4358 2682 4361 2688
rect 4334 2672 4337 2678
rect 4202 2658 4206 2661
rect 4322 2658 4326 2661
rect 4134 2572 4137 2618
rect 4142 2561 4145 2648
rect 4158 2642 4161 2658
rect 4210 2648 4214 2651
rect 4138 2558 4145 2561
rect 4134 2552 4137 2558
rect 4142 2542 4145 2548
rect 4086 2532 4089 2538
rect 4006 2442 4009 2458
rect 4014 2442 4017 2518
rect 4030 2452 4033 2478
rect 4050 2468 4054 2471
rect 4062 2462 4065 2518
rect 4080 2503 4082 2507
rect 4086 2503 4089 2507
rect 4093 2503 4096 2507
rect 4090 2488 4094 2491
rect 4110 2482 4113 2488
rect 4134 2482 4137 2498
rect 4078 2472 4081 2478
rect 4138 2468 4142 2471
rect 4118 2462 4121 2468
rect 4150 2462 4153 2598
rect 4158 2562 4161 2568
rect 4166 2552 4169 2648
rect 4186 2638 4190 2641
rect 4174 2632 4177 2638
rect 4182 2541 4185 2618
rect 4278 2562 4281 2658
rect 4302 2652 4305 2658
rect 4318 2642 4321 2648
rect 4286 2582 4289 2618
rect 4250 2558 4254 2561
rect 4210 2548 4214 2551
rect 4230 2542 4233 2558
rect 4278 2552 4281 2558
rect 4174 2538 4185 2541
rect 4194 2538 4198 2541
rect 4174 2502 4177 2538
rect 4194 2528 4198 2531
rect 4182 2522 4185 2528
rect 4166 2482 4169 2488
rect 4174 2472 4177 2478
rect 4074 2458 4078 2461
rect 4154 2458 4158 2461
rect 3986 2438 3990 2441
rect 3918 2428 3929 2431
rect 3918 2392 3921 2418
rect 3926 2392 3929 2428
rect 4006 2412 4009 2418
rect 4046 2412 4049 2418
rect 3926 2382 3929 2388
rect 3870 2362 3873 2378
rect 3878 2372 3881 2378
rect 3830 2308 3841 2311
rect 3914 2358 3918 2361
rect 3962 2358 3966 2361
rect 3846 2352 3849 2358
rect 3830 2282 3833 2308
rect 3838 2282 3841 2298
rect 3802 2278 3806 2281
rect 3790 2272 3793 2278
rect 3778 2258 3785 2261
rect 3798 2262 3801 2278
rect 3814 2262 3817 2268
rect 3846 2262 3849 2348
rect 3854 2342 3857 2348
rect 3862 2342 3865 2358
rect 3862 2292 3865 2328
rect 3870 2312 3873 2348
rect 3894 2282 3897 2338
rect 3910 2302 3913 2358
rect 3974 2352 3977 2358
rect 4018 2348 4022 2351
rect 3918 2332 3921 2348
rect 3942 2342 3945 2348
rect 3998 2342 4001 2348
rect 4030 2342 4033 2378
rect 4046 2352 4049 2398
rect 4062 2362 4065 2378
rect 4118 2372 4121 2418
rect 4146 2358 4150 2361
rect 4046 2342 4049 2348
rect 3970 2338 3974 2341
rect 3910 2282 3913 2298
rect 3998 2282 4001 2338
rect 4006 2332 4009 2338
rect 4014 2332 4017 2338
rect 4126 2332 4129 2348
rect 4142 2342 4145 2358
rect 4150 2342 4153 2348
rect 4174 2342 4177 2468
rect 4190 2462 4193 2518
rect 4198 2472 4201 2478
rect 4222 2471 4225 2518
rect 4222 2468 4230 2471
rect 4214 2462 4217 2468
rect 4238 2462 4241 2548
rect 4270 2542 4273 2548
rect 4254 2532 4257 2538
rect 4302 2532 4305 2568
rect 4326 2562 4329 2568
rect 4334 2562 4337 2668
rect 4350 2662 4353 2678
rect 4378 2668 4382 2671
rect 4350 2652 4353 2658
rect 4374 2652 4377 2658
rect 4398 2652 4401 2738
rect 4406 2682 4409 2728
rect 4406 2672 4409 2678
rect 4422 2672 4425 2858
rect 4454 2762 4457 2859
rect 4470 2852 4473 2878
rect 4582 2872 4585 2878
rect 4462 2752 4465 2778
rect 4478 2742 4481 2858
rect 4542 2852 4545 2868
rect 4558 2862 4561 2868
rect 4582 2852 4585 2858
rect 4562 2838 4566 2841
rect 4478 2682 4481 2738
rect 4454 2652 4457 2658
rect 4394 2648 4398 2651
rect 4342 2572 4345 2618
rect 4310 2542 4313 2558
rect 4322 2538 4326 2541
rect 4334 2532 4337 2538
rect 4342 2522 4345 2558
rect 4406 2552 4409 2558
rect 4438 2542 4441 2568
rect 4534 2562 4537 2747
rect 4558 2562 4561 2658
rect 4514 2558 4518 2561
rect 4470 2552 4473 2558
rect 4470 2542 4473 2548
rect 4486 2542 4489 2548
rect 4522 2538 4526 2541
rect 4350 2532 4353 2538
rect 4382 2532 4385 2538
rect 4414 2532 4417 2538
rect 4402 2528 4406 2531
rect 4450 2528 4454 2531
rect 4254 2482 4257 2508
rect 4278 2492 4281 2498
rect 4282 2478 4286 2481
rect 4326 2472 4329 2498
rect 4342 2491 4345 2518
rect 4334 2488 4345 2491
rect 4258 2468 4262 2471
rect 4334 2462 4337 2488
rect 4358 2481 4361 2518
rect 4350 2478 4361 2481
rect 4366 2482 4369 2518
rect 4342 2472 4345 2478
rect 4350 2462 4353 2478
rect 4226 2458 4230 2461
rect 4250 2458 4254 2461
rect 4198 2451 4201 2458
rect 4190 2448 4201 2451
rect 4190 2442 4193 2448
rect 4286 2442 4289 2458
rect 4346 2448 4350 2451
rect 4358 2422 4361 2468
rect 4366 2452 4369 2478
rect 4382 2472 4385 2528
rect 4390 2502 4393 2528
rect 4390 2472 4393 2498
rect 4430 2472 4433 2478
rect 4438 2472 4441 2528
rect 4446 2482 4449 2518
rect 4462 2512 4465 2528
rect 4494 2512 4497 2538
rect 4518 2482 4521 2508
rect 4430 2462 4433 2468
rect 4446 2462 4449 2468
rect 4486 2462 4489 2478
rect 4406 2452 4409 2458
rect 4414 2452 4417 2458
rect 4454 2452 4457 2458
rect 4526 2452 4529 2518
rect 4534 2481 4537 2558
rect 4546 2548 4550 2551
rect 4558 2522 4561 2558
rect 4558 2482 4561 2518
rect 4534 2478 4542 2481
rect 4574 2472 4577 2538
rect 4590 2492 4593 3158
rect 4598 2862 4601 2868
rect 4598 2792 4601 2848
rect 4598 2692 4601 2768
rect 4582 2482 4585 2488
rect 4482 2448 4486 2451
rect 4370 2438 4374 2441
rect 4318 2392 4321 2408
rect 4210 2388 4214 2391
rect 4430 2382 4433 2418
rect 4218 2368 4222 2371
rect 4274 2368 4278 2371
rect 4238 2362 4241 2368
rect 4186 2358 4190 2361
rect 4158 2332 4161 2338
rect 4166 2332 4169 2338
rect 4006 2282 4009 2328
rect 4082 2318 4086 2321
rect 4080 2303 4082 2307
rect 4086 2303 4089 2307
rect 4093 2303 4096 2307
rect 4166 2282 4169 2328
rect 4190 2322 4193 2338
rect 3874 2278 3878 2281
rect 3978 2278 3982 2281
rect 3966 2272 3969 2278
rect 3938 2268 3942 2271
rect 4090 2268 4094 2271
rect 3910 2262 3913 2268
rect 3974 2262 3977 2268
rect 3818 2258 3822 2261
rect 3606 2252 3609 2258
rect 3654 2252 3657 2258
rect 3894 2252 3897 2258
rect 3562 2248 3566 2251
rect 3626 2248 3630 2251
rect 3946 2248 3950 2251
rect 3568 2203 3570 2207
rect 3574 2203 3577 2207
rect 3581 2203 3584 2207
rect 3534 2158 3545 2161
rect 3534 2082 3537 2158
rect 3542 2142 3545 2148
rect 3558 2142 3561 2148
rect 3590 2132 3593 2178
rect 3598 2162 3601 2168
rect 3606 2142 3609 2148
rect 3622 2132 3625 2158
rect 3638 2132 3641 2218
rect 3750 2192 3753 2238
rect 3818 2228 3822 2231
rect 3870 2192 3873 2208
rect 3762 2168 3766 2171
rect 3662 2152 3665 2168
rect 3702 2162 3705 2168
rect 3790 2162 3793 2168
rect 3950 2162 3953 2238
rect 3714 2158 3718 2161
rect 3778 2158 3782 2161
rect 3810 2158 3814 2161
rect 3830 2152 3833 2158
rect 3722 2148 3726 2151
rect 3762 2148 3766 2151
rect 3794 2148 3798 2151
rect 3898 2148 3902 2151
rect 3922 2148 3926 2151
rect 3646 2142 3649 2148
rect 3670 2142 3673 2148
rect 3678 2132 3681 2138
rect 3734 2132 3737 2148
rect 3814 2142 3817 2148
rect 3822 2142 3825 2148
rect 3862 2142 3865 2148
rect 3934 2142 3937 2148
rect 3974 2142 3977 2168
rect 3982 2152 3985 2188
rect 3746 2138 3750 2141
rect 3850 2138 3854 2141
rect 3990 2141 3993 2218
rect 4006 2192 4009 2268
rect 4014 2242 4017 2248
rect 4022 2232 4025 2268
rect 4110 2262 4113 2278
rect 4118 2262 4121 2268
rect 4134 2262 4137 2268
rect 4042 2258 4046 2261
rect 4170 2258 4174 2261
rect 4070 2252 4073 2258
rect 4030 2232 4033 2248
rect 4046 2242 4049 2248
rect 4062 2242 4065 2248
rect 4030 2222 4033 2228
rect 4014 2192 4017 2198
rect 4038 2172 4041 2218
rect 4078 2212 4081 2258
rect 4122 2248 4126 2251
rect 4094 2202 4097 2248
rect 4146 2238 4150 2241
rect 4126 2222 4129 2238
rect 4158 2222 4161 2248
rect 4174 2242 4177 2248
rect 4002 2148 4006 2151
rect 3982 2138 3993 2141
rect 3782 2132 3785 2138
rect 3562 2128 3566 2131
rect 3842 2128 3846 2131
rect 3550 2092 3553 2128
rect 3518 2062 3521 2068
rect 3410 2058 3414 2061
rect 3466 2058 3470 2061
rect 3350 2022 3353 2058
rect 3382 2052 3385 2058
rect 3370 2048 3374 2051
rect 3270 1882 3273 2018
rect 3286 1942 3289 1948
rect 3270 1822 3273 1858
rect 3262 1742 3265 1748
rect 3270 1742 3273 1758
rect 3278 1752 3281 1938
rect 3294 1882 3297 1948
rect 3302 1942 3305 1958
rect 3374 1952 3377 1958
rect 3322 1948 3326 1951
rect 3346 1938 3350 1941
rect 3302 1922 3305 1938
rect 3294 1851 3297 1868
rect 3310 1862 3313 1918
rect 3318 1882 3321 1938
rect 3334 1922 3337 1938
rect 3350 1902 3353 1938
rect 3370 1928 3374 1931
rect 3358 1872 3361 1918
rect 3390 1872 3393 2058
rect 3442 2048 3446 2051
rect 3398 2012 3401 2048
rect 3454 1982 3457 2058
rect 3542 2052 3545 2078
rect 3574 2072 3577 2128
rect 3622 2092 3625 2128
rect 3646 2122 3649 2128
rect 3630 2072 3633 2118
rect 3638 2072 3641 2078
rect 3654 2072 3657 2118
rect 3694 2112 3697 2128
rect 3702 2122 3705 2128
rect 3710 2092 3713 2118
rect 3690 2078 3694 2081
rect 3678 2072 3681 2078
rect 3718 2072 3721 2078
rect 3766 2072 3769 2118
rect 3814 2092 3817 2098
rect 3782 2072 3785 2088
rect 3814 2072 3817 2088
rect 3826 2078 3830 2081
rect 3610 2068 3614 2071
rect 3698 2068 3702 2071
rect 3746 2068 3750 2071
rect 3654 2062 3657 2068
rect 3766 2062 3769 2068
rect 3846 2062 3849 2078
rect 3854 2062 3857 2138
rect 3902 2132 3905 2138
rect 3870 2128 3878 2131
rect 3914 2128 3918 2131
rect 3862 2092 3865 2098
rect 3870 2082 3873 2128
rect 3966 2122 3969 2128
rect 3878 2092 3881 2108
rect 3974 2082 3977 2098
rect 3894 2062 3897 2078
rect 3958 2072 3961 2078
rect 3594 2058 3598 2061
rect 3690 2058 3694 2061
rect 3722 2058 3726 2061
rect 3454 1962 3457 1978
rect 3494 1962 3497 2038
rect 3558 1972 3561 2058
rect 3630 2052 3633 2058
rect 3578 2048 3582 2051
rect 3618 2048 3622 2051
rect 3618 2018 3622 2021
rect 3568 2003 3570 2007
rect 3574 2003 3577 2007
rect 3581 2003 3584 2007
rect 3538 1968 3542 1971
rect 3518 1962 3521 1968
rect 3426 1948 3430 1951
rect 3414 1932 3417 1938
rect 3398 1862 3401 1868
rect 3378 1858 3382 1861
rect 3406 1861 3409 1928
rect 3422 1872 3425 1948
rect 3434 1938 3438 1941
rect 3430 1872 3433 1938
rect 3438 1922 3441 1928
rect 3406 1858 3414 1861
rect 3294 1848 3334 1851
rect 3286 1842 3289 1848
rect 3306 1818 3310 1821
rect 3326 1812 3329 1818
rect 3302 1762 3305 1788
rect 3342 1772 3345 1858
rect 3350 1842 3353 1858
rect 3350 1762 3353 1838
rect 3358 1792 3361 1828
rect 3390 1801 3393 1858
rect 3386 1798 3393 1801
rect 3398 1802 3401 1858
rect 3454 1852 3457 1918
rect 3470 1862 3473 1938
rect 3486 1872 3489 1958
rect 3518 1942 3521 1958
rect 3542 1942 3545 1948
rect 3498 1938 3502 1941
rect 3534 1932 3537 1938
rect 3494 1862 3497 1918
rect 3466 1858 3470 1861
rect 3510 1852 3513 1858
rect 3414 1842 3417 1848
rect 3518 1842 3521 1918
rect 3534 1862 3537 1928
rect 3550 1882 3553 1968
rect 3558 1942 3561 1968
rect 3614 1962 3617 1978
rect 3594 1948 3598 1951
rect 3550 1872 3553 1878
rect 3582 1872 3585 1938
rect 3606 1881 3609 1918
rect 3630 1882 3633 2048
rect 3678 1992 3681 2058
rect 3758 2051 3761 2058
rect 3774 2052 3777 2058
rect 3758 2048 3766 2051
rect 3790 2042 3793 2058
rect 3802 2048 3806 2051
rect 3774 2002 3777 2038
rect 3782 2032 3785 2038
rect 3782 1992 3785 2028
rect 3690 1988 3694 1991
rect 3654 1952 3657 1958
rect 3638 1932 3641 1948
rect 3662 1942 3665 1948
rect 3670 1942 3673 1978
rect 3706 1968 3710 1971
rect 3718 1962 3721 1968
rect 3714 1948 3718 1951
rect 3746 1948 3750 1951
rect 3746 1938 3750 1941
rect 3722 1928 3726 1931
rect 3606 1878 3614 1881
rect 3630 1872 3633 1878
rect 3574 1862 3577 1868
rect 3638 1862 3641 1928
rect 3646 1912 3649 1918
rect 3678 1882 3681 1918
rect 3686 1912 3689 1928
rect 3718 1882 3721 1908
rect 3734 1882 3737 1918
rect 3750 1882 3753 1938
rect 3758 1932 3761 1938
rect 3738 1878 3745 1881
rect 3710 1872 3713 1878
rect 3734 1862 3737 1878
rect 3674 1858 3678 1861
rect 3566 1852 3569 1858
rect 3470 1832 3473 1838
rect 3574 1822 3577 1858
rect 3598 1832 3601 1858
rect 3638 1852 3641 1858
rect 3654 1852 3657 1858
rect 3358 1772 3361 1788
rect 3290 1758 3294 1761
rect 3314 1758 3318 1761
rect 3302 1742 3305 1748
rect 3318 1742 3321 1748
rect 3326 1692 3329 1758
rect 3338 1748 3342 1751
rect 3334 1732 3337 1738
rect 3274 1678 3278 1681
rect 3342 1672 3345 1748
rect 3366 1742 3369 1788
rect 3390 1742 3393 1758
rect 3406 1742 3409 1748
rect 3414 1742 3417 1758
rect 3430 1752 3433 1818
rect 3494 1812 3497 1818
rect 3446 1762 3449 1808
rect 3466 1758 3470 1761
rect 3486 1742 3489 1798
rect 3526 1762 3529 1798
rect 3510 1752 3513 1758
rect 3506 1748 3510 1751
rect 3418 1738 3422 1741
rect 3490 1738 3494 1741
rect 3370 1728 3374 1731
rect 3382 1712 3385 1718
rect 3398 1702 3401 1718
rect 3438 1702 3441 1718
rect 3358 1662 3361 1698
rect 3402 1678 3406 1681
rect 3402 1668 3406 1671
rect 3222 1658 3230 1661
rect 3394 1658 3398 1661
rect 3214 1622 3217 1648
rect 3238 1632 3241 1638
rect 3238 1552 3241 1598
rect 3270 1592 3273 1658
rect 3310 1642 3313 1658
rect 3318 1652 3321 1658
rect 3326 1642 3329 1648
rect 3294 1592 3297 1628
rect 3302 1622 3305 1628
rect 3218 1548 3222 1551
rect 3270 1542 3273 1588
rect 3302 1562 3305 1618
rect 3310 1582 3313 1618
rect 3282 1558 3286 1561
rect 3282 1548 3286 1551
rect 3310 1542 3313 1578
rect 3318 1562 3321 1568
rect 3342 1552 3345 1658
rect 3218 1538 3222 1541
rect 3298 1538 3302 1541
rect 3114 1478 3118 1481
rect 3174 1472 3177 1488
rect 3122 1468 3126 1471
rect 3094 1462 3097 1468
rect 3114 1458 3118 1461
rect 3062 1382 3065 1418
rect 3094 1392 3097 1448
rect 3062 1352 3065 1358
rect 3110 1352 3113 1388
rect 3118 1382 3121 1458
rect 3142 1432 3145 1448
rect 3126 1362 3129 1418
rect 3142 1392 3145 1428
rect 3150 1402 3153 1448
rect 3166 1382 3169 1468
rect 3198 1462 3201 1468
rect 3186 1458 3190 1461
rect 3206 1452 3209 1458
rect 3198 1442 3201 1448
rect 3198 1382 3201 1388
rect 3134 1362 3137 1368
rect 3166 1362 3169 1378
rect 3178 1358 3182 1361
rect 3118 1352 3121 1358
rect 3034 1348 3038 1351
rect 3186 1348 3190 1351
rect 3046 1342 3049 1348
rect 3038 1312 3041 1338
rect 3048 1303 3050 1307
rect 3054 1303 3057 1307
rect 3061 1303 3064 1307
rect 3006 1272 3009 1288
rect 3014 1272 3017 1278
rect 3070 1272 3073 1318
rect 2898 1268 2902 1271
rect 2990 1262 2993 1268
rect 3030 1262 3033 1268
rect 2898 1258 2902 1261
rect 2914 1258 2918 1261
rect 2926 1252 2929 1258
rect 2890 1248 2894 1251
rect 2918 1232 2921 1248
rect 2942 1242 2945 1248
rect 2950 1242 2953 1258
rect 2958 1222 2961 1258
rect 3038 1252 3041 1258
rect 3062 1252 3065 1258
rect 2894 1192 2897 1218
rect 2990 1212 2993 1248
rect 3002 1238 3006 1241
rect 3006 1222 3009 1238
rect 2878 1168 2886 1171
rect 2862 1162 2865 1168
rect 2910 1162 2913 1188
rect 2930 1158 2937 1161
rect 2878 1142 2881 1148
rect 2910 1142 2913 1158
rect 2934 1152 2937 1158
rect 2922 1148 2926 1151
rect 2886 1092 2889 1138
rect 2902 1122 2905 1128
rect 2738 1088 2742 1091
rect 2810 1078 2814 1081
rect 2582 1068 2590 1071
rect 2582 1062 2585 1068
rect 2614 1062 2617 1068
rect 2590 1052 2593 1058
rect 2574 952 2577 988
rect 2514 948 2518 951
rect 2550 942 2553 948
rect 2582 942 2585 968
rect 2598 952 2601 1048
rect 2614 952 2617 1038
rect 2638 1012 2641 1078
rect 2678 1072 2681 1078
rect 2658 1068 2662 1071
rect 2682 1068 2686 1071
rect 2650 1058 2654 1061
rect 2694 1052 2697 1058
rect 2702 1052 2705 1058
rect 2634 998 2641 1001
rect 2638 992 2641 998
rect 2626 958 2630 961
rect 2646 952 2649 1018
rect 2606 942 2609 948
rect 2506 938 2521 941
rect 2490 928 2494 931
rect 2502 922 2505 928
rect 2446 892 2449 918
rect 2470 882 2473 908
rect 2430 878 2441 881
rect 2422 852 2425 858
rect 2414 792 2417 838
rect 2430 772 2433 868
rect 2430 752 2433 768
rect 2390 742 2393 748
rect 2382 712 2385 728
rect 2398 692 2401 738
rect 2438 732 2441 878
rect 2518 872 2521 938
rect 2534 922 2537 938
rect 2646 932 2649 938
rect 2654 932 2657 998
rect 2670 992 2673 1018
rect 2710 1002 2713 1078
rect 2774 1072 2777 1078
rect 2822 1072 2825 1078
rect 2718 1022 2721 1068
rect 2726 1062 2729 1068
rect 2750 1012 2753 1048
rect 2766 1042 2769 1058
rect 2774 1022 2777 1068
rect 2782 1062 2785 1068
rect 2798 1062 2801 1068
rect 2818 1058 2822 1061
rect 2670 952 2673 958
rect 2678 952 2681 978
rect 2710 952 2713 978
rect 2774 952 2777 998
rect 2790 992 2793 1038
rect 2586 928 2590 931
rect 2538 888 2542 891
rect 2550 872 2553 878
rect 2598 872 2601 888
rect 2482 868 2486 871
rect 2578 868 2582 871
rect 2634 868 2638 871
rect 2454 852 2457 868
rect 2462 842 2465 858
rect 2494 852 2497 858
rect 2474 838 2478 841
rect 2446 762 2449 838
rect 2502 782 2505 868
rect 2510 862 2513 868
rect 2534 852 2537 858
rect 2526 842 2529 848
rect 2518 802 2521 828
rect 2418 728 2422 731
rect 2418 688 2422 691
rect 2342 672 2345 678
rect 2358 662 2361 668
rect 2398 662 2401 678
rect 2438 672 2441 728
rect 2446 692 2449 758
rect 2478 752 2481 768
rect 2486 752 2489 758
rect 2518 752 2521 798
rect 2534 762 2537 848
rect 2606 842 2609 858
rect 2638 852 2641 858
rect 2626 848 2630 851
rect 2614 842 2617 848
rect 2544 803 2546 807
rect 2550 803 2553 807
rect 2557 803 2560 807
rect 2582 802 2585 818
rect 2578 778 2582 781
rect 2594 768 2598 771
rect 2606 761 2609 838
rect 2614 792 2617 838
rect 2598 758 2609 761
rect 2470 742 2473 748
rect 2494 732 2497 748
rect 2550 742 2553 748
rect 2454 682 2457 728
rect 2430 662 2433 668
rect 2322 658 2326 661
rect 2330 658 2342 661
rect 2382 652 2385 658
rect 2454 652 2457 678
rect 2438 592 2441 598
rect 2342 562 2345 568
rect 2318 552 2321 558
rect 2266 538 2270 541
rect 2286 522 2289 528
rect 2254 472 2257 508
rect 2166 318 2174 321
rect 2166 292 2169 318
rect 2110 272 2113 288
rect 2134 272 2137 278
rect 2142 272 2145 288
rect 2170 268 2174 271
rect 2134 262 2137 268
rect 2190 262 2193 268
rect 2002 258 2006 261
rect 2042 258 2046 261
rect 2114 258 2118 261
rect 2086 252 2089 258
rect 2094 252 2097 258
rect 2158 252 2161 258
rect 1962 248 1966 251
rect 2178 248 2182 251
rect 2198 242 2201 248
rect 1974 192 1977 198
rect 1886 82 1889 88
rect 1918 72 1921 78
rect 1870 62 1873 68
rect 1942 62 1945 158
rect 1982 142 1985 238
rect 2046 162 2049 178
rect 2002 148 2006 151
rect 2062 142 2065 148
rect 2078 142 2081 148
rect 1982 132 1985 138
rect 1950 92 1953 108
rect 1974 72 1977 128
rect 1998 92 2001 118
rect 2002 78 2006 81
rect 1982 72 1985 78
rect 2014 61 2017 138
rect 2078 112 2081 128
rect 2094 122 2097 158
rect 2102 152 2105 178
rect 2024 103 2026 107
rect 2030 103 2033 107
rect 2037 103 2040 107
rect 2046 92 2049 98
rect 2062 62 2065 88
rect 2078 82 2081 108
rect 2070 62 2073 68
rect 2094 62 2097 118
rect 2110 92 2113 238
rect 2126 182 2129 228
rect 2190 182 2193 218
rect 2206 212 2209 338
rect 2218 328 2222 331
rect 2222 292 2225 298
rect 2230 272 2233 328
rect 2238 272 2241 348
rect 2254 332 2257 458
rect 2262 452 2265 468
rect 2270 462 2273 508
rect 2278 472 2281 518
rect 2294 511 2297 528
rect 2286 508 2297 511
rect 2326 512 2329 558
rect 2350 542 2353 578
rect 2426 568 2430 571
rect 2358 558 2366 561
rect 2358 552 2361 558
rect 2390 552 2393 568
rect 2454 562 2457 608
rect 2462 582 2465 718
rect 2494 712 2497 728
rect 2510 722 2513 728
rect 2498 688 2502 691
rect 2518 682 2521 688
rect 2510 672 2513 678
rect 2490 658 2494 661
rect 2470 592 2473 618
rect 2370 548 2377 551
rect 2374 542 2377 548
rect 2462 551 2465 568
rect 2470 561 2473 588
rect 2470 558 2481 561
rect 2462 548 2470 551
rect 2382 542 2385 548
rect 2362 538 2369 541
rect 2390 538 2398 541
rect 2286 492 2289 508
rect 2306 488 2310 491
rect 2294 462 2297 478
rect 2342 472 2345 538
rect 2366 492 2369 538
rect 2382 522 2385 528
rect 2378 478 2382 481
rect 2342 462 2345 468
rect 2318 452 2321 458
rect 2290 448 2297 451
rect 2262 362 2265 368
rect 2254 272 2257 308
rect 2262 302 2265 348
rect 2278 342 2281 348
rect 2286 342 2289 378
rect 2266 268 2270 271
rect 2214 262 2217 268
rect 2230 262 2233 268
rect 2278 262 2281 338
rect 2294 331 2297 448
rect 2326 402 2329 448
rect 2342 412 2345 458
rect 2350 392 2353 468
rect 2358 462 2361 478
rect 2382 442 2385 458
rect 2390 441 2393 538
rect 2406 532 2409 548
rect 2438 542 2441 548
rect 2398 528 2406 531
rect 2398 482 2401 528
rect 2414 492 2417 508
rect 2406 482 2409 488
rect 2438 472 2441 538
rect 2402 468 2406 471
rect 2418 468 2422 471
rect 2386 438 2393 441
rect 2302 362 2305 368
rect 2414 362 2417 458
rect 2438 452 2441 458
rect 2446 431 2449 518
rect 2470 492 2473 508
rect 2478 502 2481 558
rect 2486 552 2489 648
rect 2494 642 2497 648
rect 2506 558 2510 561
rect 2494 551 2497 558
rect 2494 548 2510 551
rect 2494 532 2497 538
rect 2502 502 2505 548
rect 2510 502 2513 518
rect 2478 491 2481 498
rect 2518 492 2521 658
rect 2542 652 2545 718
rect 2550 672 2553 738
rect 2558 662 2561 758
rect 2566 662 2569 758
rect 2586 748 2590 751
rect 2574 662 2577 708
rect 2598 692 2601 758
rect 2622 742 2625 798
rect 2646 772 2649 818
rect 2654 762 2657 928
rect 2662 892 2665 898
rect 2662 842 2665 848
rect 2670 771 2673 928
rect 2678 872 2681 938
rect 2698 928 2702 931
rect 2742 922 2745 948
rect 2798 942 2801 948
rect 2806 942 2809 1058
rect 2822 962 2825 968
rect 2830 952 2833 1088
rect 2846 1022 2849 1088
rect 2910 1082 2913 1088
rect 2926 1072 2929 1088
rect 2934 1082 2937 1138
rect 2958 1132 2961 1158
rect 2966 1152 2969 1188
rect 2982 1152 2985 1198
rect 3030 1192 3033 1228
rect 3018 1188 3022 1191
rect 3006 1181 3009 1188
rect 3006 1178 3041 1181
rect 3030 1162 3033 1168
rect 3038 1162 3041 1178
rect 3054 1162 3057 1218
rect 3078 1192 3081 1338
rect 3110 1272 3113 1298
rect 3118 1272 3121 1348
rect 3126 1292 3129 1298
rect 3134 1292 3137 1348
rect 3150 1342 3153 1348
rect 3214 1332 3217 1518
rect 3246 1492 3249 1538
rect 3262 1532 3265 1538
rect 3254 1472 3257 1528
rect 3234 1468 3238 1471
rect 3246 1462 3249 1468
rect 3222 1442 3225 1448
rect 3230 1392 3233 1458
rect 3254 1352 3257 1468
rect 3262 1462 3265 1498
rect 3318 1472 3321 1548
rect 3350 1542 3353 1548
rect 3330 1538 3334 1541
rect 3334 1512 3337 1528
rect 3302 1462 3305 1468
rect 3318 1462 3321 1468
rect 3346 1458 3350 1461
rect 3270 1452 3273 1458
rect 3278 1452 3281 1458
rect 3290 1438 3294 1441
rect 3326 1412 3329 1458
rect 3342 1412 3345 1418
rect 3262 1362 3265 1378
rect 3170 1328 3174 1331
rect 3206 1322 3209 1328
rect 3162 1318 3166 1321
rect 3118 1262 3121 1268
rect 3158 1262 3161 1288
rect 3174 1282 3177 1288
rect 3182 1281 3185 1318
rect 3190 1292 3193 1308
rect 3178 1278 3185 1281
rect 3146 1258 3150 1261
rect 3102 1252 3105 1258
rect 3158 1252 3161 1258
rect 3090 1248 3094 1251
rect 3138 1248 3142 1251
rect 3166 1241 3169 1268
rect 3174 1262 3177 1268
rect 3158 1238 3169 1241
rect 3014 1142 3017 1158
rect 3094 1152 3097 1218
rect 3110 1158 3118 1161
rect 3110 1152 3113 1158
rect 3042 1148 3046 1151
rect 3126 1142 3129 1158
rect 3150 1152 3153 1198
rect 3158 1181 3161 1238
rect 3174 1192 3177 1218
rect 3214 1192 3217 1328
rect 3230 1322 3233 1348
rect 3262 1342 3265 1348
rect 3282 1338 3286 1341
rect 3294 1332 3297 1338
rect 3310 1332 3313 1348
rect 3278 1328 3286 1331
rect 3238 1282 3241 1288
rect 3234 1268 3238 1271
rect 3222 1232 3225 1258
rect 3170 1188 3174 1191
rect 3158 1178 3169 1181
rect 2994 1138 2998 1141
rect 3098 1138 3102 1141
rect 3154 1138 3158 1141
rect 2942 1122 2945 1128
rect 2974 1122 2977 1138
rect 2990 1122 2993 1128
rect 3010 1118 3014 1121
rect 3070 1112 3073 1138
rect 2958 1081 2961 1108
rect 3048 1103 3050 1107
rect 3054 1103 3057 1107
rect 3061 1103 3064 1107
rect 3070 1092 3073 1108
rect 3086 1092 3089 1118
rect 2954 1078 2961 1081
rect 2898 1068 2902 1071
rect 2886 1062 2889 1068
rect 2974 1062 2977 1088
rect 3110 1082 3113 1088
rect 3118 1072 3121 1128
rect 3134 1102 3137 1118
rect 3002 1068 3006 1071
rect 3026 1068 3030 1071
rect 3014 1062 3017 1068
rect 3054 1062 3057 1068
rect 2874 1058 2878 1061
rect 2922 1058 2926 1061
rect 3026 1058 3030 1061
rect 2838 972 2841 1018
rect 2822 942 2825 948
rect 2694 912 2697 918
rect 2694 892 2697 908
rect 2750 892 2753 938
rect 2766 922 2769 938
rect 2782 932 2785 938
rect 2806 932 2809 938
rect 2846 932 2849 1018
rect 2862 982 2865 1038
rect 2870 1032 2873 1048
rect 2878 982 2881 1048
rect 2886 992 2889 1058
rect 2902 1032 2905 1048
rect 2934 1002 2937 1058
rect 2954 1038 2966 1041
rect 2974 1032 2977 1048
rect 2990 1042 2993 1058
rect 2950 1022 2953 1028
rect 2910 962 2913 968
rect 2882 948 2886 951
rect 2870 942 2873 948
rect 2882 938 2886 941
rect 2854 932 2857 938
rect 2894 932 2897 958
rect 2906 948 2910 951
rect 2906 938 2913 941
rect 2922 938 2926 941
rect 2882 928 2886 931
rect 2714 888 2718 891
rect 2686 872 2689 878
rect 2686 802 2689 868
rect 2722 858 2726 861
rect 2702 842 2705 858
rect 2734 852 2737 858
rect 2742 852 2745 868
rect 2722 838 2726 841
rect 2670 768 2681 771
rect 2670 752 2673 758
rect 2678 752 2681 768
rect 2694 762 2697 808
rect 2702 792 2705 838
rect 2726 752 2729 808
rect 2750 772 2753 858
rect 2758 851 2761 918
rect 2838 912 2841 918
rect 2846 892 2849 928
rect 2862 922 2865 928
rect 2770 878 2830 881
rect 2770 868 2774 871
rect 2802 868 2806 871
rect 2882 868 2886 871
rect 2778 858 2782 861
rect 2758 848 2766 851
rect 2814 822 2817 838
rect 2822 832 2825 848
rect 2782 772 2785 818
rect 2814 762 2817 818
rect 2830 792 2833 858
rect 2838 852 2841 858
rect 2846 782 2849 868
rect 2910 862 2913 938
rect 2942 882 2945 1018
rect 2950 992 2953 1018
rect 2966 962 2969 968
rect 2950 942 2953 948
rect 2974 942 2977 1018
rect 2982 942 2985 1038
rect 3014 981 3017 1018
rect 3006 978 3017 981
rect 2994 958 2998 961
rect 2994 948 2998 951
rect 2958 921 2961 938
rect 2966 932 2969 938
rect 2958 918 2969 921
rect 2966 892 2969 918
rect 2966 872 2969 888
rect 2858 858 2862 861
rect 2858 848 2862 851
rect 2802 758 2806 761
rect 2734 752 2737 758
rect 2658 748 2662 751
rect 2786 748 2790 751
rect 2678 742 2681 748
rect 2694 742 2697 748
rect 2726 742 2729 748
rect 2666 738 2670 741
rect 2714 738 2718 741
rect 2738 738 2742 741
rect 2786 738 2790 741
rect 2614 732 2617 738
rect 2606 712 2609 728
rect 2622 711 2625 738
rect 2614 708 2625 711
rect 2646 712 2649 738
rect 2702 731 2705 738
rect 2702 728 2713 731
rect 2582 672 2585 678
rect 2614 672 2617 708
rect 2622 692 2625 698
rect 2654 682 2657 688
rect 2526 522 2529 618
rect 2574 612 2577 618
rect 2544 603 2546 607
rect 2550 603 2553 607
rect 2557 603 2560 607
rect 2606 592 2609 658
rect 2614 592 2617 638
rect 2630 582 2633 658
rect 2654 652 2657 668
rect 2662 662 2665 728
rect 2690 718 2694 721
rect 2678 692 2681 708
rect 2710 692 2713 728
rect 2686 682 2689 688
rect 2718 682 2721 688
rect 2662 602 2665 658
rect 2670 592 2673 678
rect 2734 672 2737 698
rect 2742 692 2745 698
rect 2750 682 2753 718
rect 2766 672 2769 728
rect 2798 712 2801 738
rect 2782 672 2785 688
rect 2806 672 2809 728
rect 2822 722 2825 738
rect 2830 692 2833 748
rect 2846 731 2849 758
rect 2870 752 2873 818
rect 2894 792 2897 818
rect 2858 748 2862 751
rect 2858 738 2862 741
rect 2878 732 2881 768
rect 2906 758 2910 761
rect 2886 742 2889 748
rect 2846 728 2857 731
rect 2846 672 2849 708
rect 2854 702 2857 728
rect 2802 668 2806 671
rect 2702 662 2705 668
rect 2686 658 2694 661
rect 2778 658 2782 661
rect 2822 658 2830 661
rect 2630 562 2633 578
rect 2662 562 2665 588
rect 2650 558 2654 561
rect 2574 552 2577 558
rect 2598 552 2601 558
rect 2538 538 2542 541
rect 2574 532 2577 538
rect 2582 532 2585 538
rect 2538 528 2542 531
rect 2542 522 2545 528
rect 2478 488 2489 491
rect 2486 482 2489 488
rect 2474 478 2478 481
rect 2454 472 2457 478
rect 2498 468 2502 471
rect 2438 428 2449 431
rect 2462 462 2465 468
rect 2510 462 2513 468
rect 2422 392 2425 428
rect 2438 362 2441 428
rect 2446 382 2449 418
rect 2446 362 2449 368
rect 2462 362 2465 458
rect 2494 451 2497 458
rect 2494 448 2518 451
rect 2534 432 2537 458
rect 2542 432 2545 468
rect 2566 452 2569 498
rect 2574 461 2577 528
rect 2598 522 2601 548
rect 2606 512 2609 538
rect 2614 532 2617 548
rect 2654 542 2657 548
rect 2634 538 2638 541
rect 2590 481 2593 508
rect 2590 478 2601 481
rect 2598 472 2601 478
rect 2586 468 2590 471
rect 2598 462 2601 468
rect 2606 462 2609 498
rect 2630 472 2633 508
rect 2638 462 2641 528
rect 2662 502 2665 558
rect 2686 552 2689 658
rect 2710 592 2713 648
rect 2726 642 2729 658
rect 2822 652 2825 658
rect 2754 648 2758 651
rect 2786 648 2790 651
rect 2702 552 2705 558
rect 2674 538 2678 541
rect 2686 532 2689 548
rect 2726 542 2729 578
rect 2758 562 2761 568
rect 2738 558 2742 561
rect 2798 561 2801 618
rect 2814 572 2817 648
rect 2830 642 2833 648
rect 2794 558 2801 561
rect 2822 562 2825 568
rect 2774 552 2777 558
rect 2830 552 2833 568
rect 2802 548 2806 551
rect 2734 542 2737 548
rect 2770 538 2774 541
rect 2802 538 2806 541
rect 2794 528 2798 531
rect 2654 462 2657 468
rect 2662 462 2665 488
rect 2670 482 2673 498
rect 2678 471 2681 508
rect 2686 492 2689 528
rect 2678 468 2686 471
rect 2574 458 2582 461
rect 2670 452 2673 468
rect 2694 462 2697 488
rect 2702 482 2705 508
rect 2822 502 2825 518
rect 2710 492 2713 498
rect 2790 492 2793 498
rect 2838 492 2841 598
rect 2846 592 2849 668
rect 2854 582 2857 618
rect 2862 542 2865 718
rect 2870 681 2873 718
rect 2894 712 2897 748
rect 2918 732 2921 858
rect 2926 852 2929 868
rect 2950 862 2953 868
rect 2958 822 2961 858
rect 2942 812 2945 818
rect 2974 792 2977 918
rect 2982 872 2985 938
rect 2982 852 2985 858
rect 2998 852 3001 938
rect 3006 862 3009 978
rect 3014 962 3017 968
rect 3038 952 3041 1018
rect 3062 992 3065 1058
rect 3094 1052 3097 1058
rect 3054 952 3057 958
rect 3030 948 3038 951
rect 3030 942 3033 948
rect 3050 938 3054 941
rect 3030 912 3033 928
rect 3048 903 3050 907
rect 3054 903 3057 907
rect 3061 903 3064 907
rect 3070 892 3073 1008
rect 3086 922 3089 1048
rect 3098 1038 3102 1041
rect 3094 952 3097 958
rect 3102 952 3105 968
rect 3106 938 3110 941
rect 3038 872 3041 878
rect 3046 872 3049 888
rect 3078 872 3081 918
rect 3026 868 3030 871
rect 3094 862 3097 938
rect 3106 928 3110 931
rect 3118 892 3121 1058
rect 3126 1052 3129 1058
rect 3142 1052 3145 1108
rect 3150 1052 3153 1068
rect 3158 1062 3161 1088
rect 3166 1072 3169 1178
rect 3186 1158 3190 1161
rect 3230 1152 3233 1238
rect 3246 1161 3249 1318
rect 3278 1282 3281 1328
rect 3318 1322 3321 1358
rect 3334 1342 3337 1348
rect 3334 1312 3337 1338
rect 3290 1288 3294 1291
rect 3278 1272 3281 1278
rect 3334 1272 3337 1308
rect 3298 1268 3302 1271
rect 3270 1252 3273 1268
rect 3314 1248 3318 1251
rect 3254 1172 3257 1248
rect 3242 1158 3249 1161
rect 3262 1162 3265 1218
rect 3186 1138 3190 1141
rect 3174 1082 3177 1098
rect 3174 1062 3177 1078
rect 3190 1072 3193 1098
rect 3198 1072 3201 1138
rect 3254 1132 3257 1138
rect 3238 1112 3241 1118
rect 3262 1112 3265 1118
rect 3270 1092 3273 1158
rect 3278 1152 3281 1188
rect 3294 1162 3297 1198
rect 3310 1142 3313 1148
rect 3318 1142 3321 1228
rect 3342 1201 3345 1318
rect 3350 1282 3353 1448
rect 3358 1372 3361 1558
rect 3366 1552 3369 1618
rect 3414 1592 3417 1638
rect 3390 1552 3393 1588
rect 3422 1562 3425 1698
rect 3438 1672 3441 1678
rect 3454 1672 3457 1708
rect 3434 1658 3441 1661
rect 3450 1658 3454 1661
rect 3430 1642 3433 1648
rect 3438 1642 3441 1658
rect 3450 1578 3454 1581
rect 3406 1552 3409 1558
rect 3366 1471 3369 1548
rect 3374 1512 3377 1518
rect 3398 1492 3401 1548
rect 3446 1542 3449 1548
rect 3426 1538 3430 1541
rect 3454 1532 3457 1538
rect 3462 1532 3465 1678
rect 3470 1662 3473 1738
rect 3494 1722 3497 1728
rect 3478 1682 3481 1718
rect 3518 1712 3521 1738
rect 3478 1672 3481 1678
rect 3526 1671 3529 1758
rect 3534 1752 3537 1818
rect 3568 1803 3570 1807
rect 3574 1803 3577 1807
rect 3581 1803 3584 1807
rect 3550 1792 3553 1798
rect 3570 1748 3574 1751
rect 3546 1738 3550 1741
rect 3574 1732 3577 1738
rect 3538 1728 3542 1731
rect 3518 1668 3529 1671
rect 3518 1662 3521 1668
rect 3534 1662 3537 1708
rect 3542 1662 3545 1678
rect 3574 1662 3577 1728
rect 3590 1702 3593 1818
rect 3598 1792 3601 1828
rect 3622 1792 3625 1818
rect 3598 1742 3601 1758
rect 3610 1748 3617 1751
rect 3614 1732 3617 1748
rect 3622 1742 3625 1758
rect 3630 1752 3633 1758
rect 3638 1748 3646 1751
rect 3638 1741 3641 1748
rect 3634 1738 3641 1741
rect 3614 1692 3617 1728
rect 3646 1712 3649 1728
rect 3654 1712 3657 1848
rect 3678 1762 3681 1818
rect 3734 1812 3737 1818
rect 3678 1742 3681 1748
rect 3638 1668 3646 1671
rect 3470 1592 3473 1658
rect 3494 1652 3497 1658
rect 3502 1602 3505 1618
rect 3494 1562 3497 1568
rect 3490 1548 3494 1551
rect 3378 1488 3382 1491
rect 3366 1468 3398 1471
rect 3406 1462 3409 1488
rect 3454 1471 3457 1528
rect 3462 1482 3465 1528
rect 3454 1468 3462 1471
rect 3394 1458 3398 1461
rect 3358 1352 3361 1368
rect 3366 1342 3369 1388
rect 3374 1362 3377 1378
rect 3378 1348 3382 1351
rect 3366 1272 3369 1288
rect 3390 1262 3393 1338
rect 3398 1302 3401 1338
rect 3406 1302 3409 1418
rect 3414 1352 3417 1428
rect 3430 1402 3433 1468
rect 3470 1462 3473 1538
rect 3486 1502 3489 1548
rect 3450 1458 3454 1461
rect 3462 1458 3470 1461
rect 3438 1402 3441 1458
rect 3450 1448 3454 1451
rect 3430 1392 3433 1398
rect 3422 1352 3425 1358
rect 3430 1352 3433 1368
rect 3454 1352 3457 1418
rect 3430 1292 3433 1318
rect 3446 1292 3449 1328
rect 3398 1282 3401 1288
rect 3422 1282 3425 1288
rect 3446 1272 3449 1288
rect 3370 1258 3374 1261
rect 3406 1252 3409 1258
rect 3422 1251 3425 1258
rect 3422 1248 3433 1251
rect 3362 1238 3366 1241
rect 3430 1232 3433 1248
rect 3438 1232 3441 1258
rect 3342 1198 3350 1201
rect 3382 1162 3385 1218
rect 3398 1161 3401 1198
rect 3342 1142 3345 1158
rect 3350 1152 3353 1158
rect 3418 1158 3422 1161
rect 3282 1138 3286 1141
rect 3258 1068 3262 1071
rect 3182 1062 3185 1068
rect 3142 962 3145 1008
rect 3154 968 3158 971
rect 3126 942 3129 958
rect 3166 952 3169 1008
rect 3174 962 3177 968
rect 3190 952 3193 1068
rect 3238 1062 3241 1068
rect 3202 1058 3206 1061
rect 3218 1058 3222 1061
rect 3206 1021 3209 1058
rect 3214 1042 3217 1048
rect 3206 1018 3217 1021
rect 3198 1002 3201 1018
rect 3174 942 3177 948
rect 3162 938 3166 941
rect 3190 941 3193 948
rect 3182 938 3193 941
rect 3198 942 3201 968
rect 3138 868 3142 871
rect 3166 862 3169 868
rect 3174 862 3177 868
rect 3106 858 3110 861
rect 3130 858 3134 861
rect 3066 848 3070 851
rect 3106 848 3110 851
rect 3122 848 3126 851
rect 3162 848 3166 851
rect 3150 842 3153 848
rect 3182 842 3185 938
rect 3206 932 3209 1008
rect 3214 892 3217 1018
rect 3222 1002 3225 1048
rect 3246 1002 3249 1068
rect 3270 1052 3273 1058
rect 3262 982 3265 988
rect 3270 961 3273 1018
rect 3278 1012 3281 1078
rect 3270 958 3278 961
rect 3226 948 3230 951
rect 3258 948 3262 951
rect 3226 938 3230 941
rect 3226 928 3230 931
rect 3238 922 3241 928
rect 3194 888 3198 891
rect 3238 872 3241 888
rect 3226 868 3230 871
rect 3214 861 3217 868
rect 3246 862 3249 948
rect 3266 938 3270 941
rect 3282 928 3286 931
rect 3294 902 3297 1128
rect 3302 1112 3305 1138
rect 3366 1132 3369 1138
rect 3338 1128 3342 1131
rect 3326 1122 3329 1128
rect 3374 1092 3377 1128
rect 3382 1112 3385 1148
rect 3410 1138 3414 1141
rect 3430 1082 3433 1228
rect 3454 1202 3457 1348
rect 3462 1272 3465 1458
rect 3494 1452 3497 1518
rect 3502 1492 3505 1568
rect 3510 1542 3513 1658
rect 3526 1652 3529 1658
rect 3522 1548 3526 1551
rect 3534 1542 3537 1658
rect 3550 1551 3553 1618
rect 3568 1603 3570 1607
rect 3574 1603 3577 1607
rect 3581 1603 3584 1607
rect 3574 1562 3577 1578
rect 3542 1548 3553 1551
rect 3590 1552 3593 1658
rect 3630 1652 3633 1668
rect 3638 1622 3641 1668
rect 3650 1658 3654 1661
rect 3654 1632 3657 1648
rect 3630 1562 3633 1568
rect 3662 1552 3665 1678
rect 3670 1672 3673 1708
rect 3678 1671 3681 1718
rect 3686 1682 3689 1738
rect 3694 1722 3697 1738
rect 3702 1712 3705 1748
rect 3726 1742 3729 1748
rect 3742 1742 3745 1878
rect 3758 1872 3761 1918
rect 3766 1902 3769 1958
rect 3774 1902 3777 1928
rect 3766 1862 3769 1878
rect 3750 1852 3753 1858
rect 3782 1852 3785 1928
rect 3790 1912 3793 2018
rect 3806 1952 3809 1988
rect 3814 1972 3817 2058
rect 3842 2038 3846 2041
rect 3854 2002 3857 2058
rect 3926 2052 3929 2058
rect 3882 2048 3886 2051
rect 3834 1988 3838 1991
rect 3814 1962 3817 1968
rect 3826 1958 3830 1961
rect 3862 1952 3865 1998
rect 3894 1958 3902 1961
rect 3870 1952 3873 1958
rect 3894 1952 3897 1958
rect 3926 1952 3929 2048
rect 3934 2002 3937 2068
rect 3950 2052 3953 2058
rect 3966 2022 3969 2048
rect 3950 1968 3966 1971
rect 3890 1948 3894 1951
rect 3822 1942 3825 1948
rect 3838 1942 3841 1948
rect 3846 1942 3849 1948
rect 3798 1902 3801 1938
rect 3838 1931 3841 1938
rect 3838 1928 3849 1931
rect 3830 1892 3833 1898
rect 3846 1892 3849 1928
rect 3854 1902 3857 1948
rect 3878 1942 3881 1948
rect 3902 1942 3905 1948
rect 3918 1942 3921 1948
rect 3934 1942 3937 1958
rect 3950 1932 3953 1968
rect 3982 1962 3985 2138
rect 3990 2102 3993 2128
rect 3998 2082 4001 2118
rect 4006 2102 4009 2148
rect 4030 2142 4033 2148
rect 4038 2082 4041 2158
rect 4046 2152 4049 2158
rect 4054 2152 4057 2178
rect 4062 2152 4065 2168
rect 4094 2162 4097 2198
rect 4126 2162 4129 2218
rect 4134 2212 4137 2218
rect 4134 2172 4137 2178
rect 4142 2172 4145 2178
rect 4082 2148 4086 2151
rect 4110 2142 4113 2148
rect 4118 2142 4121 2148
rect 4054 2132 4057 2138
rect 4062 2092 4065 2118
rect 4070 2102 4073 2138
rect 4080 2103 4082 2107
rect 4086 2103 4089 2107
rect 4093 2103 4096 2107
rect 4070 2082 4073 2098
rect 4126 2081 4129 2138
rect 4134 2122 4137 2148
rect 4158 2092 4161 2148
rect 4166 2142 4169 2218
rect 4182 2182 4185 2318
rect 4190 2262 4193 2318
rect 4198 2262 4201 2318
rect 4206 2312 4209 2358
rect 4226 2348 4230 2351
rect 4274 2348 4278 2351
rect 4214 2292 4217 2348
rect 4246 2332 4249 2338
rect 4262 2332 4265 2338
rect 4266 2328 4273 2331
rect 4246 2282 4249 2308
rect 4254 2271 4257 2318
rect 4270 2282 4273 2328
rect 4294 2292 4297 2348
rect 4314 2328 4318 2331
rect 4326 2312 4329 2368
rect 4342 2362 4345 2368
rect 4362 2358 4366 2361
rect 4438 2361 4441 2408
rect 4478 2402 4481 2448
rect 4490 2428 4494 2431
rect 4566 2422 4569 2428
rect 4518 2372 4521 2378
rect 4502 2362 4505 2368
rect 4434 2358 4441 2361
rect 4466 2358 4470 2361
rect 4334 2352 4337 2358
rect 4362 2348 4366 2351
rect 4354 2338 4361 2341
rect 4302 2292 4305 2308
rect 4250 2268 4257 2271
rect 4262 2272 4265 2278
rect 4266 2258 4270 2261
rect 4190 2232 4193 2248
rect 4198 2242 4201 2258
rect 4258 2248 4262 2251
rect 4210 2238 4214 2241
rect 4222 2232 4225 2238
rect 4286 2232 4289 2268
rect 4302 2262 4305 2278
rect 4346 2268 4350 2271
rect 4326 2262 4329 2268
rect 4314 2258 4318 2261
rect 4294 2212 4297 2258
rect 4302 2192 4305 2258
rect 4334 2252 4337 2268
rect 4346 2248 4350 2251
rect 4326 2192 4329 2238
rect 4342 2222 4345 2228
rect 4350 2192 4353 2208
rect 4254 2172 4257 2178
rect 4286 2162 4289 2178
rect 4182 2152 4185 2158
rect 4230 2152 4233 2158
rect 4202 2148 4206 2151
rect 4258 2148 4262 2151
rect 4290 2148 4294 2151
rect 4306 2148 4310 2151
rect 4214 2142 4217 2148
rect 4318 2142 4321 2148
rect 4178 2138 4182 2141
rect 4282 2138 4286 2141
rect 4198 2132 4201 2138
rect 4178 2128 4182 2131
rect 4122 2078 4129 2081
rect 4166 2082 4169 2128
rect 4014 2072 4017 2078
rect 4146 2068 4150 2071
rect 3998 2012 4001 2068
rect 4046 2062 4049 2068
rect 4018 2058 4022 2061
rect 4030 2042 4033 2048
rect 4018 2038 4022 2041
rect 3966 1952 3969 1958
rect 3958 1942 3961 1948
rect 3958 1932 3961 1938
rect 3918 1902 3921 1928
rect 3870 1882 3873 1898
rect 3918 1892 3921 1898
rect 3922 1878 3926 1881
rect 3838 1872 3841 1878
rect 3862 1872 3865 1878
rect 3886 1872 3889 1878
rect 3810 1868 3814 1871
rect 3926 1862 3929 1878
rect 3934 1872 3937 1928
rect 3982 1921 3985 1958
rect 4002 1948 4006 1951
rect 3990 1932 3993 1938
rect 3982 1918 3993 1921
rect 3942 1882 3945 1918
rect 3958 1892 3961 1908
rect 3966 1862 3969 1878
rect 3974 1872 3977 1898
rect 3982 1892 3985 1908
rect 3802 1858 3806 1861
rect 3822 1832 3825 1858
rect 3942 1852 3945 1858
rect 3890 1848 3894 1851
rect 3766 1802 3769 1818
rect 3806 1812 3809 1818
rect 3766 1762 3769 1798
rect 3782 1762 3785 1808
rect 3754 1758 3758 1761
rect 3794 1748 3798 1751
rect 3806 1742 3809 1788
rect 3706 1678 3710 1681
rect 3678 1668 3686 1671
rect 3682 1658 3686 1661
rect 3670 1652 3673 1658
rect 3678 1642 3681 1648
rect 3698 1638 3702 1641
rect 3686 1552 3689 1618
rect 3710 1592 3713 1668
rect 3718 1662 3721 1718
rect 3726 1712 3729 1738
rect 3758 1732 3761 1740
rect 3770 1718 3774 1721
rect 3742 1662 3745 1708
rect 3766 1682 3769 1698
rect 3782 1682 3785 1718
rect 3814 1702 3817 1758
rect 3838 1752 3841 1838
rect 3846 1832 3849 1848
rect 3854 1812 3857 1818
rect 3830 1742 3833 1748
rect 3782 1662 3785 1668
rect 3806 1662 3809 1678
rect 3722 1648 3726 1651
rect 3742 1622 3745 1628
rect 3718 1582 3721 1618
rect 3774 1552 3777 1658
rect 3610 1548 3614 1551
rect 3650 1548 3654 1551
rect 3786 1548 3790 1551
rect 3514 1538 3529 1541
rect 3514 1468 3518 1471
rect 3526 1461 3529 1538
rect 3542 1472 3545 1548
rect 3622 1542 3625 1548
rect 3562 1538 3566 1541
rect 3634 1538 3638 1541
rect 3706 1538 3710 1541
rect 3550 1532 3553 1538
rect 3566 1482 3569 1538
rect 3566 1472 3569 1478
rect 3526 1458 3534 1461
rect 3514 1448 3518 1451
rect 3470 1392 3473 1398
rect 3470 1382 3473 1388
rect 3486 1292 3489 1448
rect 3494 1352 3497 1438
rect 3506 1388 3510 1391
rect 3490 1268 3494 1271
rect 3502 1262 3505 1358
rect 3526 1352 3529 1458
rect 3582 1452 3585 1458
rect 3554 1418 3558 1421
rect 3534 1362 3537 1418
rect 3568 1403 3570 1407
rect 3574 1403 3577 1407
rect 3581 1403 3584 1407
rect 3590 1382 3593 1468
rect 3566 1362 3569 1378
rect 3598 1362 3601 1518
rect 3646 1492 3649 1528
rect 3662 1492 3665 1538
rect 3670 1522 3673 1528
rect 3674 1478 3678 1481
rect 3614 1472 3617 1478
rect 3702 1472 3705 1488
rect 3614 1452 3617 1458
rect 3614 1362 3617 1418
rect 3514 1348 3518 1351
rect 3526 1342 3529 1348
rect 3534 1312 3537 1348
rect 3558 1342 3561 1348
rect 3542 1332 3545 1338
rect 3558 1322 3561 1328
rect 3530 1268 3534 1271
rect 3538 1258 3542 1261
rect 3470 1252 3473 1258
rect 3482 1248 3486 1251
rect 3502 1251 3505 1258
rect 3502 1248 3510 1251
rect 3526 1251 3529 1258
rect 3550 1252 3553 1318
rect 3526 1248 3537 1251
rect 3534 1232 3537 1248
rect 3482 1188 3489 1191
rect 3438 1152 3441 1168
rect 3454 1152 3457 1158
rect 3462 1152 3465 1188
rect 3470 1152 3473 1168
rect 3314 1078 3318 1081
rect 3418 1078 3422 1081
rect 3350 1072 3353 1078
rect 3358 1070 3361 1078
rect 3398 1072 3401 1078
rect 3438 1072 3441 1148
rect 3470 1142 3473 1148
rect 3450 1138 3454 1141
rect 3478 1132 3481 1138
rect 3486 1132 3489 1188
rect 3502 1172 3505 1218
rect 3502 1152 3505 1168
rect 3534 1162 3537 1228
rect 3522 1158 3526 1161
rect 3514 1148 3518 1151
rect 3510 1142 3513 1148
rect 3534 1142 3537 1158
rect 3502 1132 3505 1138
rect 3538 1128 3542 1131
rect 3450 1078 3454 1081
rect 3310 1062 3313 1068
rect 3334 1062 3337 1068
rect 3338 1048 3342 1051
rect 3322 1018 3326 1021
rect 3334 981 3337 1038
rect 3350 1022 3353 1068
rect 3386 1068 3390 1071
rect 3486 1062 3489 1068
rect 3386 1058 3390 1061
rect 3406 1052 3409 1058
rect 3330 978 3337 981
rect 3342 982 3345 988
rect 3318 962 3321 968
rect 3326 942 3329 958
rect 3350 952 3353 958
rect 3358 942 3361 948
rect 3374 942 3377 988
rect 3382 952 3385 1048
rect 3426 1038 3430 1041
rect 3438 982 3441 1058
rect 3450 1048 3454 1051
rect 3398 972 3401 978
rect 3454 962 3457 1018
rect 3470 1012 3473 1018
rect 3486 992 3489 1058
rect 3494 1042 3497 1118
rect 3506 1078 3510 1081
rect 3506 1058 3510 1061
rect 3518 1042 3521 1048
rect 3494 1002 3497 1018
rect 3526 1012 3529 1078
rect 3534 1062 3537 1098
rect 3550 1092 3553 1158
rect 3558 1082 3561 1318
rect 3566 1272 3569 1358
rect 3606 1322 3609 1338
rect 3614 1332 3617 1348
rect 3590 1262 3593 1308
rect 3606 1282 3609 1298
rect 3602 1268 3606 1271
rect 3570 1248 3574 1251
rect 3614 1251 3617 1318
rect 3622 1302 3625 1468
rect 3630 1462 3633 1468
rect 3654 1462 3657 1468
rect 3710 1462 3713 1478
rect 3718 1472 3721 1478
rect 3726 1472 3729 1538
rect 3734 1472 3737 1540
rect 3750 1492 3753 1518
rect 3766 1502 3769 1518
rect 3774 1492 3777 1548
rect 3790 1512 3793 1538
rect 3674 1458 3678 1461
rect 3698 1458 3702 1461
rect 3670 1361 3673 1438
rect 3678 1382 3681 1448
rect 3726 1392 3729 1458
rect 3710 1362 3713 1378
rect 3670 1358 3678 1361
rect 3726 1352 3729 1368
rect 3734 1352 3737 1458
rect 3742 1452 3745 1458
rect 3750 1361 3753 1428
rect 3758 1372 3761 1418
rect 3750 1358 3758 1361
rect 3634 1348 3638 1351
rect 3666 1338 3670 1341
rect 3630 1312 3633 1338
rect 3702 1332 3705 1348
rect 3766 1342 3769 1488
rect 3798 1482 3801 1518
rect 3806 1512 3809 1538
rect 3786 1468 3790 1471
rect 3774 1462 3777 1468
rect 3798 1462 3801 1468
rect 3806 1462 3809 1508
rect 3814 1462 3817 1668
rect 3822 1652 3825 1718
rect 3830 1631 3833 1708
rect 3838 1662 3841 1738
rect 3846 1722 3849 1808
rect 3878 1802 3881 1818
rect 3862 1762 3865 1798
rect 3866 1748 3870 1751
rect 3886 1742 3889 1788
rect 3902 1772 3905 1848
rect 3990 1841 3993 1918
rect 3998 1862 4001 1918
rect 4014 1912 4017 1958
rect 4022 1932 4025 1938
rect 4038 1902 4041 2058
rect 4046 1942 4049 1958
rect 4054 1952 4057 1988
rect 4078 1962 4081 2018
rect 4094 1992 4097 2038
rect 4110 2022 4113 2068
rect 4126 2032 4129 2068
rect 4166 2062 4169 2068
rect 4190 2062 4193 2098
rect 4062 1942 4065 1948
rect 4082 1938 4086 1941
rect 4102 1932 4105 1998
rect 4118 1942 4121 1948
rect 4126 1932 4129 2028
rect 4142 1952 4145 2048
rect 4150 1972 4153 2058
rect 4198 2052 4201 2128
rect 4206 2082 4209 2138
rect 4262 2122 4265 2138
rect 4270 2132 4273 2138
rect 4222 2082 4225 2098
rect 4254 2092 4257 2108
rect 4294 2092 4297 2118
rect 4310 2112 4313 2138
rect 4326 2132 4329 2148
rect 4194 2048 4198 2051
rect 4182 2042 4185 2048
rect 4206 2032 4209 2058
rect 4234 2048 4238 2051
rect 4182 1992 4185 2018
rect 4190 1992 4193 2018
rect 4206 1982 4209 2028
rect 4254 1992 4257 2078
rect 4262 2062 4265 2088
rect 4310 2082 4313 2108
rect 4334 2092 4337 2188
rect 4358 2172 4361 2338
rect 4374 2312 4377 2358
rect 4406 2352 4409 2358
rect 4426 2348 4430 2351
rect 4514 2348 4518 2351
rect 4410 2338 4414 2341
rect 4382 2322 4385 2328
rect 4398 2322 4401 2338
rect 4494 2332 4497 2348
rect 4526 2342 4529 2388
rect 4542 2372 4545 2378
rect 4542 2352 4545 2358
rect 4518 2338 4526 2341
rect 4426 2328 4430 2331
rect 4458 2328 4462 2331
rect 4466 2318 4470 2321
rect 4390 2292 4393 2318
rect 4378 2278 4382 2281
rect 4374 2182 4377 2278
rect 4390 2252 4393 2258
rect 4342 2162 4345 2168
rect 4382 2142 4385 2148
rect 4350 2132 4353 2138
rect 4390 2121 4393 2138
rect 4398 2132 4401 2278
rect 4446 2272 4449 2318
rect 4470 2282 4473 2288
rect 4478 2272 4481 2328
rect 4494 2321 4497 2328
rect 4486 2318 4497 2321
rect 4458 2268 4462 2271
rect 4406 2262 4409 2268
rect 4442 2258 4446 2261
rect 4414 2251 4417 2258
rect 4406 2248 4417 2251
rect 4406 2192 4409 2248
rect 4430 2172 4433 2208
rect 4426 2168 4430 2171
rect 4438 2152 4441 2218
rect 4454 2202 4457 2258
rect 4478 2212 4481 2268
rect 4486 2242 4489 2318
rect 4494 2292 4497 2298
rect 4498 2258 4502 2261
rect 4502 2242 4505 2248
rect 4494 2232 4497 2238
rect 4478 2192 4481 2198
rect 4510 2162 4513 2238
rect 4518 2192 4521 2338
rect 4534 2332 4537 2338
rect 4542 2322 4545 2348
rect 4574 2342 4577 2468
rect 4590 2412 4593 2418
rect 4582 2352 4585 2358
rect 4562 2328 4566 2331
rect 4526 2252 4529 2258
rect 4538 2238 4542 2241
rect 4526 2232 4529 2238
rect 4434 2148 4438 2151
rect 4454 2142 4457 2148
rect 4434 2138 4438 2141
rect 4402 2128 4406 2131
rect 4422 2128 4430 2131
rect 4390 2118 4401 2121
rect 4398 2092 4401 2118
rect 4414 2092 4417 2128
rect 4422 2082 4425 2128
rect 4462 2122 4465 2158
rect 4474 2148 4478 2151
rect 4498 2148 4502 2151
rect 4438 2092 4441 2118
rect 4430 2082 4433 2088
rect 4370 2078 4374 2081
rect 4270 2072 4273 2078
rect 4278 2022 4281 2058
rect 4290 2048 4294 2051
rect 4302 2022 4305 2078
rect 4342 2072 4345 2078
rect 4358 2072 4361 2078
rect 4190 1962 4193 1968
rect 4162 1958 4166 1961
rect 4246 1952 4249 1968
rect 4294 1962 4297 1968
rect 4138 1948 4142 1951
rect 4194 1948 4198 1951
rect 4226 1948 4230 1951
rect 4150 1932 4153 1938
rect 4166 1932 4169 1938
rect 4074 1928 4078 1931
rect 4046 1922 4049 1928
rect 4054 1892 4057 1928
rect 4080 1903 4082 1907
rect 4086 1903 4089 1907
rect 4093 1903 4096 1907
rect 4142 1892 4145 1918
rect 4018 1878 4022 1881
rect 4082 1878 4086 1881
rect 4006 1871 4009 1878
rect 4046 1872 4049 1878
rect 4006 1868 4014 1871
rect 4098 1858 4102 1861
rect 3998 1852 4001 1858
rect 4038 1852 4041 1858
rect 4018 1848 4022 1851
rect 4110 1842 4113 1848
rect 3990 1838 4001 1841
rect 3910 1752 3913 1758
rect 3918 1752 3921 1758
rect 3934 1752 3937 1808
rect 3998 1802 4001 1838
rect 4030 1812 4033 1838
rect 3942 1742 3945 1778
rect 3966 1742 3969 1788
rect 3974 1752 3977 1798
rect 3998 1792 4001 1798
rect 4030 1792 4033 1808
rect 4054 1772 4057 1818
rect 4094 1762 4097 1788
rect 4110 1752 4113 1818
rect 4010 1748 4014 1751
rect 3982 1742 3985 1748
rect 4118 1742 4121 1878
rect 4134 1872 4137 1878
rect 4130 1858 4134 1861
rect 4138 1748 4142 1751
rect 3854 1732 3857 1738
rect 3846 1672 3849 1718
rect 3862 1681 3865 1738
rect 3858 1678 3865 1681
rect 3870 1672 3873 1738
rect 3878 1732 3881 1738
rect 3926 1732 3929 1738
rect 4046 1732 4049 1738
rect 3946 1728 3950 1731
rect 3878 1702 3881 1728
rect 3902 1672 3905 1678
rect 3874 1658 3878 1661
rect 3890 1658 3894 1661
rect 3902 1651 3905 1658
rect 3898 1648 3905 1651
rect 3838 1642 3841 1648
rect 3854 1642 3857 1648
rect 3830 1628 3841 1631
rect 3774 1422 3777 1448
rect 3806 1431 3809 1458
rect 3822 1452 3825 1518
rect 3830 1492 3833 1528
rect 3838 1492 3841 1628
rect 3854 1552 3857 1638
rect 3894 1562 3897 1568
rect 3866 1538 3870 1541
rect 3846 1472 3849 1538
rect 3862 1502 3865 1518
rect 3878 1492 3881 1538
rect 3798 1428 3809 1431
rect 3782 1402 3785 1418
rect 3782 1362 3785 1368
rect 3746 1338 3750 1341
rect 3798 1341 3801 1428
rect 3810 1418 3814 1421
rect 3814 1392 3817 1408
rect 3838 1352 3841 1358
rect 3846 1352 3849 1468
rect 3862 1382 3865 1458
rect 3870 1452 3873 1468
rect 3878 1352 3881 1358
rect 3866 1348 3870 1351
rect 3830 1342 3833 1348
rect 3798 1338 3806 1341
rect 3642 1318 3646 1321
rect 3630 1291 3633 1308
rect 3622 1288 3633 1291
rect 3622 1262 3625 1288
rect 3630 1272 3633 1278
rect 3654 1272 3657 1328
rect 3678 1302 3681 1318
rect 3686 1312 3689 1328
rect 3694 1322 3697 1328
rect 3686 1292 3689 1308
rect 3702 1292 3705 1308
rect 3718 1292 3721 1318
rect 3734 1292 3737 1338
rect 3662 1272 3665 1288
rect 3670 1272 3673 1288
rect 3718 1262 3721 1288
rect 3626 1258 3633 1261
rect 3642 1258 3646 1261
rect 3674 1258 3678 1261
rect 3610 1248 3617 1251
rect 3622 1222 3625 1228
rect 3568 1203 3570 1207
rect 3574 1203 3577 1207
rect 3581 1203 3584 1207
rect 3582 1162 3585 1168
rect 3570 1158 3577 1161
rect 3574 1151 3577 1158
rect 3574 1148 3585 1151
rect 3566 1142 3569 1148
rect 3566 1102 3569 1138
rect 3574 1132 3577 1138
rect 3582 1122 3585 1148
rect 3590 1082 3593 1158
rect 3622 1132 3625 1208
rect 3630 1142 3633 1258
rect 3654 1212 3657 1258
rect 3694 1252 3697 1258
rect 3734 1252 3737 1268
rect 3678 1212 3681 1218
rect 3654 1192 3657 1198
rect 3678 1162 3681 1188
rect 3690 1158 3694 1161
rect 3646 1142 3649 1148
rect 3618 1128 3622 1131
rect 3630 1112 3633 1128
rect 3670 1122 3673 1158
rect 3726 1142 3729 1218
rect 3734 1192 3737 1248
rect 3742 1222 3745 1278
rect 3750 1212 3753 1318
rect 3758 1292 3761 1328
rect 3758 1262 3761 1268
rect 3758 1252 3761 1258
rect 3738 1148 3742 1151
rect 3690 1138 3694 1141
rect 3714 1138 3718 1141
rect 3750 1141 3753 1158
rect 3766 1152 3769 1338
rect 3774 1282 3777 1338
rect 3786 1328 3790 1331
rect 3798 1322 3801 1338
rect 3830 1322 3833 1338
rect 3782 1302 3785 1318
rect 3798 1312 3801 1318
rect 3774 1272 3777 1278
rect 3782 1262 3785 1288
rect 3798 1282 3801 1308
rect 3846 1302 3849 1348
rect 3854 1342 3857 1348
rect 3842 1288 3846 1291
rect 3822 1272 3825 1278
rect 3870 1272 3873 1298
rect 3742 1138 3753 1141
rect 3758 1142 3761 1148
rect 3678 1132 3681 1138
rect 3618 1078 3622 1081
rect 3542 1062 3545 1068
rect 3558 1002 3561 1078
rect 3570 1068 3574 1071
rect 3582 1052 3585 1058
rect 3568 1003 3570 1007
rect 3574 1003 3577 1007
rect 3581 1003 3584 1007
rect 3402 948 3406 951
rect 3346 938 3350 941
rect 3414 941 3417 958
rect 3526 952 3529 998
rect 3542 952 3545 958
rect 3558 952 3561 968
rect 3590 962 3593 1058
rect 3426 948 3430 951
rect 3458 948 3470 951
rect 3518 942 3521 948
rect 3406 938 3417 941
rect 3258 888 3262 891
rect 3270 872 3273 898
rect 3290 888 3294 891
rect 3302 882 3305 938
rect 3390 932 3393 938
rect 3298 868 3302 871
rect 3310 862 3313 898
rect 3214 858 3222 861
rect 3274 858 3278 861
rect 3290 848 3294 851
rect 3206 842 3209 848
rect 3226 838 3230 841
rect 3014 832 3017 838
rect 2934 762 2937 768
rect 2962 758 2966 761
rect 2930 748 2934 751
rect 2974 742 2977 788
rect 2990 762 2993 788
rect 2990 742 2993 748
rect 2938 738 2942 741
rect 2910 712 2913 718
rect 2906 688 2910 691
rect 2870 678 2881 681
rect 2878 672 2881 678
rect 2942 672 2945 738
rect 2930 668 2934 671
rect 2870 662 2873 668
rect 2886 662 2889 668
rect 2870 592 2873 618
rect 2902 572 2905 648
rect 2910 612 2913 668
rect 2950 662 2953 738
rect 3006 732 3009 818
rect 3014 742 3017 778
rect 3022 752 3025 818
rect 3054 752 3057 778
rect 2994 728 2998 731
rect 2922 658 2926 661
rect 2914 608 2921 611
rect 2910 562 2913 598
rect 2918 562 2921 608
rect 2874 548 2878 551
rect 2850 538 2854 541
rect 2866 538 2870 541
rect 2898 538 2902 541
rect 2926 541 2929 658
rect 2966 652 2969 718
rect 2982 692 2985 698
rect 2990 681 2993 718
rect 3022 692 3025 738
rect 3030 732 3033 738
rect 3038 692 3041 748
rect 3062 742 3065 828
rect 3090 788 3094 791
rect 3134 762 3137 818
rect 3106 758 3110 761
rect 3106 748 3113 751
rect 3098 738 3102 741
rect 3058 728 3062 731
rect 3048 703 3050 707
rect 3054 703 3057 707
rect 3061 703 3064 707
rect 3030 682 3033 688
rect 2982 678 2993 681
rect 2974 672 2977 678
rect 2934 642 2937 648
rect 2942 592 2945 618
rect 2950 612 2953 618
rect 2966 552 2969 558
rect 2958 542 2961 548
rect 2926 538 2934 541
rect 2810 488 2814 491
rect 2866 488 2870 491
rect 2626 448 2630 451
rect 2330 358 2334 361
rect 2394 358 2398 361
rect 2450 358 2457 361
rect 2350 352 2353 358
rect 2306 348 2310 351
rect 2386 348 2390 351
rect 2442 348 2446 351
rect 2286 328 2297 331
rect 2386 338 2390 341
rect 2286 292 2289 328
rect 2298 288 2302 291
rect 2294 262 2297 278
rect 2234 248 2238 251
rect 2126 152 2129 178
rect 2166 162 2169 178
rect 2210 158 2214 161
rect 2150 152 2153 158
rect 2162 148 2166 151
rect 2202 148 2206 151
rect 2150 132 2153 148
rect 2182 142 2185 148
rect 2014 58 2022 61
rect 2082 58 2086 61
rect 1910 52 1913 58
rect 2014 52 2017 58
rect 2070 52 2073 58
rect 1862 48 1870 51
rect 2002 48 2006 51
rect 2102 42 2105 68
rect 2118 62 2121 78
rect 2134 72 2137 98
rect 2142 62 2145 118
rect 2174 92 2177 138
rect 2158 82 2161 88
rect 2182 72 2185 78
rect 2114 58 2118 61
rect 2130 58 2134 61
rect 2154 58 2158 61
rect 2142 52 2145 58
rect 2190 52 2193 78
rect 2198 62 2201 148
rect 2226 128 2230 131
rect 2206 92 2209 118
rect 2214 72 2217 88
rect 2222 72 2225 108
rect 2238 92 2241 148
rect 2246 142 2249 208
rect 2254 152 2257 238
rect 2262 232 2265 248
rect 2270 191 2273 258
rect 2266 188 2273 191
rect 2262 142 2265 188
rect 2274 158 2278 161
rect 2270 92 2273 98
rect 2286 62 2289 198
rect 2294 192 2297 258
rect 2310 232 2313 338
rect 2318 312 2321 338
rect 2326 322 2329 328
rect 2358 302 2361 338
rect 2366 322 2369 328
rect 2406 322 2409 338
rect 2414 332 2417 338
rect 2326 272 2329 288
rect 2358 282 2361 298
rect 2346 278 2350 281
rect 2326 262 2329 268
rect 2318 232 2321 258
rect 2334 232 2337 278
rect 2346 258 2350 261
rect 2350 192 2353 248
rect 2358 212 2361 268
rect 2358 182 2361 188
rect 2366 172 2369 258
rect 2350 152 2353 158
rect 2374 152 2377 308
rect 2386 288 2390 291
rect 2390 272 2393 278
rect 2382 252 2385 258
rect 2390 252 2393 268
rect 2406 262 2409 318
rect 2414 282 2417 288
rect 2446 272 2449 318
rect 2454 292 2457 358
rect 2462 342 2465 348
rect 2470 342 2473 348
rect 2478 342 2481 408
rect 2506 358 2510 361
rect 2490 348 2494 351
rect 2526 342 2529 418
rect 2544 403 2546 407
rect 2550 403 2553 407
rect 2557 403 2560 407
rect 2558 342 2561 378
rect 2590 362 2593 378
rect 2586 348 2590 351
rect 2574 342 2577 348
rect 2486 282 2489 328
rect 2418 268 2422 271
rect 2454 262 2457 268
rect 2418 258 2422 261
rect 2442 258 2446 261
rect 2398 192 2401 258
rect 2450 248 2454 251
rect 2438 192 2441 208
rect 2462 202 2465 278
rect 2486 272 2489 278
rect 2494 262 2497 288
rect 2502 261 2505 318
rect 2510 292 2513 318
rect 2534 292 2537 338
rect 2538 278 2542 281
rect 2574 271 2577 318
rect 2598 272 2601 338
rect 2606 311 2609 418
rect 2622 392 2625 428
rect 2646 392 2649 408
rect 2618 348 2622 351
rect 2630 342 2633 378
rect 2654 372 2657 418
rect 2662 382 2665 438
rect 2702 422 2705 478
rect 2710 472 2713 488
rect 2778 478 2782 481
rect 2718 472 2721 478
rect 2758 472 2761 478
rect 2822 472 2825 478
rect 2846 472 2849 478
rect 2886 472 2889 518
rect 2902 492 2905 528
rect 2894 482 2897 488
rect 2778 468 2782 471
rect 2842 468 2846 471
rect 2906 468 2910 471
rect 2830 462 2833 468
rect 2862 462 2865 468
rect 2918 462 2921 478
rect 2762 458 2766 461
rect 2810 458 2817 461
rect 2718 452 2721 458
rect 2802 448 2806 451
rect 2730 438 2734 441
rect 2654 352 2657 368
rect 2662 362 2665 378
rect 2662 342 2665 348
rect 2678 342 2681 398
rect 2710 362 2713 368
rect 2690 348 2694 351
rect 2706 348 2710 351
rect 2734 351 2737 368
rect 2742 362 2745 448
rect 2750 412 2753 448
rect 2766 392 2769 418
rect 2806 392 2809 428
rect 2814 392 2817 458
rect 2830 442 2833 448
rect 2878 442 2881 458
rect 2886 392 2889 458
rect 2926 452 2929 518
rect 2934 472 2937 538
rect 2942 522 2945 528
rect 2974 522 2977 668
rect 2982 572 2985 678
rect 3006 672 3009 678
rect 3058 668 3062 671
rect 2990 622 2993 668
rect 3014 662 3017 668
rect 3070 662 3073 738
rect 3110 732 3113 748
rect 3094 692 3097 708
rect 3078 672 3081 678
rect 3002 658 3006 661
rect 3042 648 3046 651
rect 2990 582 2993 588
rect 2982 532 2985 548
rect 2942 462 2945 498
rect 2990 492 2993 568
rect 2950 472 2953 478
rect 2978 468 2982 471
rect 2970 458 2974 461
rect 2734 348 2742 351
rect 2690 338 2694 341
rect 2738 338 2742 341
rect 2630 312 2633 338
rect 2638 332 2641 338
rect 2726 332 2729 338
rect 2718 322 2721 328
rect 2606 308 2614 311
rect 2606 292 2609 298
rect 2662 282 2665 288
rect 2630 272 2633 278
rect 2574 268 2582 271
rect 2642 268 2646 271
rect 2502 258 2510 261
rect 2470 192 2473 258
rect 2478 182 2481 258
rect 2506 248 2510 251
rect 2526 242 2529 268
rect 2510 192 2513 228
rect 2534 192 2537 268
rect 2566 252 2569 268
rect 2610 258 2614 261
rect 2618 258 2622 261
rect 2598 252 2601 258
rect 2606 241 2609 248
rect 2598 238 2609 241
rect 2578 228 2582 231
rect 2544 203 2546 207
rect 2550 203 2553 207
rect 2557 203 2560 207
rect 2598 192 2601 238
rect 2574 162 2577 168
rect 2418 158 2422 161
rect 2382 152 2385 158
rect 2314 148 2318 151
rect 2314 138 2318 141
rect 2294 132 2297 138
rect 2330 128 2334 131
rect 2294 92 2297 128
rect 2358 121 2361 148
rect 2398 142 2401 148
rect 2426 138 2430 141
rect 2370 128 2374 131
rect 2382 121 2385 138
rect 2358 118 2369 121
rect 2354 78 2358 81
rect 2366 72 2369 118
rect 2374 118 2385 121
rect 2374 92 2377 118
rect 2406 112 2409 138
rect 2414 82 2417 138
rect 2438 132 2441 148
rect 2422 112 2425 118
rect 2454 112 2457 158
rect 2466 148 2470 151
rect 2538 148 2542 151
rect 2546 148 2550 151
rect 2470 132 2473 138
rect 2486 122 2489 138
rect 2494 112 2497 148
rect 2518 122 2521 138
rect 2558 122 2561 158
rect 2590 142 2593 188
rect 2622 152 2625 248
rect 2638 242 2641 258
rect 2662 252 2665 258
rect 2678 251 2681 308
rect 2698 268 2702 271
rect 2686 262 2689 268
rect 2710 262 2713 308
rect 2726 292 2729 318
rect 2750 292 2753 358
rect 2766 352 2769 378
rect 2782 352 2785 358
rect 2814 352 2817 358
rect 2830 352 2833 358
rect 2814 342 2817 348
rect 2822 342 2825 348
rect 2794 338 2798 341
rect 2770 288 2774 291
rect 2754 278 2758 281
rect 2774 272 2777 278
rect 2782 272 2785 338
rect 2806 322 2809 328
rect 2838 322 2841 328
rect 2738 268 2742 271
rect 2782 262 2785 268
rect 2790 262 2793 318
rect 2814 292 2817 308
rect 2846 292 2849 358
rect 2862 352 2865 358
rect 2910 352 2913 358
rect 2882 348 2886 351
rect 2854 342 2857 348
rect 2882 338 2886 341
rect 2870 272 2873 338
rect 2858 268 2862 271
rect 2890 268 2894 271
rect 2874 258 2878 261
rect 2890 258 2894 261
rect 2678 248 2686 251
rect 2710 242 2713 258
rect 2722 248 2726 251
rect 2746 248 2750 251
rect 2674 238 2678 241
rect 2686 232 2689 238
rect 2638 192 2641 198
rect 2630 152 2633 188
rect 2662 182 2665 218
rect 2674 188 2678 191
rect 2662 152 2665 178
rect 2686 152 2689 158
rect 2694 152 2697 158
rect 2702 152 2705 158
rect 2734 152 2737 168
rect 2742 161 2745 218
rect 2770 168 2774 171
rect 2758 162 2761 168
rect 2742 158 2750 161
rect 2722 148 2726 151
rect 2754 148 2758 151
rect 2770 148 2774 151
rect 2614 142 2617 148
rect 2782 142 2785 258
rect 2790 162 2793 258
rect 2798 222 2801 258
rect 2822 252 2825 258
rect 2838 252 2841 258
rect 2902 252 2905 258
rect 2882 248 2886 251
rect 2798 192 2801 198
rect 2838 192 2841 238
rect 2862 202 2865 248
rect 2910 242 2913 348
rect 2918 292 2921 408
rect 2934 352 2937 458
rect 2950 448 2958 451
rect 2986 448 2990 451
rect 2942 392 2945 438
rect 2934 282 2937 338
rect 2950 292 2953 448
rect 2974 442 2977 448
rect 2998 441 3001 578
rect 3006 562 3009 568
rect 3014 492 3017 588
rect 3022 572 3025 598
rect 3030 592 3033 648
rect 3042 558 3046 561
rect 3022 542 3025 558
rect 3042 548 3046 551
rect 3070 542 3073 658
rect 3078 642 3081 668
rect 3102 662 3105 668
rect 3118 661 3121 758
rect 3130 738 3134 741
rect 3142 712 3145 758
rect 3158 741 3161 838
rect 3166 762 3169 808
rect 3238 792 3241 798
rect 3254 792 3257 808
rect 3178 758 3182 761
rect 3190 752 3193 758
rect 3154 738 3161 741
rect 3186 738 3190 741
rect 3142 682 3145 688
rect 3114 658 3121 661
rect 3134 662 3137 668
rect 3034 538 3038 541
rect 3048 503 3050 507
rect 3054 503 3057 507
rect 3061 503 3064 507
rect 3078 492 3081 598
rect 3094 582 3097 648
rect 3126 642 3129 648
rect 3142 602 3145 658
rect 3142 592 3145 598
rect 3126 562 3129 578
rect 3098 558 3102 561
rect 3114 548 3118 551
rect 3098 538 3102 541
rect 3122 538 3126 541
rect 3066 478 3070 481
rect 3030 472 3033 478
rect 3010 468 3014 471
rect 2990 438 3001 441
rect 2934 262 2937 278
rect 2958 272 2961 358
rect 2966 332 2969 428
rect 2990 392 2993 438
rect 3014 432 3017 448
rect 3030 392 3033 458
rect 3038 452 3041 478
rect 3094 472 3097 538
rect 3110 472 3113 528
rect 3150 492 3153 728
rect 3158 702 3161 718
rect 3174 692 3177 728
rect 3158 662 3161 688
rect 3166 672 3169 678
rect 3182 662 3185 718
rect 3198 692 3201 758
rect 3206 732 3209 748
rect 3214 741 3217 788
rect 3222 752 3225 758
rect 3214 738 3222 741
rect 3214 672 3217 698
rect 3222 672 3225 728
rect 3230 702 3233 758
rect 3238 721 3241 768
rect 3262 752 3265 848
rect 3270 742 3273 798
rect 3294 762 3297 768
rect 3310 761 3313 858
rect 3318 772 3321 918
rect 3334 892 3337 918
rect 3326 852 3329 868
rect 3310 758 3321 761
rect 3302 752 3305 758
rect 3278 742 3281 748
rect 3310 741 3313 748
rect 3302 738 3313 741
rect 3318 742 3321 758
rect 3342 752 3345 898
rect 3406 892 3409 938
rect 3422 932 3425 938
rect 3478 932 3481 938
rect 3486 932 3489 938
rect 3494 932 3497 938
rect 3458 928 3462 931
rect 3526 931 3529 948
rect 3534 942 3537 948
rect 3558 942 3561 948
rect 3598 942 3601 1078
rect 3638 1072 3641 1078
rect 3610 1068 3614 1071
rect 3662 1062 3665 1108
rect 3686 1092 3689 1128
rect 3694 1102 3697 1138
rect 3742 1132 3745 1138
rect 3750 1122 3753 1128
rect 3706 1118 3710 1121
rect 3674 1068 3678 1071
rect 3698 1068 3702 1071
rect 3650 1058 3654 1061
rect 3698 1058 3702 1061
rect 3674 1048 3678 1051
rect 3702 1042 3705 1048
rect 3646 972 3649 1018
rect 3662 992 3665 998
rect 3678 962 3681 968
rect 3702 962 3705 968
rect 3626 958 3630 961
rect 3642 958 3646 961
rect 3626 948 3630 951
rect 3666 948 3670 951
rect 3546 938 3550 941
rect 3626 938 3630 941
rect 3518 928 3529 931
rect 3586 928 3590 931
rect 3358 872 3361 878
rect 3350 862 3353 868
rect 3374 861 3377 878
rect 3390 872 3393 878
rect 3414 872 3417 928
rect 3374 858 3382 861
rect 3350 802 3353 858
rect 3414 852 3417 868
rect 3422 852 3425 918
rect 3462 882 3465 888
rect 3450 868 3454 871
rect 3478 862 3481 898
rect 3518 882 3521 928
rect 3614 922 3617 928
rect 3622 918 3630 921
rect 3622 892 3625 918
rect 3646 902 3649 948
rect 3654 932 3657 938
rect 3530 888 3534 891
rect 3610 888 3614 891
rect 3534 872 3537 878
rect 3542 862 3545 878
rect 3566 872 3569 878
rect 3646 872 3649 888
rect 3666 878 3670 881
rect 3678 872 3681 948
rect 3686 942 3689 958
rect 3710 942 3713 1098
rect 3734 1082 3737 1088
rect 3718 1062 3721 1068
rect 3726 1022 3729 1078
rect 3742 1052 3745 1058
rect 3750 1022 3753 1058
rect 3758 1042 3761 1048
rect 3734 972 3737 998
rect 3722 968 3726 971
rect 3734 952 3737 958
rect 3718 942 3721 948
rect 3742 942 3745 1008
rect 3750 992 3753 998
rect 3766 962 3769 1078
rect 3774 1062 3777 1258
rect 3806 1232 3809 1248
rect 3790 1192 3793 1218
rect 3782 1152 3785 1188
rect 3794 1158 3801 1161
rect 3786 1148 3790 1151
rect 3798 1142 3801 1158
rect 3806 1152 3809 1188
rect 3786 1128 3790 1131
rect 3782 1072 3785 1118
rect 3790 1072 3793 1098
rect 3798 1082 3801 1138
rect 3822 1132 3825 1158
rect 3838 1152 3841 1268
rect 3878 1262 3881 1268
rect 3850 1248 3854 1251
rect 3886 1232 3889 1478
rect 3894 1452 3897 1518
rect 3902 1492 3905 1648
rect 3910 1532 3913 1718
rect 3958 1712 3961 1718
rect 3926 1672 3929 1678
rect 3950 1662 3953 1698
rect 4046 1681 4049 1718
rect 4054 1702 4057 1740
rect 4090 1718 4094 1721
rect 4058 1698 4065 1701
rect 4046 1678 4057 1681
rect 4054 1672 4057 1678
rect 3970 1668 3985 1671
rect 3958 1662 3961 1668
rect 3970 1658 3974 1661
rect 3926 1652 3929 1658
rect 3982 1652 3985 1668
rect 4022 1662 4025 1668
rect 4046 1662 4049 1668
rect 4062 1662 4065 1698
rect 4070 1672 4073 1718
rect 4080 1703 4082 1707
rect 4086 1703 4089 1707
rect 4093 1703 4096 1707
rect 4150 1672 4153 1878
rect 4158 1862 4161 1918
rect 4174 1862 4177 1928
rect 4206 1902 4209 1918
rect 4214 1882 4217 1928
rect 4198 1872 4201 1878
rect 4206 1862 4209 1878
rect 4230 1872 4233 1878
rect 4238 1872 4241 1948
rect 4302 1941 4305 1968
rect 4318 1962 4321 2068
rect 4342 2022 4345 2068
rect 4382 2062 4385 2078
rect 4446 2072 4449 2118
rect 4470 2092 4473 2148
rect 4498 2138 4502 2141
rect 4486 2132 4489 2138
rect 4470 2072 4473 2088
rect 4478 2072 4481 2128
rect 4486 2092 4489 2098
rect 4510 2082 4513 2118
rect 4518 2092 4521 2128
rect 4550 2122 4553 2248
rect 4558 2192 4561 2318
rect 4574 2262 4577 2298
rect 4582 2272 4585 2348
rect 4566 2242 4569 2248
rect 4574 2222 4577 2258
rect 4566 2072 4569 2138
rect 4590 2132 4593 2148
rect 4590 2092 4593 2128
rect 4598 2092 4601 2618
rect 4442 2068 4446 2071
rect 4570 2068 4574 2071
rect 4390 2062 4393 2068
rect 4378 2058 4382 2061
rect 4354 2048 4358 2051
rect 4406 2032 4409 2058
rect 4454 2052 4457 2058
rect 4462 2032 4465 2068
rect 4494 2062 4497 2068
rect 4510 2062 4513 2068
rect 4510 2048 4518 2051
rect 4326 1992 4329 2018
rect 4398 1982 4401 2018
rect 4282 1938 4305 1941
rect 4254 1922 4257 1938
rect 4294 1922 4297 1928
rect 4246 1892 4249 1908
rect 4222 1862 4225 1868
rect 4246 1852 4249 1868
rect 4254 1862 4257 1868
rect 4262 1862 4265 1868
rect 4270 1862 4273 1868
rect 4278 1862 4281 1878
rect 4162 1838 4166 1841
rect 4166 1752 4169 1768
rect 4174 1752 4177 1818
rect 4222 1792 4225 1818
rect 4206 1752 4209 1758
rect 4222 1742 4225 1778
rect 4246 1752 4249 1788
rect 4278 1752 4281 1848
rect 4286 1842 4289 1868
rect 4294 1862 4297 1898
rect 4310 1892 4313 1928
rect 4326 1882 4329 1948
rect 4318 1852 4321 1878
rect 4286 1792 4289 1838
rect 4310 1832 4313 1848
rect 4318 1782 4321 1848
rect 4310 1752 4313 1768
rect 4170 1738 4174 1741
rect 4194 1738 4198 1741
rect 4250 1738 4254 1741
rect 4098 1668 4102 1671
rect 4122 1658 4126 1661
rect 3990 1652 3993 1658
rect 4014 1652 4017 1658
rect 4078 1652 4081 1658
rect 3934 1642 3937 1648
rect 3950 1642 3953 1648
rect 3926 1562 3929 1578
rect 3982 1552 3985 1588
rect 3990 1552 3993 1648
rect 4014 1572 4017 1618
rect 4038 1561 4041 1618
rect 4034 1558 4041 1561
rect 3946 1548 3950 1551
rect 4010 1548 4014 1551
rect 3974 1542 3977 1548
rect 3998 1542 4001 1548
rect 3946 1538 3950 1541
rect 3970 1538 3974 1541
rect 3902 1472 3905 1478
rect 3910 1472 3913 1518
rect 3918 1492 3921 1528
rect 3918 1472 3921 1488
rect 3914 1458 3918 1461
rect 3926 1452 3929 1518
rect 3942 1462 3945 1528
rect 3950 1472 3953 1538
rect 4006 1532 4009 1538
rect 3998 1512 4001 1528
rect 3990 1482 3993 1498
rect 3998 1482 4001 1488
rect 4006 1482 4009 1518
rect 4022 1472 4025 1478
rect 4030 1462 4033 1548
rect 4046 1542 4049 1548
rect 4038 1522 4041 1538
rect 4038 1462 4041 1468
rect 4054 1462 4057 1648
rect 4070 1582 4073 1588
rect 4078 1552 4081 1648
rect 4134 1622 4137 1668
rect 4118 1552 4121 1618
rect 4126 1612 4129 1618
rect 4142 1602 4145 1668
rect 4174 1662 4177 1718
rect 4182 1692 4185 1738
rect 4154 1648 4158 1651
rect 4190 1641 4193 1718
rect 4198 1682 4201 1698
rect 4186 1638 4193 1641
rect 4166 1572 4169 1578
rect 4098 1548 4102 1551
rect 4154 1548 4158 1551
rect 4134 1542 4137 1548
rect 4150 1532 4153 1538
rect 4066 1528 4070 1531
rect 4174 1531 4177 1618
rect 4198 1592 4201 1668
rect 4206 1652 4209 1668
rect 4230 1652 4233 1718
rect 4238 1692 4241 1738
rect 4246 1682 4249 1698
rect 4246 1662 4249 1668
rect 4234 1618 4238 1621
rect 4254 1592 4257 1678
rect 4262 1672 4265 1748
rect 4318 1742 4321 1748
rect 4290 1738 4294 1741
rect 4290 1728 4294 1731
rect 4278 1722 4281 1728
rect 4286 1592 4289 1718
rect 4302 1662 4305 1718
rect 4326 1712 4329 1718
rect 4334 1692 4337 1758
rect 4342 1742 4345 1978
rect 4394 1968 4398 1971
rect 4406 1962 4409 2018
rect 4350 1932 4353 1948
rect 4350 1862 4353 1898
rect 4358 1872 4361 1938
rect 4366 1902 4369 1938
rect 4374 1912 4377 1948
rect 4362 1868 4366 1871
rect 4358 1858 4374 1861
rect 4358 1851 4361 1858
rect 4354 1848 4361 1851
rect 4366 1802 4369 1848
rect 4382 1842 4385 1918
rect 4398 1892 4401 1948
rect 4406 1942 4409 1948
rect 4414 1942 4417 1948
rect 4406 1932 4409 1938
rect 4422 1912 4425 2008
rect 4494 1972 4497 1978
rect 4406 1892 4409 1908
rect 4430 1902 4433 1928
rect 4442 1918 4446 1921
rect 4438 1892 4441 1908
rect 4462 1882 4465 1948
rect 4494 1942 4497 1948
rect 4486 1932 4489 1938
rect 4474 1928 4478 1931
rect 4450 1878 4454 1881
rect 4470 1881 4473 1918
rect 4510 1912 4513 2048
rect 4534 2012 4537 2058
rect 4542 2042 4545 2068
rect 4598 2062 4601 2078
rect 4562 2058 4566 2061
rect 4550 2042 4553 2048
rect 4566 1962 4569 2018
rect 4582 2012 4585 2058
rect 4530 1938 4534 1941
rect 4518 1922 4521 1928
rect 4510 1892 4513 1898
rect 4470 1878 4481 1881
rect 4434 1868 4438 1871
rect 4398 1862 4401 1868
rect 4414 1852 4417 1868
rect 4390 1772 4393 1778
rect 4398 1762 4401 1838
rect 4362 1748 4366 1751
rect 4394 1748 4398 1751
rect 4350 1742 4353 1748
rect 4374 1742 4377 1748
rect 4374 1732 4377 1738
rect 4366 1702 4369 1718
rect 4314 1678 4318 1681
rect 4358 1672 4361 1678
rect 4298 1638 4302 1641
rect 4294 1582 4297 1618
rect 4238 1572 4241 1578
rect 4202 1568 4206 1571
rect 4222 1562 4225 1568
rect 4186 1548 4190 1551
rect 4210 1548 4214 1551
rect 4170 1528 4177 1531
rect 4062 1472 4065 1508
rect 4080 1503 4082 1507
rect 4086 1503 4089 1507
rect 4093 1503 4096 1507
rect 4126 1492 4129 1508
rect 4134 1502 4137 1528
rect 4182 1522 4185 1538
rect 4118 1472 4121 1488
rect 4142 1472 4145 1518
rect 4198 1492 4201 1548
rect 4230 1542 4233 1548
rect 4114 1468 4118 1471
rect 4062 1462 4065 1468
rect 3970 1458 3974 1461
rect 4010 1458 4014 1461
rect 4026 1458 4030 1461
rect 3958 1452 3961 1458
rect 3986 1448 3990 1451
rect 3942 1392 3945 1418
rect 3982 1392 3985 1438
rect 4006 1392 4009 1448
rect 3926 1382 3929 1388
rect 3926 1352 3929 1378
rect 3898 1348 3905 1351
rect 3946 1348 3950 1351
rect 3902 1262 3905 1348
rect 3966 1342 3969 1348
rect 3974 1342 3977 1368
rect 3990 1352 3993 1358
rect 3998 1342 4001 1358
rect 3910 1332 3913 1338
rect 3962 1328 3966 1331
rect 3934 1272 3937 1318
rect 3942 1312 3945 1328
rect 3950 1312 3953 1328
rect 4014 1322 4017 1358
rect 4054 1352 4057 1458
rect 4134 1452 4137 1468
rect 4150 1452 4153 1458
rect 4158 1452 4161 1458
rect 4166 1452 4169 1468
rect 4178 1458 4182 1461
rect 4206 1452 4209 1498
rect 4238 1492 4241 1548
rect 4254 1522 4257 1558
rect 4262 1492 4265 1548
rect 4286 1542 4289 1558
rect 4294 1542 4297 1558
rect 4318 1552 4321 1668
rect 4366 1662 4369 1668
rect 4382 1662 4385 1678
rect 4366 1592 4369 1658
rect 4374 1632 4377 1658
rect 4382 1621 4385 1658
rect 4406 1652 4409 1708
rect 4414 1692 4417 1758
rect 4422 1752 4425 1858
rect 4446 1812 4449 1868
rect 4462 1842 4465 1878
rect 4478 1872 4481 1878
rect 4486 1872 4489 1888
rect 4514 1878 4518 1881
rect 4502 1872 4505 1878
rect 4470 1852 4473 1868
rect 4478 1862 4481 1868
rect 4438 1792 4441 1798
rect 4430 1742 4433 1778
rect 4454 1772 4457 1818
rect 4446 1722 4449 1768
rect 4454 1752 4457 1758
rect 4486 1752 4489 1848
rect 4494 1742 4497 1868
rect 4526 1862 4529 1888
rect 4542 1882 4545 1938
rect 4550 1932 4553 1948
rect 4558 1922 4561 1948
rect 4566 1942 4569 1958
rect 4582 1932 4585 1938
rect 4558 1882 4561 1918
rect 4558 1871 4561 1878
rect 4554 1868 4561 1871
rect 4542 1862 4545 1868
rect 4566 1862 4569 1928
rect 4558 1842 4561 1848
rect 4534 1762 4537 1818
rect 4558 1792 4561 1828
rect 4426 1678 4430 1681
rect 4414 1672 4417 1678
rect 4450 1668 4454 1671
rect 4462 1662 4465 1698
rect 4486 1662 4489 1728
rect 4502 1692 4505 1758
rect 4518 1742 4521 1748
rect 4542 1742 4545 1748
rect 4566 1742 4569 1858
rect 4574 1852 4577 1918
rect 4582 1882 4585 1888
rect 4598 1862 4601 1868
rect 4498 1668 4502 1671
rect 4526 1662 4529 1668
rect 4534 1662 4537 1738
rect 4574 1732 4577 1758
rect 4590 1752 4593 1818
rect 4554 1658 4558 1661
rect 4414 1652 4417 1658
rect 4522 1648 4526 1651
rect 4538 1638 4542 1641
rect 4374 1618 4385 1621
rect 4374 1572 4377 1618
rect 4326 1552 4329 1568
rect 4398 1562 4401 1568
rect 4426 1558 4430 1561
rect 4462 1558 4470 1561
rect 4350 1552 4353 1558
rect 4462 1552 4465 1558
rect 4486 1552 4489 1618
rect 4510 1562 4513 1598
rect 4410 1548 4414 1551
rect 4474 1548 4478 1551
rect 4274 1538 4278 1541
rect 4286 1522 4289 1528
rect 4278 1492 4281 1508
rect 4310 1492 4313 1548
rect 4266 1478 4270 1481
rect 4246 1472 4249 1478
rect 4234 1468 4238 1471
rect 4254 1462 4257 1468
rect 4262 1462 4265 1468
rect 4238 1458 4246 1461
rect 4130 1448 4134 1451
rect 4174 1442 4177 1448
rect 4190 1432 4193 1438
rect 4026 1348 4030 1351
rect 4038 1312 4041 1348
rect 4046 1342 4049 1348
rect 4054 1342 4057 1348
rect 4046 1322 4049 1338
rect 4062 1312 4065 1348
rect 3998 1292 4001 1298
rect 3942 1272 3945 1278
rect 3974 1272 3977 1278
rect 4014 1270 4017 1278
rect 3950 1262 3953 1268
rect 3914 1258 3918 1261
rect 3930 1258 3934 1261
rect 3970 1258 3974 1261
rect 3902 1242 3905 1258
rect 3914 1248 3918 1251
rect 3862 1162 3865 1208
rect 3894 1152 3897 1188
rect 3926 1162 3929 1218
rect 3942 1172 3945 1188
rect 3914 1158 3918 1161
rect 3902 1152 3905 1158
rect 3842 1148 3846 1151
rect 3806 1078 3814 1081
rect 3830 1072 3833 1128
rect 3846 1112 3849 1138
rect 3870 1132 3873 1148
rect 3886 1132 3889 1148
rect 3910 1142 3913 1158
rect 3890 1128 3894 1131
rect 3854 1112 3857 1118
rect 3850 1088 3854 1091
rect 3878 1082 3881 1088
rect 3774 1052 3777 1058
rect 3782 972 3785 1068
rect 3790 1062 3793 1068
rect 3830 1052 3833 1068
rect 3838 1062 3841 1068
rect 3862 1062 3865 1068
rect 3878 1062 3881 1068
rect 3894 1062 3897 1128
rect 3902 1072 3905 1078
rect 3918 1072 3921 1098
rect 3926 1082 3929 1158
rect 3914 1068 3918 1071
rect 3794 1048 3798 1051
rect 3842 1048 3846 1051
rect 3798 962 3801 968
rect 3754 948 3758 951
rect 3782 942 3785 948
rect 3798 942 3801 948
rect 3746 938 3750 941
rect 3694 922 3697 928
rect 3694 892 3697 908
rect 3710 892 3713 938
rect 3774 932 3777 938
rect 3806 932 3809 998
rect 3910 981 3913 1068
rect 3918 1052 3921 1058
rect 3926 1042 3929 1058
rect 3934 1052 3937 1118
rect 3942 1102 3945 1138
rect 3950 1081 3953 1218
rect 3966 1172 3969 1248
rect 3990 1242 3993 1258
rect 4022 1242 4025 1268
rect 4030 1252 4033 1268
rect 3966 1122 3969 1148
rect 3974 1142 3977 1208
rect 3994 1158 3998 1161
rect 4006 1152 4009 1158
rect 4038 1152 4041 1308
rect 4054 1262 4057 1268
rect 4062 1262 4065 1268
rect 4046 1252 4049 1258
rect 4058 1248 4062 1251
rect 4046 1202 4049 1218
rect 4070 1212 4073 1418
rect 4090 1388 4094 1391
rect 4138 1358 4142 1361
rect 4166 1352 4169 1358
rect 4182 1352 4185 1408
rect 4198 1392 4201 1398
rect 4098 1328 4102 1331
rect 4080 1303 4082 1307
rect 4086 1303 4089 1307
rect 4093 1303 4096 1307
rect 4118 1292 4121 1348
rect 4126 1292 4129 1338
rect 4150 1332 4153 1338
rect 4174 1332 4177 1348
rect 4138 1318 4142 1321
rect 4150 1272 4153 1328
rect 4166 1302 4169 1318
rect 4090 1268 4094 1271
rect 4078 1262 4081 1268
rect 4014 1142 4017 1148
rect 4042 1138 4049 1141
rect 3942 1078 3953 1081
rect 3942 1052 3945 1078
rect 3974 1072 3977 1138
rect 3990 1092 3993 1128
rect 4030 1102 4033 1128
rect 3990 1082 3993 1088
rect 3954 1068 3958 1071
rect 4014 1062 4017 1068
rect 3962 1058 3966 1061
rect 3986 1058 3990 1061
rect 4006 1052 4009 1058
rect 4038 1052 4041 1108
rect 4046 1082 4049 1138
rect 4062 1082 4065 1188
rect 4070 1162 4073 1168
rect 4054 1071 4057 1078
rect 4050 1068 4057 1071
rect 4062 1062 4065 1068
rect 4046 1052 4049 1058
rect 3946 1018 3950 1021
rect 3902 978 3913 981
rect 3862 962 3865 968
rect 3874 958 3878 961
rect 3830 952 3833 958
rect 3902 952 3905 978
rect 3910 962 3913 968
rect 3934 962 3937 968
rect 3842 948 3846 951
rect 3814 922 3817 928
rect 3742 918 3750 921
rect 3742 892 3745 918
rect 3782 892 3785 898
rect 3806 892 3809 898
rect 3698 868 3702 871
rect 3430 858 3438 861
rect 3386 848 3390 851
rect 3246 732 3249 738
rect 3286 732 3289 738
rect 3266 728 3270 731
rect 3238 718 3249 721
rect 3238 692 3241 708
rect 3246 672 3249 718
rect 3270 682 3273 688
rect 3294 672 3297 708
rect 3210 668 3214 671
rect 3166 562 3169 658
rect 3182 642 3185 648
rect 3190 602 3193 668
rect 3222 662 3225 668
rect 3258 658 3262 661
rect 3278 651 3281 668
rect 3286 662 3289 668
rect 3278 648 3289 651
rect 3206 612 3209 648
rect 3222 592 3225 618
rect 3238 582 3241 648
rect 3270 581 3273 648
rect 3278 592 3281 638
rect 3286 592 3289 648
rect 3302 592 3305 738
rect 3318 662 3321 738
rect 3334 722 3337 748
rect 3342 732 3345 738
rect 3326 672 3329 708
rect 3342 692 3345 718
rect 3350 672 3353 798
rect 3366 751 3369 848
rect 3398 792 3401 848
rect 3362 748 3369 751
rect 3366 712 3369 718
rect 3374 692 3377 768
rect 3382 752 3385 758
rect 3398 742 3401 748
rect 3394 738 3398 741
rect 3358 672 3361 678
rect 3350 662 3353 668
rect 3310 622 3313 648
rect 3334 622 3337 648
rect 3318 582 3321 588
rect 3270 578 3281 581
rect 3186 558 3190 561
rect 3206 552 3209 558
rect 3194 548 3198 551
rect 3066 458 3070 461
rect 3078 392 3081 398
rect 3066 358 3073 361
rect 2978 338 2982 341
rect 2966 312 2969 328
rect 2982 272 2985 278
rect 2990 272 2993 338
rect 3006 322 3009 358
rect 3014 292 3017 358
rect 3030 352 3033 358
rect 3030 272 3033 348
rect 3038 332 3041 338
rect 3048 303 3050 307
rect 3054 303 3057 307
rect 3061 303 3064 307
rect 3070 292 3073 358
rect 3086 352 3089 468
rect 3094 462 3097 468
rect 3102 412 3105 458
rect 3118 452 3121 488
rect 3126 472 3129 478
rect 3134 462 3137 468
rect 3126 448 3134 451
rect 3110 392 3113 448
rect 3098 348 3102 351
rect 3078 282 3081 348
rect 3086 332 3089 338
rect 3086 292 3089 318
rect 3110 292 3113 308
rect 3126 292 3129 448
rect 3158 422 3161 448
rect 3158 382 3161 418
rect 3166 412 3169 548
rect 3182 532 3185 548
rect 3174 528 3182 531
rect 3174 472 3177 528
rect 3190 522 3193 538
rect 3182 492 3185 508
rect 3206 472 3209 528
rect 3222 492 3225 578
rect 3266 558 3270 561
rect 3266 548 3270 551
rect 3230 542 3233 548
rect 3246 542 3249 548
rect 3250 538 3254 541
rect 3246 482 3249 488
rect 3234 478 3238 481
rect 3254 472 3257 478
rect 3182 402 3185 448
rect 3142 352 3145 358
rect 3150 352 3153 378
rect 3162 368 3166 371
rect 3190 362 3193 448
rect 3198 422 3201 458
rect 3198 392 3201 398
rect 3170 348 3174 351
rect 3134 322 3137 348
rect 3038 272 3041 278
rect 3090 268 3094 271
rect 2926 252 2929 258
rect 2934 192 2937 218
rect 2890 188 2894 191
rect 2790 142 2793 148
rect 2806 142 2809 158
rect 2842 148 2846 151
rect 2714 138 2718 141
rect 2778 138 2782 141
rect 2810 138 2817 141
rect 2594 128 2598 131
rect 2642 128 2646 131
rect 2574 92 2577 108
rect 2598 92 2601 118
rect 2614 92 2617 128
rect 2638 102 2641 118
rect 2430 82 2433 88
rect 2470 82 2473 88
rect 2386 78 2390 81
rect 2310 62 2313 68
rect 2366 62 2369 68
rect 2390 62 2393 78
rect 2502 72 2505 78
rect 2534 72 2537 78
rect 2622 72 2625 78
rect 2630 72 2633 88
rect 2402 68 2406 71
rect 2418 68 2422 71
rect 2586 68 2590 71
rect 2526 62 2529 68
rect 2242 58 2246 61
rect 2330 58 2334 61
rect 2254 52 2257 58
rect 2454 52 2457 58
rect 2194 48 2198 51
rect 2242 48 2246 51
rect 2534 51 2537 58
rect 2530 48 2537 51
rect 2334 42 2337 48
rect 2486 42 2489 48
rect 2034 38 2038 41
rect 2558 41 2561 58
rect 2574 52 2577 68
rect 2638 62 2641 98
rect 2694 92 2697 98
rect 2718 92 2721 128
rect 2670 88 2689 91
rect 2650 78 2654 81
rect 2662 72 2665 88
rect 2670 82 2673 88
rect 2686 82 2689 88
rect 2734 82 2737 98
rect 2678 52 2681 78
rect 2766 72 2769 78
rect 2790 72 2793 138
rect 2814 132 2817 138
rect 2854 132 2857 178
rect 2878 162 2881 168
rect 2926 162 2929 168
rect 2862 142 2865 148
rect 2918 142 2921 158
rect 2942 152 2945 268
rect 2954 248 2958 251
rect 2966 242 2969 248
rect 2958 238 2966 241
rect 2958 192 2961 238
rect 2958 152 2961 168
rect 2974 162 2977 168
rect 2946 148 2950 151
rect 2982 142 2985 188
rect 2990 162 2993 268
rect 3102 252 3105 288
rect 3122 268 3126 271
rect 3002 248 3006 251
rect 3046 248 3054 251
rect 3014 242 3017 248
rect 2998 161 3001 218
rect 3022 192 3025 198
rect 3046 192 3049 248
rect 3118 232 3121 268
rect 2998 158 3006 161
rect 3026 158 3030 161
rect 2990 152 2993 158
rect 3054 152 3057 228
rect 3062 142 3065 198
rect 3086 192 3089 218
rect 3126 202 3129 248
rect 3134 191 3137 298
rect 3150 292 3153 328
rect 3190 302 3193 358
rect 3198 272 3201 378
rect 3206 342 3209 468
rect 3218 448 3222 451
rect 3230 442 3233 468
rect 3270 462 3273 528
rect 3278 492 3281 578
rect 3302 552 3305 558
rect 3318 542 3321 548
rect 3294 522 3297 528
rect 3294 482 3297 488
rect 3318 482 3321 538
rect 3290 468 3294 471
rect 3258 458 3262 461
rect 3306 458 3310 461
rect 3298 448 3302 451
rect 3238 352 3241 408
rect 3262 392 3265 448
rect 3270 372 3273 448
rect 3318 442 3321 468
rect 3326 462 3329 598
rect 3334 462 3337 608
rect 3350 542 3353 658
rect 3366 552 3369 678
rect 3382 662 3385 668
rect 3374 572 3377 648
rect 3350 532 3353 538
rect 3342 512 3345 528
rect 3358 522 3361 548
rect 3374 541 3377 568
rect 3390 561 3393 718
rect 3398 661 3401 738
rect 3406 732 3409 798
rect 3414 792 3417 838
rect 3430 832 3433 858
rect 3498 848 3502 851
rect 3438 822 3441 828
rect 3414 758 3422 761
rect 3414 672 3417 758
rect 3430 752 3433 758
rect 3462 752 3465 758
rect 3494 752 3497 818
rect 3510 812 3513 858
rect 3542 802 3545 858
rect 3550 832 3553 848
rect 3550 792 3553 818
rect 3510 752 3513 758
rect 3422 742 3425 748
rect 3438 742 3441 748
rect 3438 672 3441 708
rect 3426 668 3430 671
rect 3398 658 3409 661
rect 3418 658 3422 661
rect 3398 642 3401 648
rect 3398 592 3401 618
rect 3386 558 3393 561
rect 3406 552 3409 658
rect 3454 652 3457 698
rect 3462 692 3465 738
rect 3470 732 3473 738
rect 3478 702 3481 738
rect 3486 722 3489 748
rect 3486 672 3489 718
rect 3502 692 3505 698
rect 3518 692 3521 788
rect 3526 722 3529 738
rect 3534 702 3537 758
rect 3558 742 3561 868
rect 3566 862 3569 868
rect 3590 862 3593 868
rect 3638 862 3641 868
rect 3642 858 3646 861
rect 3654 852 3657 858
rect 3578 848 3582 851
rect 3610 848 3614 851
rect 3666 848 3670 851
rect 3568 803 3570 807
rect 3574 803 3577 807
rect 3581 803 3584 807
rect 3566 731 3569 768
rect 3590 732 3593 808
rect 3598 752 3601 758
rect 3622 752 3625 848
rect 3654 792 3657 828
rect 3678 762 3681 868
rect 3690 848 3694 851
rect 3686 752 3689 798
rect 3698 748 3702 751
rect 3602 738 3606 741
rect 3558 728 3569 731
rect 3582 728 3590 731
rect 3558 692 3561 728
rect 3582 692 3585 728
rect 3614 722 3617 748
rect 3622 732 3625 738
rect 3638 732 3641 740
rect 3590 672 3593 718
rect 3606 692 3609 698
rect 3614 692 3617 708
rect 3638 672 3641 728
rect 3670 722 3673 728
rect 3658 678 3662 681
rect 3534 668 3542 671
rect 3666 668 3670 671
rect 3478 662 3481 668
rect 3510 662 3513 668
rect 3446 648 3454 651
rect 3490 648 3494 651
rect 3446 592 3449 648
rect 3478 592 3481 638
rect 3454 582 3457 588
rect 3366 538 3377 541
rect 3358 492 3361 518
rect 3346 458 3350 461
rect 3302 392 3305 398
rect 3246 342 3249 348
rect 3206 302 3209 338
rect 3222 272 3225 318
rect 3254 312 3257 348
rect 3238 272 3241 278
rect 3146 268 3150 271
rect 3186 268 3190 271
rect 3226 268 3233 271
rect 3130 188 3137 191
rect 3150 192 3153 248
rect 3078 142 3081 188
rect 3162 168 3166 171
rect 3110 162 3113 168
rect 3098 158 3102 161
rect 3130 148 3134 151
rect 2946 138 2950 141
rect 2782 62 2785 68
rect 2754 58 2758 61
rect 2786 58 2798 61
rect 2702 52 2705 58
rect 2582 48 2598 51
rect 2806 51 2809 108
rect 2814 62 2817 68
rect 2830 61 2833 108
rect 2854 72 2857 128
rect 2878 92 2881 98
rect 2910 82 2913 98
rect 2918 92 2921 108
rect 2926 82 2929 98
rect 2842 68 2846 71
rect 2882 68 2886 71
rect 2942 62 2945 128
rect 2974 82 2977 98
rect 2998 92 3001 138
rect 3038 112 3041 138
rect 3048 103 3050 107
rect 3054 103 3057 107
rect 3061 103 3064 107
rect 3086 92 3089 148
rect 3130 138 3134 141
rect 3142 141 3145 158
rect 3174 152 3177 268
rect 3230 262 3233 268
rect 3246 262 3249 298
rect 3262 292 3265 358
rect 3278 342 3281 348
rect 3294 342 3297 358
rect 3302 332 3305 348
rect 3294 292 3297 298
rect 3194 258 3198 261
rect 3218 258 3222 261
rect 3254 252 3257 258
rect 3218 248 3222 251
rect 3206 241 3209 248
rect 3206 238 3217 241
rect 3214 192 3217 238
rect 3186 158 3190 161
rect 3138 138 3145 141
rect 3166 142 3169 148
rect 3134 92 3137 108
rect 3098 78 3102 81
rect 2830 58 2838 61
rect 2938 58 2942 61
rect 2958 52 2961 68
rect 2982 62 2985 68
rect 3038 62 3041 68
rect 3070 62 3073 78
rect 3102 72 3105 78
rect 3142 72 3145 78
rect 3158 72 3161 98
rect 3182 92 3185 138
rect 3190 132 3193 158
rect 3230 152 3233 168
rect 3246 162 3249 198
rect 3294 192 3297 248
rect 3302 222 3305 328
rect 3310 272 3313 438
rect 3318 292 3321 358
rect 3342 342 3345 378
rect 3358 332 3361 458
rect 3366 392 3369 538
rect 3374 452 3377 498
rect 3382 492 3385 548
rect 3414 542 3417 558
rect 3402 538 3406 541
rect 3390 472 3393 528
rect 3398 492 3401 498
rect 3406 492 3409 538
rect 3390 382 3393 468
rect 3402 448 3406 451
rect 3414 392 3417 528
rect 3430 502 3433 558
rect 3454 542 3457 548
rect 3470 542 3473 558
rect 3422 472 3425 498
rect 3438 472 3441 478
rect 3430 462 3433 468
rect 3438 462 3441 468
rect 3454 462 3457 478
rect 3462 472 3465 488
rect 3478 472 3481 548
rect 3486 542 3489 558
rect 3494 542 3497 558
rect 3510 552 3513 648
rect 3534 562 3537 668
rect 3542 592 3545 658
rect 3550 622 3553 648
rect 3568 603 3570 607
rect 3574 603 3577 607
rect 3581 603 3584 607
rect 3586 558 3590 561
rect 3518 532 3521 558
rect 3542 552 3545 558
rect 3542 542 3545 548
rect 3598 542 3601 668
rect 3686 662 3689 748
rect 3694 672 3697 718
rect 3710 682 3713 888
rect 3750 882 3753 888
rect 3774 882 3777 888
rect 3734 872 3737 878
rect 3822 872 3825 878
rect 3830 872 3833 938
rect 3846 932 3849 938
rect 3726 862 3729 868
rect 3758 862 3761 868
rect 3798 862 3801 868
rect 3718 792 3721 818
rect 3726 772 3729 848
rect 3762 838 3766 841
rect 3782 832 3785 848
rect 3754 758 3758 761
rect 3782 752 3785 758
rect 3798 752 3801 858
rect 3806 852 3809 868
rect 3826 858 3830 861
rect 3838 852 3841 858
rect 3806 832 3809 848
rect 3738 748 3742 751
rect 3726 742 3729 748
rect 3746 738 3750 741
rect 3794 738 3798 741
rect 3774 732 3777 738
rect 3806 731 3809 828
rect 3822 752 3825 838
rect 3834 788 3838 791
rect 3846 772 3849 898
rect 3854 762 3857 878
rect 3862 872 3865 878
rect 3862 832 3865 858
rect 3870 842 3873 868
rect 3870 792 3873 828
rect 3834 758 3838 761
rect 3798 728 3809 731
rect 3798 712 3801 728
rect 3806 712 3809 718
rect 3830 692 3833 708
rect 3810 688 3814 691
rect 3714 668 3718 671
rect 3750 662 3753 688
rect 3790 678 3798 681
rect 3766 662 3769 668
rect 3630 652 3633 658
rect 3674 648 3678 651
rect 3606 552 3609 648
rect 3614 642 3617 648
rect 3618 558 3622 561
rect 3518 491 3521 528
rect 3510 488 3521 491
rect 3502 462 3505 488
rect 3446 458 3454 461
rect 3466 458 3470 461
rect 3490 458 3494 461
rect 3366 322 3369 348
rect 3374 342 3377 378
rect 3398 362 3401 368
rect 3382 342 3385 358
rect 3406 342 3409 358
rect 3394 328 3398 331
rect 3366 292 3369 318
rect 3386 278 3390 281
rect 3346 268 3350 271
rect 3378 268 3382 271
rect 3318 242 3321 248
rect 3334 242 3337 268
rect 3390 262 3393 268
rect 3346 258 3350 261
rect 3334 172 3337 238
rect 3258 158 3262 161
rect 3274 158 3278 161
rect 3238 152 3241 158
rect 3286 152 3289 168
rect 3318 162 3321 168
rect 3198 142 3201 148
rect 3226 138 3230 141
rect 3270 122 3273 148
rect 3294 141 3297 158
rect 3334 152 3337 158
rect 3290 138 3297 141
rect 3342 142 3345 228
rect 3350 162 3353 258
rect 3366 192 3369 248
rect 3350 152 3353 158
rect 3222 92 3225 108
rect 3270 102 3273 108
rect 3278 102 3281 138
rect 3194 78 3198 81
rect 3166 72 3169 78
rect 3206 72 3209 78
rect 3230 72 3233 98
rect 3270 82 3273 98
rect 3278 92 3281 98
rect 3294 92 3297 118
rect 3258 78 3262 81
rect 3026 58 3030 61
rect 3006 52 3009 58
rect 3038 52 3041 58
rect 3126 52 3129 58
rect 3254 52 3257 68
rect 3278 52 3281 68
rect 3302 62 3305 88
rect 3310 71 3313 108
rect 3358 92 3361 168
rect 3366 152 3369 158
rect 3374 142 3377 228
rect 3398 192 3401 308
rect 3406 292 3409 318
rect 3414 292 3417 348
rect 3430 292 3433 358
rect 3438 332 3441 358
rect 3446 352 3449 458
rect 3454 392 3457 448
rect 3462 362 3465 458
rect 3478 448 3486 451
rect 3462 352 3465 358
rect 3454 338 3462 341
rect 3454 322 3457 338
rect 3438 281 3441 288
rect 3470 282 3473 338
rect 3478 292 3481 448
rect 3490 348 3494 351
rect 3510 341 3513 488
rect 3542 472 3545 508
rect 3582 492 3585 528
rect 3558 462 3561 468
rect 3606 461 3609 538
rect 3630 502 3633 518
rect 3622 482 3625 488
rect 3602 458 3609 461
rect 3622 462 3625 468
rect 3630 462 3633 498
rect 3646 462 3649 548
rect 3654 542 3657 638
rect 3670 562 3673 568
rect 3662 532 3665 558
rect 3678 542 3681 598
rect 3686 592 3689 608
rect 3702 582 3705 658
rect 3698 568 3702 571
rect 3710 552 3713 558
rect 3718 552 3721 648
rect 3726 642 3729 658
rect 3678 462 3681 468
rect 3526 442 3529 458
rect 3566 421 3569 458
rect 3558 418 3569 421
rect 3518 372 3521 418
rect 3558 362 3561 418
rect 3568 403 3570 407
rect 3574 403 3577 407
rect 3581 403 3584 407
rect 3598 402 3601 458
rect 3606 392 3609 418
rect 3662 381 3665 458
rect 3670 452 3673 458
rect 3690 448 3694 451
rect 3670 392 3673 428
rect 3702 422 3705 548
rect 3718 532 3721 548
rect 3734 542 3737 638
rect 3742 572 3745 618
rect 3758 601 3761 658
rect 3750 598 3761 601
rect 3726 522 3729 528
rect 3742 482 3745 488
rect 3750 462 3753 598
rect 3766 591 3769 608
rect 3790 602 3793 678
rect 3798 672 3801 678
rect 3806 661 3809 678
rect 3838 672 3841 738
rect 3846 722 3849 748
rect 3858 728 3862 731
rect 3878 692 3881 918
rect 3886 862 3889 948
rect 3902 942 3905 948
rect 3910 942 3913 948
rect 3950 942 3953 948
rect 3894 932 3897 938
rect 3950 882 3953 938
rect 3958 882 3961 1048
rect 3982 1002 3985 1048
rect 4006 1031 4009 1048
rect 4002 1028 4009 1031
rect 4006 992 4009 1008
rect 4070 1002 4073 1158
rect 4078 1142 4081 1238
rect 4102 1172 4105 1248
rect 4110 1192 4113 1258
rect 4102 1152 4105 1168
rect 4118 1142 4121 1148
rect 4126 1142 4129 1228
rect 4110 1132 4113 1138
rect 4134 1132 4137 1268
rect 4142 1252 4145 1258
rect 4142 1212 4145 1218
rect 4150 1202 4153 1268
rect 4158 1252 4161 1278
rect 4166 1262 4169 1268
rect 4182 1252 4185 1258
rect 4190 1252 4193 1388
rect 4206 1332 4209 1448
rect 4222 1432 4225 1438
rect 4230 1422 4233 1458
rect 4238 1452 4241 1458
rect 4286 1422 4289 1468
rect 4294 1462 4297 1488
rect 4306 1458 4310 1461
rect 4294 1452 4297 1458
rect 4234 1388 4238 1391
rect 4246 1362 4249 1368
rect 4266 1358 4270 1361
rect 4230 1352 4233 1358
rect 4286 1352 4289 1388
rect 4318 1361 4321 1548
rect 4346 1528 4350 1531
rect 4342 1472 4345 1478
rect 4310 1358 4321 1361
rect 4330 1468 4334 1471
rect 4214 1292 4217 1348
rect 4226 1338 4230 1341
rect 4230 1272 4233 1318
rect 4254 1292 4257 1348
rect 4278 1342 4281 1348
rect 4274 1328 4278 1331
rect 4238 1282 4241 1288
rect 4278 1282 4281 1318
rect 4146 1178 4150 1181
rect 4146 1158 4150 1161
rect 4150 1142 4153 1158
rect 4166 1152 4169 1238
rect 4194 1228 4198 1231
rect 4174 1222 4177 1228
rect 4182 1152 4185 1178
rect 4198 1161 4201 1218
rect 4206 1182 4209 1268
rect 4266 1258 4270 1261
rect 4278 1252 4281 1258
rect 4286 1232 4289 1348
rect 4294 1252 4297 1258
rect 4214 1222 4217 1228
rect 4302 1222 4305 1318
rect 4310 1272 4313 1358
rect 4318 1342 4321 1348
rect 4326 1332 4329 1468
rect 4338 1458 4342 1461
rect 4358 1442 4361 1448
rect 4334 1392 4337 1438
rect 4366 1371 4369 1538
rect 4390 1532 4393 1538
rect 4382 1482 4385 1518
rect 4398 1492 4401 1498
rect 4406 1482 4409 1538
rect 4446 1482 4449 1548
rect 4510 1542 4513 1558
rect 4566 1552 4569 1718
rect 4574 1682 4577 1728
rect 4590 1692 4593 1728
rect 4594 1678 4598 1681
rect 4582 1662 4585 1668
rect 4518 1548 4526 1551
rect 4466 1538 4470 1541
rect 4490 1538 4494 1541
rect 4454 1532 4457 1538
rect 4394 1468 4398 1471
rect 4434 1468 4438 1471
rect 4374 1462 4377 1468
rect 4414 1462 4417 1468
rect 4382 1452 4385 1458
rect 4422 1452 4425 1458
rect 4434 1448 4438 1451
rect 4446 1382 4449 1478
rect 4454 1442 4457 1528
rect 4462 1472 4465 1478
rect 4494 1472 4497 1478
rect 4486 1462 4489 1468
rect 4502 1462 4505 1468
rect 4462 1412 4465 1458
rect 4470 1452 4473 1458
rect 4478 1452 4481 1458
rect 4518 1452 4521 1548
rect 4534 1492 4537 1538
rect 4542 1472 4545 1518
rect 4550 1492 4553 1548
rect 4558 1532 4561 1538
rect 4570 1528 4574 1531
rect 4554 1468 4558 1471
rect 4586 1468 4590 1471
rect 4506 1448 4510 1451
rect 4470 1401 4473 1448
rect 4462 1398 4473 1401
rect 4462 1392 4465 1398
rect 4366 1368 4374 1371
rect 4318 1292 4321 1298
rect 4326 1272 4329 1308
rect 4334 1302 4337 1368
rect 4374 1362 4377 1368
rect 4350 1352 4353 1358
rect 4342 1342 4345 1348
rect 4350 1291 4353 1348
rect 4358 1311 4361 1348
rect 4390 1342 4393 1378
rect 4494 1362 4497 1368
rect 4410 1358 4414 1361
rect 4474 1348 4478 1351
rect 4398 1332 4401 1348
rect 4430 1342 4433 1348
rect 4454 1342 4457 1348
rect 4486 1332 4489 1358
rect 4510 1352 4513 1438
rect 4518 1392 4521 1448
rect 4526 1392 4529 1468
rect 4538 1458 4542 1461
rect 4550 1452 4553 1458
rect 4566 1442 4569 1448
rect 4518 1352 4521 1358
rect 4498 1348 4502 1351
rect 4510 1342 4513 1348
rect 4502 1338 4510 1341
rect 4358 1308 4366 1311
rect 4350 1288 4361 1291
rect 4334 1232 4337 1258
rect 4342 1252 4345 1268
rect 4214 1162 4217 1208
rect 4198 1158 4209 1161
rect 4194 1148 4198 1151
rect 4166 1142 4169 1148
rect 4174 1132 4177 1138
rect 4138 1128 4142 1131
rect 4154 1128 4158 1131
rect 4080 1103 4082 1107
rect 4086 1103 4089 1107
rect 4093 1103 4096 1107
rect 4110 1082 4113 1128
rect 4082 1078 4086 1081
rect 4098 1068 4102 1071
rect 4118 1062 4121 1128
rect 4126 1092 4129 1098
rect 4190 1082 4193 1148
rect 4206 1142 4209 1158
rect 4222 1142 4225 1178
rect 4254 1172 4257 1218
rect 4226 1138 4230 1141
rect 4234 1128 4238 1131
rect 4198 1082 4201 1118
rect 4138 1078 4142 1081
rect 4158 1072 4161 1078
rect 4166 1072 4169 1078
rect 4070 962 4073 998
rect 3978 948 3982 951
rect 3942 872 3945 878
rect 3966 862 3969 918
rect 3990 892 3993 958
rect 4094 952 4097 958
rect 4002 948 4006 951
rect 4014 942 4017 948
rect 4054 942 4057 948
rect 4022 932 4025 938
rect 4034 928 4038 931
rect 3982 872 3985 878
rect 3986 868 3993 871
rect 3990 862 3993 868
rect 3890 858 3894 861
rect 3938 858 3942 861
rect 3982 852 3985 858
rect 3914 848 3918 851
rect 3962 848 3966 851
rect 3886 842 3889 848
rect 3962 838 3966 841
rect 3906 788 3910 791
rect 3886 682 3889 758
rect 3942 752 3945 838
rect 3990 832 3993 848
rect 3978 788 3982 791
rect 3998 772 4001 888
rect 4022 882 4025 928
rect 4038 892 4041 908
rect 4046 902 4049 918
rect 4014 832 4017 868
rect 4022 862 4025 878
rect 4038 842 4041 848
rect 4046 812 4049 868
rect 4058 858 4062 861
rect 4070 861 4073 948
rect 4090 938 4094 941
rect 4080 903 4082 907
rect 4086 903 4089 907
rect 4093 903 4096 907
rect 4102 872 4105 1038
rect 4118 952 4121 1048
rect 4134 1012 4137 1068
rect 4182 1062 4185 1068
rect 4202 1058 4206 1061
rect 4214 1042 4217 1118
rect 4194 1028 4198 1031
rect 4222 1031 4225 1068
rect 4238 1052 4241 1128
rect 4254 1102 4257 1168
rect 4274 1158 4278 1161
rect 4294 1152 4297 1198
rect 4350 1182 4353 1278
rect 4358 1272 4361 1288
rect 4374 1272 4377 1278
rect 4390 1262 4393 1268
rect 4406 1262 4409 1288
rect 4438 1262 4441 1268
rect 4358 1258 4366 1261
rect 4310 1162 4313 1178
rect 4350 1152 4353 1178
rect 4358 1152 4361 1258
rect 4374 1192 4377 1258
rect 4382 1252 4385 1258
rect 4398 1222 4401 1258
rect 4422 1252 4425 1258
rect 4430 1241 4433 1258
rect 4446 1252 4449 1318
rect 4466 1268 4470 1271
rect 4462 1252 4465 1258
rect 4478 1252 4481 1298
rect 4486 1272 4489 1328
rect 4494 1262 4497 1278
rect 4502 1272 4505 1338
rect 4550 1292 4553 1428
rect 4574 1392 4577 1418
rect 4574 1362 4577 1368
rect 4562 1348 4566 1351
rect 4582 1332 4585 1458
rect 4582 1292 4585 1328
rect 4590 1292 4593 1348
rect 4598 1342 4601 1348
rect 4538 1278 4542 1281
rect 4518 1272 4521 1278
rect 4554 1268 4558 1271
rect 4422 1238 4433 1241
rect 4390 1192 4393 1218
rect 4398 1202 4401 1218
rect 4282 1148 4286 1151
rect 4314 1148 4318 1151
rect 4262 1142 4265 1148
rect 4282 1138 4286 1141
rect 4294 1091 4297 1148
rect 4314 1138 4318 1141
rect 4338 1138 4342 1141
rect 4326 1132 4329 1138
rect 4334 1102 4337 1118
rect 4286 1088 4297 1091
rect 4258 1068 4262 1071
rect 4270 1062 4273 1088
rect 4278 1072 4281 1078
rect 4214 1028 4225 1031
rect 4138 958 4142 961
rect 4150 961 4153 1018
rect 4150 958 4161 961
rect 4130 948 4134 951
rect 4118 932 4121 938
rect 4126 882 4129 948
rect 4150 942 4153 948
rect 4142 881 4145 918
rect 4142 878 4150 881
rect 4126 872 4129 878
rect 4110 862 4113 868
rect 4126 862 4129 868
rect 4070 858 4081 861
rect 4090 858 4094 861
rect 4078 852 4081 858
rect 4066 848 4070 851
rect 4134 802 4137 868
rect 4158 862 4161 958
rect 4182 952 4185 1018
rect 4170 948 4174 951
rect 4190 942 4193 948
rect 4206 932 4209 1008
rect 4202 918 4206 921
rect 4174 882 4177 888
rect 4214 882 4217 1028
rect 4246 1002 4249 1048
rect 4286 1032 4289 1088
rect 4294 1072 4297 1078
rect 4302 1072 4305 1098
rect 4350 1092 4353 1148
rect 4326 1062 4329 1088
rect 4338 1078 4345 1081
rect 4342 1072 4345 1078
rect 4334 1062 4337 1068
rect 4338 1058 4345 1061
rect 4310 1052 4313 1058
rect 4298 1028 4302 1031
rect 4254 1002 4257 1018
rect 4230 942 4233 978
rect 4262 962 4265 1028
rect 4286 962 4289 968
rect 4318 962 4321 1018
rect 4242 948 4246 951
rect 4242 938 4246 941
rect 4186 878 4190 881
rect 4202 878 4209 881
rect 4206 872 4209 878
rect 4170 868 4174 871
rect 4154 848 4158 851
rect 4006 762 4009 768
rect 4014 752 4017 758
rect 4046 752 4049 788
rect 4166 782 4169 868
rect 4190 852 4193 868
rect 4214 862 4217 878
rect 4222 872 4225 918
rect 4230 862 4233 918
rect 4238 882 4241 898
rect 4246 882 4249 888
rect 4198 842 4201 858
rect 4214 842 4217 848
rect 4222 842 4225 848
rect 4238 832 4241 868
rect 4246 842 4249 848
rect 4254 822 4257 948
rect 4262 902 4265 958
rect 4294 952 4297 958
rect 4326 952 4329 1058
rect 4286 942 4289 948
rect 4314 938 4318 941
rect 4302 932 4305 938
rect 4326 932 4329 948
rect 4334 912 4337 1048
rect 4342 952 4345 1058
rect 4350 1022 4353 1058
rect 4358 962 4361 1148
rect 4366 1062 4369 1068
rect 4382 1062 4385 1108
rect 4390 1052 4393 1158
rect 4398 1152 4401 1198
rect 4406 1142 4409 1238
rect 4422 1192 4425 1238
rect 4430 1152 4433 1158
rect 4446 1152 4449 1178
rect 4478 1162 4481 1248
rect 4494 1242 4497 1248
rect 4502 1222 4505 1268
rect 4514 1248 4518 1251
rect 4510 1192 4513 1208
rect 4534 1192 4537 1258
rect 4542 1242 4545 1268
rect 4562 1258 4566 1261
rect 4530 1158 4534 1161
rect 4462 1152 4465 1158
rect 4398 1112 4401 1118
rect 4422 1082 4425 1148
rect 4430 1102 4433 1118
rect 4410 1078 4414 1081
rect 4398 1052 4401 1068
rect 4422 1062 4425 1068
rect 4438 1062 4441 1138
rect 4406 1052 4409 1058
rect 4446 1052 4449 1148
rect 4490 1138 4494 1141
rect 4454 1092 4457 1138
rect 4478 1082 4481 1138
rect 4486 1092 4489 1118
rect 4502 1112 4505 1138
rect 4454 1072 4457 1078
rect 4478 1072 4481 1078
rect 4462 1062 4465 1068
rect 4486 1062 4489 1068
rect 4494 1062 4497 1098
rect 4518 1072 4521 1158
rect 4434 1048 4438 1051
rect 4454 1051 4457 1058
rect 4454 1048 4465 1051
rect 4462 1042 4465 1048
rect 4382 1032 4385 1038
rect 4374 1012 4377 1018
rect 4382 1001 4385 1008
rect 4374 998 4385 1001
rect 4374 962 4377 998
rect 4386 988 4390 991
rect 4398 962 4401 968
rect 4354 948 4358 951
rect 4270 872 4273 898
rect 4278 872 4281 878
rect 4294 862 4297 868
rect 4266 858 4270 861
rect 4198 772 4201 778
rect 4110 762 4113 768
rect 3954 748 3958 751
rect 4002 748 4006 751
rect 4022 742 4025 748
rect 4030 742 4033 748
rect 4110 742 4113 748
rect 3914 738 3918 741
rect 4066 738 4070 741
rect 4146 738 4150 741
rect 3926 732 3929 738
rect 4050 728 4054 731
rect 3902 682 3905 718
rect 3950 672 3953 678
rect 3890 668 3894 671
rect 3802 658 3809 661
rect 3814 652 3817 658
rect 3842 648 3846 651
rect 3822 622 3825 648
rect 3862 642 3865 668
rect 3758 588 3769 591
rect 3758 562 3761 588
rect 3854 582 3857 618
rect 3870 602 3873 658
rect 3902 642 3905 648
rect 3922 638 3926 641
rect 3934 612 3937 658
rect 3930 578 3934 581
rect 3842 568 3849 571
rect 3838 562 3841 568
rect 3758 512 3761 558
rect 3766 552 3769 558
rect 3782 542 3785 548
rect 3790 542 3793 558
rect 3810 548 3814 551
rect 3798 532 3801 548
rect 3806 512 3809 548
rect 3830 542 3833 558
rect 3818 538 3822 541
rect 3838 531 3841 548
rect 3846 542 3849 568
rect 3854 562 3857 568
rect 3866 558 3870 561
rect 3878 552 3881 578
rect 3858 548 3862 551
rect 3834 528 3841 531
rect 3806 482 3809 488
rect 3758 462 3761 478
rect 3814 472 3817 478
rect 3714 458 3718 461
rect 3746 458 3750 461
rect 3822 461 3825 518
rect 3854 492 3857 538
rect 3890 528 3894 531
rect 3878 521 3881 528
rect 3878 518 3889 521
rect 3886 492 3889 518
rect 3878 482 3881 488
rect 3814 458 3825 461
rect 3858 478 3862 481
rect 3830 462 3833 478
rect 3842 468 3846 471
rect 3870 471 3873 478
rect 3870 468 3878 471
rect 3882 468 3886 471
rect 3854 462 3857 468
rect 3782 452 3785 458
rect 3798 442 3801 458
rect 3718 422 3721 428
rect 3770 418 3774 421
rect 3662 378 3673 381
rect 3530 358 3534 361
rect 3518 352 3521 358
rect 3510 338 3521 341
rect 3502 332 3505 338
rect 3430 278 3441 281
rect 3406 252 3409 268
rect 3414 242 3417 268
rect 3422 251 3425 268
rect 3430 262 3433 278
rect 3422 248 3430 251
rect 3438 251 3441 268
rect 3446 261 3449 278
rect 3470 272 3473 278
rect 3494 272 3497 278
rect 3502 272 3505 328
rect 3510 292 3513 318
rect 3518 292 3521 338
rect 3542 321 3545 338
rect 3550 332 3553 348
rect 3558 342 3561 358
rect 3542 318 3553 321
rect 3526 282 3529 288
rect 3458 268 3462 271
rect 3446 258 3454 261
rect 3434 248 3441 251
rect 3470 242 3473 268
rect 3510 248 3518 251
rect 3534 251 3537 318
rect 3550 282 3553 318
rect 3566 312 3569 318
rect 3574 302 3577 328
rect 3566 292 3569 298
rect 3542 262 3545 278
rect 3550 272 3553 278
rect 3530 248 3537 251
rect 3438 202 3441 238
rect 3486 222 3489 248
rect 3510 222 3513 248
rect 3374 92 3377 118
rect 3382 112 3385 148
rect 3322 78 3326 81
rect 3346 78 3350 81
rect 3310 68 3318 71
rect 3366 62 3369 68
rect 3382 62 3385 108
rect 3390 72 3393 78
rect 3398 72 3401 88
rect 3342 52 3345 58
rect 3414 52 3417 148
rect 3422 142 3425 148
rect 3430 102 3433 148
rect 3438 112 3441 138
rect 3454 132 3457 158
rect 3486 152 3489 198
rect 3462 142 3465 148
rect 3478 142 3481 148
rect 3438 82 3441 108
rect 3446 92 3449 98
rect 3470 92 3473 118
rect 3494 92 3497 198
rect 3518 162 3521 208
rect 3550 182 3553 268
rect 3558 242 3561 268
rect 3574 232 3577 298
rect 3590 262 3593 338
rect 3598 272 3601 278
rect 3606 262 3609 368
rect 3634 358 3638 361
rect 3622 332 3625 358
rect 3630 352 3633 358
rect 3654 352 3657 358
rect 3618 288 3622 291
rect 3622 251 3625 258
rect 3594 248 3625 251
rect 3630 252 3633 318
rect 3646 282 3649 338
rect 3662 292 3665 328
rect 3654 272 3657 278
rect 3662 262 3665 278
rect 3650 248 3662 251
rect 3568 203 3570 207
rect 3574 203 3577 207
rect 3581 203 3584 207
rect 3590 152 3593 238
rect 3522 148 3526 151
rect 3510 142 3513 148
rect 3534 142 3537 148
rect 3534 132 3537 138
rect 3518 112 3521 118
rect 3526 92 3529 108
rect 3542 92 3545 138
rect 3550 132 3553 148
rect 3574 142 3577 148
rect 3562 128 3566 131
rect 3606 122 3609 128
rect 3590 92 3593 98
rect 3614 92 3617 238
rect 3622 192 3625 198
rect 3422 72 3425 78
rect 3478 72 3481 78
rect 3550 72 3553 78
rect 3598 72 3601 88
rect 3622 82 3625 148
rect 3630 132 3633 178
rect 3642 158 3646 161
rect 3654 82 3657 178
rect 3662 152 3665 218
rect 3670 192 3673 378
rect 3678 352 3681 398
rect 3678 332 3681 338
rect 3686 332 3689 368
rect 3718 362 3721 418
rect 3814 412 3817 458
rect 3894 452 3897 498
rect 3902 492 3905 558
rect 3950 552 3953 658
rect 3958 562 3961 668
rect 3966 562 3969 718
rect 4102 712 4105 738
rect 4130 728 4134 731
rect 4158 722 4161 748
rect 4166 732 4169 758
rect 4186 748 4190 751
rect 4080 703 4082 707
rect 4086 703 4089 707
rect 4093 703 4096 707
rect 3994 688 3998 691
rect 4030 672 4033 678
rect 3982 662 3985 668
rect 4002 658 4006 661
rect 4014 652 4017 668
rect 4038 662 4041 668
rect 4038 652 4041 658
rect 4046 652 4049 678
rect 4070 672 4073 678
rect 4110 672 4113 698
rect 4106 668 4110 671
rect 4058 658 4062 661
rect 4050 648 4057 651
rect 3974 612 3977 648
rect 3998 622 4001 648
rect 4018 618 4022 621
rect 4014 592 4017 608
rect 3910 502 3913 548
rect 3934 542 3937 548
rect 3950 542 3953 548
rect 3922 538 3929 541
rect 3926 532 3929 538
rect 3942 531 3945 538
rect 3934 528 3945 531
rect 3918 481 3921 528
rect 3934 522 3937 528
rect 3950 512 3953 518
rect 3914 478 3921 481
rect 3910 472 3913 478
rect 3918 462 3921 468
rect 3942 462 3945 508
rect 3954 458 3958 461
rect 3942 452 3945 458
rect 3950 452 3953 458
rect 3822 442 3825 448
rect 3934 442 3937 448
rect 3958 442 3961 448
rect 3842 438 3846 441
rect 3734 362 3737 408
rect 3830 392 3833 438
rect 3926 372 3929 418
rect 3934 392 3937 408
rect 3806 362 3809 368
rect 3842 358 3849 361
rect 3722 348 3726 351
rect 3738 348 3742 351
rect 3750 348 3758 351
rect 3694 342 3697 348
rect 3694 292 3697 298
rect 3702 282 3705 348
rect 3710 332 3713 338
rect 3742 332 3745 338
rect 3710 292 3713 308
rect 3750 302 3753 348
rect 3766 342 3769 358
rect 3750 292 3753 298
rect 3686 272 3689 278
rect 3678 262 3681 268
rect 3718 262 3721 278
rect 3738 268 3742 271
rect 3706 258 3710 261
rect 3722 258 3726 261
rect 3678 192 3681 208
rect 3710 162 3713 248
rect 3734 192 3737 258
rect 3698 158 3702 161
rect 3686 152 3689 158
rect 3734 152 3737 188
rect 3698 148 3702 151
rect 3718 142 3721 148
rect 3710 132 3713 138
rect 3670 92 3673 98
rect 3506 68 3510 71
rect 3626 68 3630 71
rect 3674 68 3678 71
rect 3426 58 3430 61
rect 3438 52 3441 68
rect 3454 62 3457 68
rect 3462 62 3465 68
rect 3478 62 3481 68
rect 3638 62 3641 68
rect 3498 58 3502 61
rect 3530 58 3534 61
rect 3526 52 3529 58
rect 3574 52 3577 58
rect 2802 48 2809 51
rect 2906 48 2910 51
rect 2954 48 2958 51
rect 2970 48 2974 51
rect 3050 48 3054 51
rect 3122 48 3126 51
rect 3178 48 3182 51
rect 3218 48 3222 51
rect 3242 48 3246 51
rect 3290 48 3294 51
rect 3302 48 3310 51
rect 3402 48 3406 51
rect 3610 48 3614 51
rect 2582 41 2585 48
rect 2558 38 2585 41
rect 3014 42 3017 48
rect 3302 42 3305 48
rect 3414 42 3417 48
rect 3654 42 3657 58
rect 3114 28 3118 31
rect 3338 28 3342 31
rect 1382 -22 1393 -19
rect 3082 18 3086 21
rect 1398 -18 1401 18
rect 1398 -22 1402 -18
rect 1414 -19 1418 -18
rect 1422 -19 1425 18
rect 1520 3 1522 7
rect 1526 3 1529 7
rect 1533 3 1536 7
rect 1414 -22 1425 -19
rect 1550 -19 1554 -18
rect 1558 -19 1561 18
rect 1550 -22 1561 -19
rect 1574 -19 1578 -18
rect 1582 -19 1585 18
rect 3678 12 3681 68
rect 3694 52 3697 118
rect 3702 72 3705 78
rect 3718 62 3721 68
rect 3706 58 3710 61
rect 3698 48 3702 51
rect 3726 22 3729 138
rect 3734 92 3737 138
rect 3742 62 3745 228
rect 3758 192 3761 268
rect 3766 192 3769 338
rect 3774 332 3777 348
rect 3774 212 3777 258
rect 3782 242 3785 338
rect 3814 332 3817 348
rect 3838 342 3841 348
rect 3790 252 3793 328
rect 3814 312 3817 328
rect 3822 292 3825 318
rect 3830 272 3833 288
rect 3838 272 3841 328
rect 3846 292 3849 358
rect 3942 352 3945 408
rect 3950 402 3953 418
rect 3890 348 3894 351
rect 3854 332 3857 348
rect 3854 282 3857 318
rect 3862 292 3865 338
rect 3842 268 3846 271
rect 3858 268 3862 271
rect 3774 152 3777 208
rect 3798 202 3801 268
rect 3830 262 3833 268
rect 3822 252 3825 258
rect 3858 248 3862 251
rect 3870 242 3873 328
rect 3878 262 3881 298
rect 3886 272 3889 348
rect 3950 342 3953 348
rect 3958 342 3961 408
rect 3966 401 3969 558
rect 4054 552 4057 648
rect 4062 592 4065 618
rect 4062 552 4065 558
rect 3986 548 3990 551
rect 4042 548 4046 551
rect 4082 548 4086 551
rect 3974 532 3977 538
rect 3986 528 3990 531
rect 3998 522 4001 548
rect 3974 452 3977 498
rect 3982 482 3985 488
rect 3990 452 3993 518
rect 4006 502 4009 548
rect 4030 532 4033 548
rect 4054 542 4057 548
rect 4094 542 4097 668
rect 4106 648 4110 651
rect 4118 642 4121 668
rect 4126 662 4129 718
rect 4166 702 4169 728
rect 4158 672 4161 678
rect 4174 672 4177 718
rect 4190 712 4193 738
rect 4206 692 4209 818
rect 4238 792 4241 808
rect 4214 762 4217 778
rect 4262 772 4265 778
rect 4234 768 4238 771
rect 4214 752 4217 758
rect 4222 752 4225 768
rect 4242 758 4246 761
rect 4238 692 4241 728
rect 4246 692 4249 738
rect 4254 682 4257 688
rect 4262 682 4265 748
rect 4142 668 4150 671
rect 4186 668 4190 671
rect 4126 552 4129 618
rect 4142 612 4145 668
rect 4186 658 4190 661
rect 4150 582 4153 658
rect 4166 612 4169 658
rect 4198 651 4201 678
rect 4186 648 4201 651
rect 4206 642 4209 678
rect 4234 668 4238 671
rect 4258 668 4262 671
rect 4114 548 4118 551
rect 4042 538 4046 541
rect 4002 488 4006 491
rect 4022 472 4025 528
rect 4054 492 4057 538
rect 4062 492 4065 498
rect 4058 478 4062 481
rect 4070 481 4073 538
rect 4126 532 4129 538
rect 4134 532 4137 558
rect 4154 548 4158 551
rect 4166 542 4169 608
rect 4182 542 4185 608
rect 4142 532 4145 538
rect 4162 528 4166 531
rect 4080 503 4082 507
rect 4086 503 4089 507
rect 4093 503 4096 507
rect 4102 482 4105 488
rect 4070 478 4081 481
rect 4010 468 4014 471
rect 4050 468 4054 471
rect 3998 462 4001 468
rect 4038 462 4041 468
rect 4022 442 4025 448
rect 3966 398 3974 401
rect 4006 362 4009 398
rect 4022 372 4025 438
rect 4038 402 4041 418
rect 4046 391 4049 398
rect 4042 388 4049 391
rect 4070 382 4073 468
rect 3966 352 3969 358
rect 3994 348 3998 351
rect 3942 332 3945 338
rect 3914 328 3918 331
rect 3910 322 3913 328
rect 3894 282 3897 288
rect 3910 262 3913 308
rect 3966 292 3969 348
rect 3974 342 3977 348
rect 3982 342 3985 348
rect 3990 331 3993 338
rect 3986 328 3993 331
rect 4006 332 4009 338
rect 3982 292 3985 328
rect 3990 322 3993 328
rect 3938 278 3942 281
rect 3942 262 3945 268
rect 3950 262 3953 288
rect 3958 272 3961 278
rect 3930 258 3934 261
rect 3966 252 3969 278
rect 3998 272 4001 308
rect 3974 242 3977 248
rect 3754 138 3758 141
rect 3782 132 3785 188
rect 3810 168 3814 171
rect 3794 158 3798 161
rect 3822 152 3825 158
rect 3838 152 3841 238
rect 3854 162 3857 198
rect 3862 192 3865 218
rect 3794 148 3798 151
rect 3830 142 3833 148
rect 3838 142 3841 148
rect 3750 112 3753 128
rect 3754 78 3758 81
rect 3766 72 3769 78
rect 3774 32 3777 128
rect 3782 112 3785 128
rect 3798 112 3801 138
rect 3846 132 3849 158
rect 3870 152 3873 168
rect 3858 148 3862 151
rect 3890 148 3894 151
rect 3890 138 3894 141
rect 3902 112 3905 218
rect 3910 192 3913 208
rect 3958 192 3961 218
rect 3938 178 3942 181
rect 3990 172 3993 268
rect 4014 262 4017 358
rect 4042 348 4046 351
rect 4022 342 4025 348
rect 4054 341 4057 358
rect 4062 352 4065 368
rect 4054 338 4062 341
rect 4078 341 4081 478
rect 4110 472 4113 528
rect 4174 502 4177 518
rect 4122 478 4126 481
rect 4150 472 4153 498
rect 4118 462 4121 468
rect 4142 462 4145 468
rect 4118 392 4121 458
rect 4158 452 4161 498
rect 4174 462 4177 488
rect 4190 472 4193 588
rect 4198 552 4201 568
rect 4206 542 4209 638
rect 4214 602 4217 668
rect 4278 662 4281 858
rect 4302 852 4305 878
rect 4326 872 4329 878
rect 4334 872 4337 908
rect 4374 902 4377 918
rect 4370 868 4374 871
rect 4318 862 4321 868
rect 4382 861 4385 958
rect 4414 952 4417 958
rect 4390 912 4393 948
rect 4430 942 4433 958
rect 4438 952 4441 1018
rect 4454 992 4457 1008
rect 4458 968 4462 971
rect 4446 962 4449 968
rect 4470 962 4473 978
rect 4474 958 4478 961
rect 4442 948 4449 951
rect 4410 928 4414 931
rect 4414 872 4417 898
rect 4446 892 4449 948
rect 4486 951 4489 1058
rect 4510 1052 4513 1058
rect 4494 992 4497 1018
rect 4510 952 4513 958
rect 4486 948 4494 951
rect 4454 942 4457 948
rect 4478 942 4481 948
rect 4478 892 4481 908
rect 4486 902 4489 948
rect 4502 932 4505 938
rect 4518 902 4521 1068
rect 4526 1052 4529 1148
rect 4550 1132 4553 1148
rect 4558 1142 4561 1158
rect 4542 1128 4550 1131
rect 4542 1072 4545 1128
rect 4558 1092 4561 1128
rect 4538 1068 4542 1071
rect 4538 1058 4542 1061
rect 4526 1042 4529 1048
rect 4530 968 4534 971
rect 4526 922 4529 928
rect 4482 878 4486 881
rect 4434 868 4438 871
rect 4374 858 4385 861
rect 4410 858 4414 861
rect 4286 792 4289 818
rect 4294 762 4297 838
rect 4326 832 4329 858
rect 4322 788 4326 791
rect 4350 772 4353 818
rect 4374 812 4377 858
rect 4386 848 4390 851
rect 4422 842 4425 868
rect 4438 822 4441 858
rect 4454 852 4457 868
rect 4502 862 4505 868
rect 4518 862 4521 878
rect 4466 858 4470 861
rect 4510 852 4513 858
rect 4430 792 4433 818
rect 4382 772 4385 778
rect 4414 762 4417 768
rect 4286 742 4289 748
rect 4294 732 4297 758
rect 4286 682 4289 688
rect 4294 682 4297 718
rect 4310 702 4313 748
rect 4318 682 4321 738
rect 4342 732 4345 748
rect 4350 732 4353 758
rect 4358 742 4361 748
rect 4406 742 4409 748
rect 4378 738 4382 741
rect 4394 738 4398 741
rect 4398 732 4401 738
rect 4374 711 4377 728
rect 4382 722 4385 728
rect 4374 708 4385 711
rect 4374 702 4377 708
rect 4366 682 4369 688
rect 4294 672 4297 678
rect 4282 658 4286 661
rect 4222 582 4225 658
rect 4230 622 4233 658
rect 4246 592 4249 648
rect 4270 642 4273 658
rect 4302 592 4305 678
rect 4362 668 4366 671
rect 4342 662 4345 668
rect 4374 662 4377 668
rect 4310 642 4313 658
rect 4318 652 4321 658
rect 4198 532 4201 538
rect 4222 532 4225 578
rect 4198 462 4201 478
rect 4214 462 4217 518
rect 4130 448 4137 451
rect 4202 448 4206 451
rect 4074 338 4081 341
rect 4022 292 4025 308
rect 4030 302 4033 338
rect 4030 272 4033 298
rect 4038 262 4041 288
rect 4002 258 4006 261
rect 3934 151 3937 158
rect 3934 148 3942 151
rect 3910 132 3913 138
rect 3866 78 3870 81
rect 3790 72 3793 78
rect 3878 72 3881 88
rect 3842 68 3846 71
rect 3862 62 3865 68
rect 3886 62 3889 108
rect 3918 82 3921 138
rect 3926 132 3929 148
rect 3942 142 3945 148
rect 3950 142 3953 158
rect 4006 152 4009 168
rect 3982 142 3985 148
rect 4014 142 4017 258
rect 4022 222 4025 248
rect 4046 192 4049 338
rect 4074 328 4078 331
rect 4090 328 4094 331
rect 4080 303 4082 307
rect 4086 303 4089 307
rect 4093 303 4096 307
rect 4054 282 4057 288
rect 4054 212 4057 258
rect 4062 242 4065 268
rect 4070 262 4073 298
rect 4102 292 4105 338
rect 4110 322 4113 358
rect 4118 352 4121 358
rect 4126 302 4129 368
rect 4134 331 4137 448
rect 4174 412 4177 418
rect 4146 368 4150 371
rect 4142 342 4145 348
rect 4166 342 4169 368
rect 4190 352 4193 438
rect 4214 412 4217 448
rect 4206 392 4209 398
rect 4230 382 4233 558
rect 4238 492 4241 578
rect 4302 572 4305 588
rect 4246 532 4249 548
rect 4254 542 4257 548
rect 4262 522 4265 548
rect 4278 532 4281 568
rect 4286 542 4289 548
rect 4294 532 4297 548
rect 4246 472 4249 518
rect 4254 472 4257 478
rect 4270 472 4273 518
rect 4294 512 4297 528
rect 4294 462 4297 508
rect 4310 492 4313 638
rect 4318 592 4321 648
rect 4350 642 4353 648
rect 4334 632 4337 638
rect 4326 582 4329 618
rect 4350 592 4353 628
rect 4382 612 4385 708
rect 4414 692 4417 698
rect 4406 662 4409 668
rect 4422 662 4425 768
rect 4430 732 4433 748
rect 4438 742 4441 818
rect 4454 762 4457 848
rect 4518 792 4521 838
rect 4534 832 4537 858
rect 4542 772 4545 1038
rect 4550 1032 4553 1068
rect 4566 992 4569 1168
rect 4574 1092 4577 1148
rect 4582 1142 4585 1188
rect 4598 1172 4601 1258
rect 4590 1070 4593 1118
rect 4598 1032 4601 1068
rect 4554 958 4558 961
rect 4562 948 4566 951
rect 4550 932 4553 938
rect 4574 922 4577 968
rect 4550 882 4553 888
rect 4562 878 4566 881
rect 4582 872 4585 878
rect 4550 868 4558 871
rect 4470 762 4473 768
rect 4446 721 4449 738
rect 4438 718 4449 721
rect 4398 622 4401 658
rect 4390 572 4393 578
rect 4406 572 4409 658
rect 4414 632 4417 648
rect 4430 642 4433 658
rect 4438 652 4441 718
rect 4454 681 4457 748
rect 4470 742 4473 748
rect 4478 731 4481 748
rect 4470 728 4481 731
rect 4450 678 4457 681
rect 4446 672 4449 678
rect 4462 652 4465 708
rect 4450 648 4454 651
rect 4326 561 4329 568
rect 4318 558 4329 561
rect 4374 558 4393 561
rect 4318 552 4321 558
rect 4374 552 4377 558
rect 4318 532 4321 538
rect 4326 482 4329 548
rect 4342 482 4345 528
rect 4366 512 4369 538
rect 4374 532 4377 538
rect 4382 521 4385 548
rect 4374 518 4385 521
rect 4374 492 4377 518
rect 4390 492 4393 558
rect 4406 552 4409 558
rect 4430 552 4433 638
rect 4470 631 4473 728
rect 4478 692 4481 718
rect 4486 712 4489 738
rect 4498 728 4502 731
rect 4510 722 4513 738
rect 4478 642 4481 648
rect 4470 628 4481 631
rect 4438 552 4441 558
rect 4454 552 4457 588
rect 4462 552 4465 568
rect 4414 502 4417 538
rect 4442 518 4446 521
rect 4454 511 4457 548
rect 4470 542 4473 618
rect 4478 592 4481 628
rect 4486 592 4489 658
rect 4494 652 4497 668
rect 4506 658 4510 661
rect 4494 642 4497 648
rect 4478 542 4481 588
rect 4502 552 4505 578
rect 4518 552 4521 768
rect 4538 748 4542 751
rect 4526 692 4529 728
rect 4534 722 4537 738
rect 4542 732 4545 738
rect 4542 692 4545 708
rect 4550 702 4553 868
rect 4574 822 4577 858
rect 4590 842 4593 848
rect 4570 718 4574 721
rect 4598 712 4601 738
rect 4570 678 4574 681
rect 4530 668 4534 671
rect 4542 658 4550 661
rect 4526 652 4529 658
rect 4526 562 4529 648
rect 4542 592 4545 658
rect 4558 602 4561 668
rect 4578 618 4582 621
rect 4574 592 4577 608
rect 4550 552 4553 568
rect 4558 562 4561 568
rect 4514 548 4518 551
rect 4578 548 4582 551
rect 4462 532 4465 538
rect 4446 508 4457 511
rect 4470 512 4473 538
rect 4398 492 4401 498
rect 4430 492 4433 508
rect 4446 492 4449 508
rect 4362 488 4366 491
rect 4382 482 4385 488
rect 4346 478 4350 481
rect 4302 462 4305 468
rect 4238 452 4241 458
rect 4278 452 4281 458
rect 4238 362 4241 418
rect 4254 352 4257 448
rect 4262 392 4265 408
rect 4278 392 4281 448
rect 4310 422 4313 478
rect 4414 472 4417 488
rect 4462 482 4465 488
rect 4338 468 4345 471
rect 4322 458 4326 461
rect 4318 442 4321 448
rect 4330 428 4334 431
rect 4342 392 4345 468
rect 4402 468 4406 471
rect 4350 462 4353 468
rect 4494 462 4497 538
rect 4510 532 4513 538
rect 4502 482 4505 488
rect 4514 478 4518 481
rect 4518 462 4521 468
rect 4490 458 4494 461
rect 4366 442 4369 458
rect 4390 412 4393 448
rect 4322 358 4326 361
rect 4302 352 4305 358
rect 4242 348 4246 351
rect 4282 348 4286 351
rect 4346 348 4350 351
rect 4378 348 4382 351
rect 4134 328 4145 331
rect 4110 282 4113 288
rect 4114 268 4118 271
rect 4062 212 4065 238
rect 4026 148 4030 151
rect 3970 138 3974 141
rect 3994 138 3998 141
rect 4026 138 4030 141
rect 4046 132 4049 178
rect 4054 162 4057 188
rect 4078 152 4081 248
rect 4086 202 4089 268
rect 4126 262 4129 298
rect 4142 292 4145 328
rect 4134 262 4137 268
rect 4086 172 4089 198
rect 4102 192 4105 258
rect 4110 162 4113 258
rect 4150 232 4153 278
rect 4158 272 4161 328
rect 4158 242 4161 268
rect 4166 252 4169 258
rect 4118 162 4121 188
rect 4094 142 4097 158
rect 4118 142 4121 148
rect 4126 142 4129 228
rect 4142 172 4145 188
rect 4134 152 4137 158
rect 4154 148 4158 151
rect 4166 142 4169 228
rect 4174 162 4177 348
rect 4190 342 4193 348
rect 4222 342 4225 348
rect 4182 292 4185 328
rect 4190 322 4193 328
rect 4198 322 4201 338
rect 4230 332 4233 348
rect 4270 342 4273 348
rect 4310 342 4313 348
rect 4246 332 4249 338
rect 4210 328 4214 331
rect 4290 328 4294 331
rect 4198 292 4201 308
rect 4246 292 4249 308
rect 4186 278 4190 281
rect 4206 272 4209 278
rect 4222 272 4225 278
rect 4226 258 4230 261
rect 4182 232 4185 248
rect 4214 212 4217 258
rect 4190 152 4193 158
rect 4198 152 4201 158
rect 4206 142 4209 148
rect 4154 138 4158 141
rect 3954 128 3958 131
rect 3894 72 3897 78
rect 3926 72 3929 78
rect 3958 72 3961 78
rect 3914 68 3918 71
rect 3982 62 3985 128
rect 4014 92 4017 128
rect 4070 102 4073 138
rect 4110 128 4118 131
rect 4080 103 4082 107
rect 4086 103 4089 107
rect 4093 103 4096 107
rect 4034 68 4038 71
rect 3802 58 3806 61
rect 3906 58 3910 61
rect 3922 58 3926 61
rect 3938 58 3942 61
rect 3782 52 3785 58
rect 3810 48 3814 51
rect 3826 48 3830 51
rect 3798 42 3801 48
rect 3846 32 3849 58
rect 3854 52 3857 58
rect 3938 48 3942 51
rect 3950 22 3953 58
rect 3990 52 3993 68
rect 3998 62 4001 68
rect 4034 58 4038 61
rect 3970 48 3974 51
rect 4046 42 4049 98
rect 4102 92 4105 108
rect 4070 82 4073 88
rect 4110 82 4113 128
rect 4190 112 4193 138
rect 4214 131 4217 208
rect 4222 192 4225 198
rect 4238 192 4241 238
rect 4246 202 4249 248
rect 4254 242 4257 268
rect 4262 252 4265 328
rect 4270 262 4273 328
rect 4286 292 4289 318
rect 4290 288 4294 291
rect 4254 152 4257 208
rect 4278 152 4281 248
rect 4294 152 4297 168
rect 4302 162 4305 248
rect 4310 192 4313 328
rect 4318 292 4321 348
rect 4390 341 4393 348
rect 4382 338 4393 341
rect 4350 302 4353 338
rect 4358 322 4361 328
rect 4342 292 4345 298
rect 4350 292 4353 298
rect 4358 292 4361 318
rect 4374 312 4377 338
rect 4382 292 4385 338
rect 4390 332 4393 338
rect 4398 292 4401 458
rect 4426 448 4430 451
rect 4438 442 4441 448
rect 4470 392 4473 458
rect 4478 442 4481 458
rect 4526 451 4529 548
rect 4578 538 4582 541
rect 4554 528 4558 531
rect 4534 472 4537 528
rect 4542 482 4545 518
rect 4550 492 4553 498
rect 4574 472 4577 478
rect 4534 462 4537 468
rect 4558 452 4561 458
rect 4522 448 4529 451
rect 4538 448 4542 451
rect 4518 412 4521 448
rect 4558 392 4561 438
rect 4438 362 4441 368
rect 4502 362 4505 368
rect 4570 358 4574 361
rect 4410 348 4414 351
rect 4530 348 4534 351
rect 4414 312 4417 338
rect 4422 332 4425 348
rect 4446 332 4449 348
rect 4494 342 4497 348
rect 4550 342 4553 348
rect 4478 332 4481 338
rect 4490 328 4494 331
rect 4518 302 4521 318
rect 4318 262 4321 268
rect 4350 262 4353 268
rect 4402 258 4406 261
rect 4326 162 4329 258
rect 4342 192 4345 218
rect 4322 158 4326 161
rect 4234 148 4238 151
rect 4350 151 4353 258
rect 4346 148 4353 151
rect 4358 252 4361 258
rect 4382 252 4385 258
rect 4390 252 4393 258
rect 4414 251 4417 298
rect 4446 272 4449 298
rect 4422 262 4425 268
rect 4454 262 4457 278
rect 4470 262 4473 298
rect 4478 262 4481 288
rect 4518 282 4521 288
rect 4506 278 4510 281
rect 4486 272 4489 278
rect 4506 268 4510 271
rect 4534 262 4537 338
rect 4542 332 4545 338
rect 4550 271 4553 338
rect 4546 268 4553 271
rect 4414 248 4422 251
rect 4358 152 4361 248
rect 4406 222 4409 238
rect 4414 192 4417 228
rect 4366 162 4369 168
rect 4382 162 4385 178
rect 4438 152 4441 258
rect 4454 192 4457 238
rect 4214 128 4222 131
rect 4230 112 4233 138
rect 4238 112 4241 148
rect 4266 138 4270 141
rect 4290 138 4294 141
rect 4270 112 4273 128
rect 4302 102 4305 128
rect 4318 122 4321 148
rect 4342 142 4345 148
rect 4350 131 4353 138
rect 4346 128 4353 131
rect 4358 132 4361 138
rect 4210 88 4214 91
rect 4158 72 4161 88
rect 4286 82 4289 88
rect 4310 82 4313 88
rect 4326 82 4329 108
rect 4366 82 4369 148
rect 4398 142 4401 148
rect 4414 132 4417 138
rect 4410 128 4414 131
rect 4422 122 4425 148
rect 4446 142 4449 188
rect 4470 162 4473 218
rect 4494 192 4497 218
rect 4454 152 4457 158
rect 4470 142 4473 148
rect 4434 128 4438 131
rect 4478 112 4481 138
rect 4338 78 4342 81
rect 4382 78 4390 81
rect 4190 72 4193 78
rect 4058 68 4062 71
rect 4122 68 4126 71
rect 4178 68 4182 71
rect 4246 62 4249 78
rect 4258 68 4262 71
rect 4130 58 4134 61
rect 4154 58 4158 61
rect 4046 32 4049 38
rect 4054 32 4057 58
rect 4070 52 4073 58
rect 4182 52 4185 58
rect 4278 52 4281 68
rect 4294 62 4297 78
rect 4374 72 4377 78
rect 4322 68 4326 71
rect 4366 62 4369 68
rect 4342 52 4345 58
rect 4226 48 4230 51
rect 4374 42 4377 58
rect 4382 52 4385 78
rect 4394 68 4398 71
rect 4418 58 4422 61
rect 4406 42 4409 58
rect 4430 52 4433 98
rect 4446 72 4449 78
rect 4454 72 4457 88
rect 4474 78 4478 81
rect 4442 68 4446 71
rect 4478 62 4481 68
rect 4470 52 4473 58
rect 4494 52 4497 58
rect 4502 52 4505 218
rect 4518 212 4521 258
rect 4518 192 4521 208
rect 4542 202 4545 258
rect 4558 192 4561 308
rect 4566 292 4569 348
rect 4510 162 4513 168
rect 4542 152 4545 158
rect 4514 148 4518 151
rect 4530 128 4534 131
rect 4526 62 4529 118
rect 4542 92 4545 138
rect 4534 82 4537 88
rect 4554 68 4558 71
rect 4562 58 4566 61
rect 4550 42 4553 58
rect 4578 48 4582 51
rect 4570 38 4574 41
rect 4146 28 4150 31
rect 4490 28 4494 31
rect 4050 18 4054 21
rect 4162 18 4166 21
rect 4262 12 4265 18
rect 2544 3 2546 7
rect 2550 3 2553 7
rect 2557 3 2560 7
rect 3568 3 3570 7
rect 3574 3 3577 7
rect 3581 3 3584 7
rect 1574 -22 1585 -19
<< m3contact >>
rect 30 4358 34 4362
rect 6 4348 10 4352
rect 70 4348 74 4352
rect 110 4348 114 4352
rect 30 4338 34 4342
rect 54 4338 58 4342
rect 30 4268 34 4272
rect 54 4268 58 4272
rect 102 4338 106 4342
rect 498 4403 502 4407
rect 505 4403 509 4407
rect 1522 4403 1526 4407
rect 1529 4403 1533 4407
rect 1998 4398 2002 4402
rect 2546 4403 2550 4407
rect 2553 4403 2557 4407
rect 1582 4378 1586 4382
rect 2022 4378 2026 4382
rect 774 4368 778 4372
rect 1510 4368 1514 4372
rect 190 4358 194 4362
rect 726 4358 730 4362
rect 758 4358 762 4362
rect 798 4358 802 4362
rect 406 4348 410 4352
rect 462 4348 466 4352
rect 542 4348 546 4352
rect 614 4348 618 4352
rect 286 4338 290 4342
rect 358 4338 362 4342
rect 582 4338 586 4342
rect 78 4328 82 4332
rect 190 4328 194 4332
rect 270 4328 274 4332
rect 126 4318 130 4322
rect 46 4258 50 4262
rect 6 4248 10 4252
rect 30 4248 34 4252
rect 6 4148 10 4152
rect 30 4138 34 4142
rect 6 3968 10 3972
rect 38 4018 42 4022
rect 54 4138 58 4142
rect 230 4288 234 4292
rect 110 4268 114 4272
rect 142 4268 146 4272
rect 190 4258 194 4262
rect 134 4178 138 4182
rect 110 4158 114 4162
rect 86 4148 90 4152
rect 70 4018 74 4022
rect 54 3948 58 3952
rect 70 3938 74 3942
rect 206 4248 210 4252
rect 350 4308 354 4312
rect 358 4298 362 4302
rect 350 4278 354 4282
rect 254 4268 258 4272
rect 294 4268 298 4272
rect 406 4298 410 4302
rect 438 4298 442 4302
rect 414 4288 418 4292
rect 382 4278 386 4282
rect 430 4258 434 4262
rect 534 4288 538 4292
rect 454 4278 458 4282
rect 262 4248 266 4252
rect 302 4248 306 4252
rect 374 4248 378 4252
rect 174 4198 178 4202
rect 230 4198 234 4202
rect 174 4158 178 4162
rect 214 4158 218 4162
rect 254 4188 258 4192
rect 254 4168 258 4172
rect 246 4158 250 4162
rect 366 4238 370 4242
rect 270 4208 274 4212
rect 510 4238 514 4242
rect 430 4228 434 4232
rect 454 4228 458 4232
rect 462 4228 466 4232
rect 478 4228 482 4232
rect 446 4198 450 4202
rect 366 4188 370 4192
rect 326 4168 330 4172
rect 318 4158 322 4162
rect 230 4138 234 4142
rect 182 4128 186 4132
rect 198 4128 202 4132
rect 222 4128 226 4132
rect 238 4128 242 4132
rect 270 4138 274 4142
rect 286 4138 290 4142
rect 302 4138 306 4142
rect 310 4138 314 4142
rect 206 4108 210 4112
rect 110 4098 114 4102
rect 142 4098 146 4102
rect 182 4098 186 4102
rect 182 4078 186 4082
rect 182 4068 186 4072
rect 198 4068 202 4072
rect 110 4018 114 4022
rect 46 3928 50 3932
rect 78 3928 82 3932
rect 102 3928 106 3932
rect 94 3878 98 3882
rect 78 3868 82 3872
rect 6 3848 10 3852
rect 30 3758 34 3762
rect 6 3748 10 3752
rect 14 3748 18 3752
rect 30 3738 34 3742
rect 38 3688 42 3692
rect 54 3738 58 3742
rect 86 3728 90 3732
rect 86 3678 90 3682
rect 6 3668 10 3672
rect 54 3658 58 3662
rect 70 3648 74 3652
rect 6 3548 10 3552
rect 62 3548 66 3552
rect 22 3538 26 3542
rect 70 3538 74 3542
rect 222 4088 226 4092
rect 230 4078 234 4082
rect 214 4068 218 4072
rect 286 4128 290 4132
rect 294 4128 298 4132
rect 294 4098 298 4102
rect 190 4058 194 4062
rect 206 4058 210 4062
rect 230 4058 234 4062
rect 238 4058 242 4062
rect 166 3978 170 3982
rect 126 3948 130 3952
rect 206 3948 210 3952
rect 206 3928 210 3932
rect 246 4048 250 4052
rect 254 4018 258 4022
rect 334 4138 338 4142
rect 430 4178 434 4182
rect 382 4158 386 4162
rect 326 4128 330 4132
rect 350 4128 354 4132
rect 398 4128 402 4132
rect 318 4108 322 4112
rect 318 4078 322 4082
rect 310 4068 314 4072
rect 334 4098 338 4102
rect 382 4108 386 4112
rect 350 4088 354 4092
rect 382 4078 386 4082
rect 374 4068 378 4072
rect 342 4048 346 4052
rect 310 4028 314 4032
rect 326 4028 330 4032
rect 270 4008 274 4012
rect 286 4008 290 4012
rect 254 3988 258 3992
rect 270 3968 274 3972
rect 342 4018 346 4022
rect 318 4008 322 4012
rect 262 3948 266 3952
rect 294 3948 298 3952
rect 286 3938 290 3942
rect 294 3938 298 3942
rect 310 3918 314 3922
rect 214 3878 218 3882
rect 334 3958 338 3962
rect 326 3928 330 3932
rect 366 4058 370 4062
rect 358 4048 362 4052
rect 374 4018 378 4022
rect 350 3988 354 3992
rect 350 3978 354 3982
rect 374 3948 378 3952
rect 446 4148 450 4152
rect 430 4118 434 4122
rect 498 4203 502 4207
rect 505 4203 509 4207
rect 446 4088 450 4092
rect 422 4038 426 4042
rect 406 4028 410 4032
rect 390 3968 394 3972
rect 494 4128 498 4132
rect 470 4098 474 4102
rect 590 4328 594 4332
rect 614 4328 618 4332
rect 614 4318 618 4322
rect 638 4348 642 4352
rect 702 4348 706 4352
rect 742 4348 746 4352
rect 654 4338 658 4342
rect 726 4338 730 4342
rect 630 4288 634 4292
rect 670 4318 674 4322
rect 686 4318 690 4322
rect 678 4308 682 4312
rect 646 4288 650 4292
rect 542 4268 546 4272
rect 582 4268 586 4272
rect 614 4268 618 4272
rect 662 4278 666 4282
rect 590 4258 594 4262
rect 582 4238 586 4242
rect 678 4248 682 4252
rect 710 4308 714 4312
rect 670 4238 674 4242
rect 702 4238 706 4242
rect 598 4228 602 4232
rect 630 4228 634 4232
rect 622 4198 626 4202
rect 542 4188 546 4192
rect 694 4188 698 4192
rect 710 4178 714 4182
rect 694 4168 698 4172
rect 558 4158 562 4162
rect 566 4158 570 4162
rect 606 4158 610 4162
rect 534 4108 538 4112
rect 526 4078 530 4082
rect 534 4068 538 4072
rect 478 4058 482 4062
rect 462 4048 466 4052
rect 454 3978 458 3982
rect 446 3968 450 3972
rect 414 3948 418 3952
rect 358 3938 362 3942
rect 398 3938 402 3942
rect 326 3918 330 3922
rect 334 3918 338 3922
rect 374 3928 378 3932
rect 358 3898 362 3902
rect 382 3918 386 3922
rect 158 3858 162 3862
rect 118 3748 122 3752
rect 102 3728 106 3732
rect 118 3728 122 3732
rect 134 3718 138 3722
rect 214 3838 218 3842
rect 302 3848 306 3852
rect 238 3798 242 3802
rect 270 3798 274 3802
rect 334 3866 338 3870
rect 366 3868 370 3872
rect 414 3908 418 3912
rect 526 4028 530 4032
rect 534 4028 538 4032
rect 498 4003 502 4007
rect 505 4003 509 4007
rect 486 3988 490 3992
rect 510 3988 514 3992
rect 486 3978 490 3982
rect 462 3928 466 3932
rect 454 3918 458 3922
rect 486 3908 490 3912
rect 518 3938 522 3942
rect 510 3898 514 3902
rect 462 3888 466 3892
rect 350 3858 354 3862
rect 374 3858 378 3862
rect 390 3838 394 3842
rect 510 3838 514 3842
rect 318 3788 322 3792
rect 326 3788 330 3792
rect 174 3758 178 3762
rect 254 3738 258 3742
rect 158 3728 162 3732
rect 134 3678 138 3682
rect 110 3668 114 3672
rect 134 3668 138 3672
rect 94 3658 98 3662
rect 126 3658 130 3662
rect 110 3648 114 3652
rect 126 3558 130 3562
rect 30 3528 34 3532
rect 86 3518 90 3522
rect 30 3468 34 3472
rect 78 3478 82 3482
rect 54 3468 58 3472
rect 46 3458 50 3462
rect 6 3448 10 3452
rect 30 3368 34 3372
rect 30 3358 34 3362
rect 6 3348 10 3352
rect 54 3348 58 3352
rect 30 3338 34 3342
rect 54 3338 58 3342
rect 126 3528 130 3532
rect 142 3478 146 3482
rect 366 3738 370 3742
rect 270 3718 274 3722
rect 262 3678 266 3682
rect 222 3668 226 3672
rect 286 3668 290 3672
rect 326 3658 330 3662
rect 342 3658 346 3662
rect 382 3658 386 3662
rect 190 3648 194 3652
rect 198 3568 202 3572
rect 286 3558 290 3562
rect 318 3558 322 3562
rect 374 3568 378 3572
rect 498 3803 502 3807
rect 505 3803 509 3807
rect 430 3798 434 3802
rect 502 3768 506 3772
rect 422 3738 426 3742
rect 446 3728 450 3732
rect 518 3728 522 3732
rect 638 4148 642 4152
rect 670 4138 674 4142
rect 558 4128 562 4132
rect 638 4128 642 4132
rect 654 4128 658 4132
rect 606 4118 610 4122
rect 598 4108 602 4112
rect 606 4078 610 4082
rect 574 4058 578 4062
rect 598 4058 602 4062
rect 686 4108 690 4112
rect 686 4078 690 4082
rect 630 4048 634 4052
rect 662 4048 666 4052
rect 558 4028 562 4032
rect 566 4018 570 4022
rect 622 3988 626 3992
rect 702 4148 706 4152
rect 718 4158 722 4162
rect 782 4348 786 4352
rect 798 4348 802 4352
rect 918 4348 922 4352
rect 782 4328 786 4332
rect 798 4328 802 4332
rect 734 4318 738 4322
rect 766 4318 770 4322
rect 734 4288 738 4292
rect 838 4318 842 4322
rect 806 4278 810 4282
rect 830 4258 834 4262
rect 806 4248 810 4252
rect 750 4238 754 4242
rect 806 4238 810 4242
rect 790 4228 794 4232
rect 734 4148 738 4152
rect 774 4148 778 4152
rect 726 4138 730 4142
rect 750 4138 754 4142
rect 702 4088 706 4092
rect 726 4118 730 4122
rect 718 4098 722 4102
rect 718 4088 722 4092
rect 758 4098 762 4102
rect 750 4078 754 4082
rect 710 4038 714 4042
rect 702 4008 706 4012
rect 702 3988 706 3992
rect 630 3968 634 3972
rect 550 3948 554 3952
rect 598 3928 602 3932
rect 614 3928 618 3932
rect 806 4168 810 4172
rect 790 4158 794 4162
rect 814 4148 818 4152
rect 806 4138 810 4142
rect 846 4308 850 4312
rect 846 4288 850 4292
rect 862 4328 866 4332
rect 926 4328 930 4332
rect 942 4358 946 4362
rect 1534 4358 1538 4362
rect 974 4348 978 4352
rect 942 4338 946 4342
rect 982 4338 986 4342
rect 958 4318 962 4322
rect 966 4288 970 4292
rect 1002 4303 1006 4307
rect 1009 4303 1013 4307
rect 894 4278 898 4282
rect 918 4278 922 4282
rect 990 4278 994 4282
rect 998 4278 1002 4282
rect 1046 4278 1050 4282
rect 1062 4278 1066 4282
rect 862 4268 866 4272
rect 838 4208 842 4212
rect 822 4128 826 4132
rect 814 4118 818 4122
rect 822 4108 826 4112
rect 766 4088 770 4092
rect 782 4088 786 4092
rect 830 4098 834 4102
rect 830 4088 834 4092
rect 766 4078 770 4082
rect 798 4078 802 4082
rect 822 4078 826 4082
rect 870 4258 874 4262
rect 878 4248 882 4252
rect 854 4228 858 4232
rect 934 4268 938 4272
rect 966 4268 970 4272
rect 902 4258 906 4262
rect 958 4258 962 4262
rect 1038 4268 1042 4272
rect 1030 4258 1034 4262
rect 1046 4258 1050 4262
rect 1054 4248 1058 4252
rect 886 4218 890 4222
rect 910 4218 914 4222
rect 870 4188 874 4192
rect 878 4178 882 4182
rect 926 4158 930 4162
rect 854 4148 858 4152
rect 870 4148 874 4152
rect 894 4138 898 4142
rect 910 4138 914 4142
rect 878 4118 882 4122
rect 846 4078 850 4082
rect 838 4068 842 4072
rect 846 4068 850 4072
rect 782 4058 786 4062
rect 830 4058 834 4062
rect 886 4078 890 4082
rect 894 4078 898 4082
rect 902 4068 906 4072
rect 918 4058 922 4062
rect 942 4238 946 4242
rect 966 4238 970 4242
rect 950 4188 954 4192
rect 1038 4178 1042 4182
rect 1046 4178 1050 4182
rect 958 4168 962 4172
rect 966 4168 970 4172
rect 1014 4148 1018 4152
rect 942 4118 946 4122
rect 1134 4338 1138 4342
rect 1086 4328 1090 4332
rect 1102 4278 1106 4282
rect 1150 4278 1154 4282
rect 1118 4268 1122 4272
rect 1134 4268 1138 4272
rect 1094 4258 1098 4262
rect 1134 4258 1138 4262
rect 1158 4268 1162 4272
rect 1126 4248 1130 4252
rect 1118 4238 1122 4242
rect 1150 4238 1154 4242
rect 1086 4218 1090 4222
rect 1110 4218 1114 4222
rect 1094 4198 1098 4202
rect 1094 4178 1098 4182
rect 1070 4158 1074 4162
rect 1062 4148 1066 4152
rect 1078 4148 1082 4152
rect 1054 4138 1058 4142
rect 1070 4138 1074 4142
rect 1086 4138 1090 4142
rect 1022 4128 1026 4132
rect 1070 4128 1074 4132
rect 974 4118 978 4122
rect 958 4108 962 4112
rect 990 4108 994 4112
rect 966 4098 970 4102
rect 982 4088 986 4092
rect 1002 4103 1006 4107
rect 1009 4103 1013 4107
rect 1030 4118 1034 4122
rect 1038 4118 1042 4122
rect 958 4078 962 4082
rect 998 4078 1002 4082
rect 934 4068 938 4072
rect 974 4068 978 4072
rect 990 4068 994 4072
rect 942 4058 946 4062
rect 950 4058 954 4062
rect 758 4048 762 4052
rect 766 4048 770 4052
rect 782 4048 786 4052
rect 790 4048 794 4052
rect 806 4048 810 4052
rect 862 4048 866 4052
rect 926 4048 930 4052
rect 846 4038 850 4042
rect 886 4038 890 4042
rect 734 4028 738 4032
rect 766 4028 770 4032
rect 726 3928 730 3932
rect 630 3918 634 3922
rect 582 3908 586 3912
rect 558 3898 562 3902
rect 574 3898 578 3902
rect 558 3878 562 3882
rect 542 3868 546 3872
rect 630 3898 634 3902
rect 790 3998 794 4002
rect 854 3988 858 3992
rect 910 4008 914 4012
rect 894 3978 898 3982
rect 894 3958 898 3962
rect 790 3948 794 3952
rect 814 3948 818 3952
rect 830 3948 834 3952
rect 766 3938 770 3942
rect 750 3918 754 3922
rect 774 3898 778 3902
rect 606 3888 610 3892
rect 694 3888 698 3892
rect 710 3888 714 3892
rect 766 3888 770 3892
rect 638 3878 642 3882
rect 686 3878 690 3882
rect 726 3878 730 3882
rect 574 3868 578 3872
rect 718 3868 722 3872
rect 806 3938 810 3942
rect 806 3928 810 3932
rect 806 3878 810 3882
rect 558 3738 562 3742
rect 550 3718 554 3722
rect 502 3678 506 3682
rect 542 3668 546 3672
rect 446 3558 450 3562
rect 414 3548 418 3552
rect 414 3538 418 3542
rect 438 3538 442 3542
rect 630 3858 634 3862
rect 766 3858 770 3862
rect 614 3798 618 3802
rect 662 3848 666 3852
rect 710 3848 714 3852
rect 630 3778 634 3782
rect 678 3778 682 3782
rect 646 3758 650 3762
rect 790 3858 794 3862
rect 854 3918 858 3922
rect 838 3898 842 3902
rect 854 3898 858 3902
rect 1062 4058 1066 4062
rect 1134 4188 1138 4192
rect 1142 4158 1146 4162
rect 1126 4148 1130 4152
rect 1086 4068 1090 4072
rect 1046 4048 1050 4052
rect 1094 4038 1098 4042
rect 1126 4118 1130 4122
rect 1166 4188 1170 4192
rect 1158 4118 1162 4122
rect 1134 4068 1138 4072
rect 1110 4028 1114 4032
rect 1110 4018 1114 4022
rect 1030 3998 1034 4002
rect 1038 3988 1042 3992
rect 950 3958 954 3962
rect 950 3948 954 3952
rect 1054 3948 1058 3952
rect 1038 3938 1042 3942
rect 1002 3903 1006 3907
rect 1009 3903 1013 3907
rect 942 3888 946 3892
rect 926 3878 930 3882
rect 910 3868 914 3872
rect 950 3868 954 3872
rect 982 3868 986 3872
rect 846 3858 850 3862
rect 902 3858 906 3862
rect 814 3848 818 3852
rect 830 3848 834 3852
rect 854 3848 858 3852
rect 926 3848 930 3852
rect 870 3838 874 3842
rect 974 3818 978 3822
rect 750 3758 754 3762
rect 726 3748 730 3752
rect 758 3748 762 3752
rect 614 3738 618 3742
rect 766 3738 770 3742
rect 662 3718 666 3722
rect 590 3688 594 3692
rect 702 3718 706 3722
rect 670 3688 674 3692
rect 734 3718 738 3722
rect 498 3603 502 3607
rect 505 3603 509 3607
rect 494 3578 498 3582
rect 486 3568 490 3572
rect 454 3548 458 3552
rect 558 3568 562 3572
rect 526 3558 530 3562
rect 566 3548 570 3552
rect 574 3538 578 3542
rect 230 3528 234 3532
rect 318 3528 322 3532
rect 190 3518 194 3522
rect 230 3488 234 3492
rect 374 3488 378 3492
rect 310 3478 314 3482
rect 374 3478 378 3482
rect 78 3468 82 3472
rect 94 3468 98 3472
rect 118 3468 122 3472
rect 286 3468 290 3472
rect 126 3458 130 3462
rect 222 3458 226 3462
rect 254 3458 258 3462
rect 286 3458 290 3462
rect 302 3458 306 3462
rect 174 3448 178 3452
rect 366 3458 370 3462
rect 206 3368 210 3372
rect 110 3358 114 3362
rect 142 3348 146 3352
rect 366 3358 370 3362
rect 110 3328 114 3332
rect 70 3298 74 3302
rect 62 3268 66 3272
rect 110 3268 114 3272
rect 86 3258 90 3262
rect 102 3218 106 3222
rect 38 3168 42 3172
rect 86 3168 90 3172
rect 102 3158 106 3162
rect 14 3148 18 3152
rect 30 3148 34 3152
rect 6 3138 10 3142
rect 62 3148 66 3152
rect 78 3148 82 3152
rect 46 3128 50 3132
rect 94 3128 98 3132
rect 6 3078 10 3082
rect 38 3068 42 3072
rect 14 3058 18 3062
rect 30 3058 34 3062
rect 54 3118 58 3122
rect 78 3068 82 3072
rect 38 3038 42 3042
rect 6 2948 10 2952
rect 14 2948 18 2952
rect 126 3248 130 3252
rect 302 3348 306 3352
rect 342 3338 346 3342
rect 366 3338 370 3342
rect 390 3468 394 3472
rect 190 3328 194 3332
rect 270 3328 274 3332
rect 374 3328 378 3332
rect 182 3318 186 3322
rect 230 3318 234 3322
rect 174 3298 178 3302
rect 142 3148 146 3152
rect 126 3138 130 3142
rect 150 3138 154 3142
rect 230 3288 234 3292
rect 238 3278 242 3282
rect 294 3308 298 3312
rect 534 3488 538 3492
rect 422 3478 426 3482
rect 446 3478 450 3482
rect 478 3478 482 3482
rect 438 3468 442 3472
rect 510 3468 514 3472
rect 446 3448 450 3452
rect 470 3448 474 3452
rect 494 3448 498 3452
rect 518 3448 522 3452
rect 454 3438 458 3442
rect 502 3438 506 3442
rect 498 3403 502 3407
rect 505 3403 509 3407
rect 430 3378 434 3382
rect 318 3318 322 3322
rect 358 3318 362 3322
rect 398 3318 402 3322
rect 406 3318 410 3322
rect 262 3288 266 3292
rect 302 3288 306 3292
rect 238 3268 242 3272
rect 310 3268 314 3272
rect 326 3268 330 3272
rect 206 3258 210 3262
rect 270 3258 274 3262
rect 286 3258 290 3262
rect 214 3248 218 3252
rect 230 3248 234 3252
rect 214 3218 218 3222
rect 246 3178 250 3182
rect 238 3168 242 3172
rect 294 3248 298 3252
rect 382 3288 386 3292
rect 398 3278 402 3282
rect 422 3308 426 3312
rect 558 3478 562 3482
rect 558 3378 562 3382
rect 582 3378 586 3382
rect 542 3368 546 3372
rect 566 3358 570 3362
rect 662 3668 666 3672
rect 630 3658 634 3662
rect 726 3658 730 3662
rect 622 3648 626 3652
rect 774 3638 778 3642
rect 614 3628 618 3632
rect 774 3628 778 3632
rect 742 3568 746 3572
rect 766 3568 770 3572
rect 742 3558 746 3562
rect 630 3548 634 3552
rect 646 3548 650 3552
rect 758 3548 762 3552
rect 902 3798 906 3802
rect 1070 3878 1074 3882
rect 1022 3768 1026 3772
rect 790 3758 794 3762
rect 934 3748 938 3752
rect 806 3688 810 3692
rect 782 3548 786 3552
rect 790 3548 794 3552
rect 670 3528 674 3532
rect 606 3488 610 3492
rect 726 3508 730 3512
rect 662 3478 666 3482
rect 750 3488 754 3492
rect 734 3468 738 3472
rect 750 3468 754 3472
rect 662 3458 666 3462
rect 726 3438 730 3442
rect 526 3338 530 3342
rect 590 3338 594 3342
rect 470 3328 474 3332
rect 438 3308 442 3312
rect 454 3278 458 3282
rect 598 3318 602 3322
rect 534 3308 538 3312
rect 606 3298 610 3302
rect 694 3378 698 3382
rect 654 3368 658 3372
rect 638 3348 642 3352
rect 678 3348 682 3352
rect 630 3338 634 3342
rect 622 3288 626 3292
rect 510 3278 514 3282
rect 446 3268 450 3272
rect 470 3268 474 3272
rect 486 3268 490 3272
rect 374 3258 378 3262
rect 542 3258 546 3262
rect 558 3248 562 3252
rect 342 3238 346 3242
rect 382 3238 386 3242
rect 294 3168 298 3172
rect 334 3168 338 3172
rect 350 3168 354 3172
rect 198 3158 202 3162
rect 238 3158 242 3162
rect 254 3158 258 3162
rect 270 3158 274 3162
rect 278 3158 282 3162
rect 342 3158 346 3162
rect 382 3158 386 3162
rect 406 3158 410 3162
rect 190 3148 194 3152
rect 182 3138 186 3142
rect 190 3138 194 3142
rect 150 3088 154 3092
rect 174 3108 178 3112
rect 254 3148 258 3152
rect 246 3128 250 3132
rect 262 3128 266 3132
rect 262 3118 266 3122
rect 182 3088 186 3092
rect 246 3088 250 3092
rect 222 3078 226 3082
rect 246 3078 250 3082
rect 174 3068 178 3072
rect 158 3058 162 3062
rect 110 3048 114 3052
rect 190 3048 194 3052
rect 150 3028 154 3032
rect 118 2988 122 2992
rect 262 3108 266 3112
rect 498 3203 502 3207
rect 505 3203 509 3207
rect 294 3148 298 3152
rect 326 3148 330 3152
rect 342 3148 346 3152
rect 374 3148 378 3152
rect 398 3148 402 3152
rect 446 3148 450 3152
rect 470 3148 474 3152
rect 486 3148 490 3152
rect 278 3138 282 3142
rect 350 3138 354 3142
rect 366 3138 370 3142
rect 382 3138 386 3142
rect 310 3128 314 3132
rect 334 3128 338 3132
rect 318 3108 322 3112
rect 286 3058 290 3062
rect 262 3048 266 3052
rect 270 3048 274 3052
rect 278 3048 282 3052
rect 310 3038 314 3042
rect 270 3028 274 3032
rect 310 2958 314 2962
rect 246 2948 250 2952
rect 30 2878 34 2882
rect 62 2878 66 2882
rect 70 2878 74 2882
rect 86 2868 90 2872
rect 110 2868 114 2872
rect 126 2868 130 2872
rect 150 2938 154 2942
rect 174 2928 178 2932
rect 166 2918 170 2922
rect 326 3088 330 3092
rect 366 3118 370 3122
rect 422 3138 426 3142
rect 454 3138 458 3142
rect 430 3128 434 3132
rect 454 3128 458 3132
rect 406 3118 410 3122
rect 430 3108 434 3112
rect 438 3108 442 3112
rect 566 3158 570 3162
rect 502 3148 506 3152
rect 534 3148 538 3152
rect 622 3248 626 3252
rect 646 3338 650 3342
rect 726 3358 730 3362
rect 678 3328 682 3332
rect 710 3328 714 3332
rect 654 3298 658 3302
rect 526 3138 530 3142
rect 510 3118 514 3122
rect 398 3078 402 3082
rect 334 3068 338 3072
rect 390 3068 394 3072
rect 326 3048 330 3052
rect 318 2928 322 2932
rect 310 2918 314 2922
rect 158 2878 162 2882
rect 62 2858 66 2862
rect 142 2858 146 2862
rect 6 2848 10 2852
rect 110 2848 114 2852
rect 14 2748 18 2752
rect 46 2748 50 2752
rect 142 2748 146 2752
rect 6 2728 10 2732
rect 22 2738 26 2742
rect 70 2738 74 2742
rect 94 2728 98 2732
rect 70 2718 74 2722
rect 78 2708 82 2712
rect 14 2688 18 2692
rect 22 2668 26 2672
rect 46 2668 50 2672
rect 70 2668 74 2672
rect 118 2668 122 2672
rect 190 2848 194 2852
rect 158 2728 162 2732
rect 142 2688 146 2692
rect 190 2708 194 2712
rect 142 2678 146 2682
rect 78 2658 82 2662
rect 102 2658 106 2662
rect 134 2658 138 2662
rect 6 2648 10 2652
rect 6 2558 10 2562
rect 46 2558 50 2562
rect 70 2548 74 2552
rect 22 2538 26 2542
rect 70 2538 74 2542
rect 222 2668 226 2672
rect 182 2658 186 2662
rect 262 2888 266 2892
rect 302 2898 306 2902
rect 270 2858 274 2862
rect 286 2858 290 2862
rect 270 2848 274 2852
rect 342 3048 346 3052
rect 398 3048 402 3052
rect 550 3128 554 3132
rect 582 3128 586 3132
rect 542 3118 546 3122
rect 598 3108 602 3112
rect 726 3318 730 3322
rect 870 3738 874 3742
rect 910 3728 914 3732
rect 870 3678 874 3682
rect 1022 3718 1026 3722
rect 1002 3703 1006 3707
rect 1009 3703 1013 3707
rect 990 3678 994 3682
rect 910 3668 914 3672
rect 926 3668 930 3672
rect 1038 3838 1042 3842
rect 1062 3758 1066 3762
rect 1110 3838 1114 3842
rect 1102 3788 1106 3792
rect 1286 4338 1290 4342
rect 1318 4338 1322 4342
rect 1270 4278 1274 4282
rect 1390 4318 1394 4322
rect 1502 4338 1506 4342
rect 1510 4318 1514 4322
rect 1422 4278 1426 4282
rect 1478 4278 1482 4282
rect 1182 4268 1186 4272
rect 1222 4268 1226 4272
rect 1238 4268 1242 4272
rect 1254 4268 1258 4272
rect 1502 4268 1506 4272
rect 1198 4258 1202 4262
rect 1206 4248 1210 4252
rect 1238 4258 1242 4262
rect 1222 4218 1226 4222
rect 1270 4258 1274 4262
rect 1254 4248 1258 4252
rect 1246 4228 1250 4232
rect 1278 4228 1282 4232
rect 1238 4208 1242 4212
rect 1214 4198 1218 4202
rect 1286 4178 1290 4182
rect 1262 4168 1266 4172
rect 1238 4158 1242 4162
rect 1318 4158 1322 4162
rect 1334 4158 1338 4162
rect 1206 4138 1210 4142
rect 1182 4128 1186 4132
rect 1198 4088 1202 4092
rect 1246 4128 1250 4132
rect 1262 4098 1266 4102
rect 1318 4138 1322 4142
rect 1302 4128 1306 4132
rect 1326 4128 1330 4132
rect 1286 4098 1290 4102
rect 1270 4088 1274 4092
rect 1278 4088 1282 4092
rect 1326 4088 1330 4092
rect 1302 4078 1306 4082
rect 1302 4058 1306 4062
rect 1294 4038 1298 4042
rect 1302 4028 1306 4032
rect 1318 3988 1322 3992
rect 1158 3948 1162 3952
rect 1262 3948 1266 3952
rect 1294 3948 1298 3952
rect 1182 3918 1186 3922
rect 1222 3908 1226 3912
rect 1310 3908 1314 3912
rect 1126 3898 1130 3902
rect 1150 3878 1154 3882
rect 1190 3878 1194 3882
rect 1166 3868 1170 3872
rect 1270 3888 1274 3892
rect 1310 3878 1314 3882
rect 1510 4258 1514 4262
rect 1350 4248 1354 4252
rect 1406 4248 1410 4252
rect 1478 4238 1482 4242
rect 1726 4368 1730 4372
rect 1910 4368 1914 4372
rect 1702 4358 1706 4362
rect 1734 4358 1738 4362
rect 1766 4358 1770 4362
rect 2158 4358 2162 4362
rect 2182 4358 2186 4362
rect 2238 4358 2242 4362
rect 2334 4358 2338 4362
rect 2422 4358 2426 4362
rect 2462 4358 2466 4362
rect 2670 4358 2674 4362
rect 2694 4358 2698 4362
rect 2974 4358 2978 4362
rect 2990 4358 2994 4362
rect 3014 4358 3018 4362
rect 1734 4348 1738 4352
rect 1566 4328 1570 4332
rect 1518 4218 1522 4222
rect 1522 4203 1526 4207
rect 1529 4203 1533 4207
rect 1494 4168 1498 4172
rect 1438 4158 1442 4162
rect 1398 4138 1402 4142
rect 1430 4138 1434 4142
rect 1438 4128 1442 4132
rect 1414 4108 1418 4112
rect 1430 4108 1434 4112
rect 1414 4088 1418 4092
rect 1414 4058 1418 4062
rect 1390 4018 1394 4022
rect 1398 4008 1402 4012
rect 1374 3958 1378 3962
rect 1414 3958 1418 3962
rect 1342 3948 1346 3952
rect 1406 3948 1410 3952
rect 1262 3868 1266 3872
rect 1286 3868 1290 3872
rect 1214 3858 1218 3862
rect 1182 3838 1186 3842
rect 1134 3788 1138 3792
rect 1118 3778 1122 3782
rect 1134 3778 1138 3782
rect 1198 3848 1202 3852
rect 1206 3848 1210 3852
rect 1222 3848 1226 3852
rect 1270 3798 1274 3802
rect 1142 3748 1146 3752
rect 1214 3748 1218 3752
rect 1166 3738 1170 3742
rect 1190 3738 1194 3742
rect 1110 3698 1114 3702
rect 1142 3678 1146 3682
rect 1046 3668 1050 3672
rect 918 3658 922 3662
rect 982 3658 986 3662
rect 1030 3658 1034 3662
rect 838 3648 842 3652
rect 1158 3708 1162 3712
rect 1158 3698 1162 3702
rect 1334 3868 1338 3872
rect 1382 3868 1386 3872
rect 1326 3858 1330 3862
rect 1406 3848 1410 3852
rect 1574 4258 1578 4262
rect 1590 4258 1594 4262
rect 1606 4238 1610 4242
rect 1622 4158 1626 4162
rect 1470 4128 1474 4132
rect 1518 4128 1522 4132
rect 1566 4128 1570 4132
rect 1486 4098 1490 4102
rect 1550 4098 1554 4102
rect 1542 4088 1546 4092
rect 1518 4078 1522 4082
rect 1502 4068 1506 4072
rect 1526 4068 1530 4072
rect 1878 4347 1882 4351
rect 1902 4348 1906 4352
rect 1710 4338 1714 4342
rect 1758 4338 1762 4342
rect 1694 4318 1698 4322
rect 1766 4328 1770 4332
rect 1798 4328 1802 4332
rect 1886 4328 1890 4332
rect 1718 4278 1722 4282
rect 1846 4278 1850 4282
rect 1662 4228 1666 4232
rect 1750 4268 1754 4272
rect 1822 4268 1826 4272
rect 1782 4238 1786 4242
rect 1806 4238 1810 4242
rect 1702 4228 1706 4232
rect 1678 4218 1682 4222
rect 1798 4188 1802 4192
rect 1790 4178 1794 4182
rect 1750 4158 1754 4162
rect 1670 4148 1674 4152
rect 1638 4098 1642 4102
rect 1654 4098 1658 4102
rect 1638 4088 1642 4092
rect 1614 4078 1618 4082
rect 1486 4058 1490 4062
rect 1494 4048 1498 4052
rect 1462 4038 1466 4042
rect 1494 4038 1498 4042
rect 1502 4038 1506 4042
rect 1486 4018 1490 4022
rect 1522 4003 1526 4007
rect 1529 4003 1533 4007
rect 1542 3998 1546 4002
rect 1542 3978 1546 3982
rect 1534 3958 1538 3962
rect 1614 4048 1618 4052
rect 1606 4018 1610 4022
rect 1646 3978 1650 3982
rect 1350 3838 1354 3842
rect 1374 3838 1378 3842
rect 1422 3838 1426 3842
rect 1294 3768 1298 3772
rect 1326 3768 1330 3772
rect 1470 3858 1474 3862
rect 1438 3798 1442 3802
rect 1398 3778 1402 3782
rect 1478 3778 1482 3782
rect 1390 3768 1394 3772
rect 1286 3758 1290 3762
rect 1358 3758 1362 3762
rect 1278 3738 1282 3742
rect 1198 3718 1202 3722
rect 1214 3718 1218 3722
rect 1262 3718 1266 3722
rect 1174 3688 1178 3692
rect 1182 3688 1186 3692
rect 1230 3708 1234 3712
rect 1206 3668 1210 3672
rect 1350 3748 1354 3752
rect 1310 3728 1314 3732
rect 1294 3718 1298 3722
rect 1302 3688 1306 3692
rect 1286 3678 1290 3682
rect 1430 3768 1434 3772
rect 1438 3768 1442 3772
rect 1470 3758 1474 3762
rect 1510 3918 1514 3922
rect 1502 3908 1506 3912
rect 1542 3908 1546 3912
rect 1502 3898 1506 3902
rect 1526 3878 1530 3882
rect 1590 3878 1594 3882
rect 1622 3868 1626 3872
rect 1566 3858 1570 3862
rect 1522 3803 1526 3807
rect 1529 3803 1533 3807
rect 1502 3768 1506 3772
rect 1486 3758 1490 3762
rect 1558 3758 1562 3762
rect 1606 3758 1610 3762
rect 1550 3748 1554 3752
rect 1382 3738 1386 3742
rect 1406 3738 1410 3742
rect 1446 3738 1450 3742
rect 1366 3728 1370 3732
rect 1350 3668 1354 3672
rect 1246 3658 1250 3662
rect 1054 3648 1058 3652
rect 1126 3648 1130 3652
rect 1150 3648 1154 3652
rect 862 3628 866 3632
rect 886 3548 890 3552
rect 1246 3588 1250 3592
rect 1142 3558 1146 3562
rect 1174 3558 1178 3562
rect 1374 3638 1378 3642
rect 1422 3728 1426 3732
rect 1454 3698 1458 3702
rect 1446 3678 1450 3682
rect 1502 3728 1506 3732
rect 1478 3718 1482 3722
rect 1518 3698 1522 3702
rect 1438 3668 1442 3672
rect 1470 3668 1474 3672
rect 1438 3618 1442 3622
rect 1414 3588 1418 3592
rect 1390 3558 1394 3562
rect 1522 3603 1526 3607
rect 1529 3603 1533 3607
rect 1086 3547 1090 3551
rect 1254 3548 1258 3552
rect 1390 3548 1394 3552
rect 1510 3547 1514 3551
rect 1534 3548 1538 3552
rect 1574 3738 1578 3742
rect 1694 4118 1698 4122
rect 1686 4108 1690 4112
rect 1718 4148 1722 4152
rect 1710 4138 1714 4142
rect 1774 4138 1778 4142
rect 1742 4128 1746 4132
rect 1758 4128 1762 4132
rect 1718 4108 1722 4112
rect 1702 4098 1706 4102
rect 1742 4098 1746 4102
rect 1678 4078 1682 4082
rect 1662 4068 1666 4072
rect 1710 4068 1714 4072
rect 1886 4258 1890 4262
rect 1814 4218 1818 4222
rect 1822 4208 1826 4212
rect 1894 4228 1898 4232
rect 1838 4198 1842 4202
rect 1814 4178 1818 4182
rect 1806 4158 1810 4162
rect 2014 4348 2018 4352
rect 1966 4328 1970 4332
rect 1910 4288 1914 4292
rect 1950 4278 1954 4282
rect 1966 4268 1970 4272
rect 1998 4258 2002 4262
rect 1974 4248 1978 4252
rect 1966 4218 1970 4222
rect 1990 4238 1994 4242
rect 2078 4328 2082 4332
rect 2026 4303 2030 4307
rect 2033 4303 2037 4307
rect 2134 4338 2138 4342
rect 2078 4298 2082 4302
rect 2134 4298 2138 4302
rect 2022 4288 2026 4292
rect 2086 4288 2090 4292
rect 2094 4288 2098 4292
rect 2118 4288 2122 4292
rect 2030 4268 2034 4272
rect 2014 4218 2018 4222
rect 1998 4208 2002 4212
rect 1942 4188 1946 4192
rect 1926 4178 1930 4182
rect 1854 4148 1858 4152
rect 1862 4148 1866 4152
rect 1822 4138 1826 4142
rect 1838 4138 1842 4142
rect 1886 4138 1890 4142
rect 1790 4108 1794 4112
rect 1766 4078 1770 4082
rect 1782 4078 1786 4082
rect 1814 4078 1818 4082
rect 1774 4068 1778 4072
rect 1806 4068 1810 4072
rect 1846 4078 1850 4082
rect 1870 4068 1874 4072
rect 1742 4058 1746 4062
rect 1790 4058 1794 4062
rect 1854 4058 1858 4062
rect 1862 4058 1866 4062
rect 1662 3968 1666 3972
rect 1822 4038 1826 4042
rect 1822 4018 1826 4022
rect 1782 4008 1786 4012
rect 1766 3988 1770 3992
rect 1822 3988 1826 3992
rect 1782 3958 1786 3962
rect 1814 3958 1818 3962
rect 1694 3928 1698 3932
rect 1782 3938 1786 3942
rect 1878 4048 1882 4052
rect 1926 4148 1930 4152
rect 1942 4148 1946 4152
rect 1910 4138 1914 4142
rect 1966 4138 1970 4142
rect 1974 4128 1978 4132
rect 1982 4118 1986 4122
rect 1958 4058 1962 4062
rect 1934 4048 1938 4052
rect 1950 4048 1954 4052
rect 1974 4048 1978 4052
rect 1950 4038 1954 4042
rect 1926 4018 1930 4022
rect 1918 3998 1922 4002
rect 1902 3958 1906 3962
rect 2006 4168 2010 4172
rect 2078 4228 2082 4232
rect 2038 4218 2042 4222
rect 2118 4218 2122 4222
rect 2030 4208 2034 4212
rect 2046 4168 2050 4172
rect 2014 4148 2018 4152
rect 2022 4148 2026 4152
rect 2026 4103 2030 4107
rect 2033 4103 2037 4107
rect 1998 4078 2002 4082
rect 1982 4008 1986 4012
rect 2006 4058 2010 4062
rect 1998 4038 2002 4042
rect 1990 3988 1994 3992
rect 1966 3958 1970 3962
rect 1982 3958 1986 3962
rect 2014 3958 2018 3962
rect 1806 3938 1810 3942
rect 1814 3938 1818 3942
rect 1846 3938 1850 3942
rect 1854 3938 1858 3942
rect 1734 3908 1738 3912
rect 1766 3908 1770 3912
rect 1718 3878 1722 3882
rect 1726 3878 1730 3882
rect 1686 3848 1690 3852
rect 1750 3838 1754 3842
rect 1694 3788 1698 3792
rect 1686 3758 1690 3762
rect 1670 3748 1674 3752
rect 1678 3738 1682 3742
rect 1750 3748 1754 3752
rect 1726 3698 1730 3702
rect 1790 3858 1794 3862
rect 1774 3848 1778 3852
rect 1838 3928 1842 3932
rect 1894 3938 1898 3942
rect 1902 3938 1906 3942
rect 1878 3928 1882 3932
rect 1886 3928 1890 3932
rect 1878 3918 1882 3922
rect 1862 3878 1866 3882
rect 1854 3848 1858 3852
rect 1862 3848 1866 3852
rect 1830 3838 1834 3842
rect 1806 3788 1810 3792
rect 1766 3747 1770 3751
rect 1910 3868 1914 3872
rect 1870 3788 1874 3792
rect 1854 3768 1858 3772
rect 1758 3738 1762 3742
rect 1814 3728 1818 3732
rect 1830 3728 1834 3732
rect 1878 3758 1882 3762
rect 1854 3738 1858 3742
rect 1878 3738 1882 3742
rect 1854 3728 1858 3732
rect 1838 3708 1842 3712
rect 1806 3698 1810 3702
rect 1750 3688 1754 3692
rect 1838 3688 1842 3692
rect 1950 3928 1954 3932
rect 1974 3928 1978 3932
rect 1918 3808 1922 3812
rect 1934 3858 1938 3862
rect 1950 3838 1954 3842
rect 2070 4148 2074 4152
rect 2102 4198 2106 4202
rect 2094 4178 2098 4182
rect 2110 4148 2114 4152
rect 2086 4138 2090 4142
rect 2078 4128 2082 4132
rect 2054 4068 2058 4072
rect 2062 4068 2066 4072
rect 2070 4058 2074 4062
rect 2086 4048 2090 4052
rect 2142 4188 2146 4192
rect 2118 4128 2122 4132
rect 2142 4128 2146 4132
rect 2142 4118 2146 4122
rect 2118 4078 2122 4082
rect 2158 4348 2162 4352
rect 2286 4348 2290 4352
rect 2166 4338 2170 4342
rect 2174 4328 2178 4332
rect 2206 4328 2210 4332
rect 2214 4328 2218 4332
rect 2238 4328 2242 4332
rect 2166 4248 2170 4252
rect 2230 4268 2234 4272
rect 2182 4238 2186 4242
rect 2166 4228 2170 4232
rect 2182 4198 2186 4202
rect 2182 4168 2186 4172
rect 2158 4148 2162 4152
rect 2206 4248 2210 4252
rect 2206 4208 2210 4212
rect 2214 4208 2218 4212
rect 2206 4168 2210 4172
rect 2214 4158 2218 4162
rect 2222 4138 2226 4142
rect 2182 4128 2186 4132
rect 2174 4118 2178 4122
rect 2222 4108 2226 4112
rect 2302 4338 2306 4342
rect 2310 4328 2314 4332
rect 2406 4328 2410 4332
rect 2294 4268 2298 4272
rect 2326 4268 2330 4272
rect 3478 4368 3482 4372
rect 3502 4368 3506 4372
rect 3570 4403 3574 4407
rect 3577 4403 3581 4407
rect 3630 4398 3634 4402
rect 3686 4398 3690 4402
rect 3702 4398 3706 4402
rect 3750 4398 3754 4402
rect 3254 4358 3258 4362
rect 3310 4358 3314 4362
rect 3334 4358 3338 4362
rect 3414 4358 3418 4362
rect 3438 4358 3442 4362
rect 3486 4358 3490 4362
rect 3598 4358 3602 4362
rect 3622 4358 3626 4362
rect 2526 4348 2530 4352
rect 2606 4348 2610 4352
rect 2830 4348 2834 4352
rect 2422 4338 2426 4342
rect 2598 4338 2602 4342
rect 2654 4338 2658 4342
rect 2678 4338 2682 4342
rect 2726 4338 2730 4342
rect 2318 4258 2322 4262
rect 2246 4238 2250 4242
rect 2270 4248 2274 4252
rect 2254 4228 2258 4232
rect 2246 4218 2250 4222
rect 2302 4248 2306 4252
rect 2350 4248 2354 4252
rect 2310 4238 2314 4242
rect 2286 4228 2290 4232
rect 2334 4208 2338 4212
rect 2262 4198 2266 4202
rect 2294 4198 2298 4202
rect 2326 4198 2330 4202
rect 2246 4188 2250 4192
rect 2278 4188 2282 4192
rect 2238 4178 2242 4182
rect 2326 4178 2330 4182
rect 2310 4138 2314 4142
rect 2246 4128 2250 4132
rect 2254 4128 2258 4132
rect 2262 4118 2266 4122
rect 2182 4078 2186 4082
rect 2230 4078 2234 4082
rect 2254 4078 2258 4082
rect 2190 4068 2194 4072
rect 2270 4108 2274 4112
rect 2110 4048 2114 4052
rect 2134 4048 2138 4052
rect 2150 4048 2154 4052
rect 2206 4048 2210 4052
rect 2110 4038 2114 4042
rect 2134 4038 2138 4042
rect 2126 4018 2130 4022
rect 2110 4008 2114 4012
rect 2094 3968 2098 3972
rect 2206 4038 2210 4042
rect 2222 4038 2226 4042
rect 2302 4098 2306 4102
rect 2286 4058 2290 4062
rect 2206 4018 2210 4022
rect 2150 3968 2154 3972
rect 2006 3948 2010 3952
rect 2094 3948 2098 3952
rect 2134 3948 2138 3952
rect 1998 3908 2002 3912
rect 2026 3903 2030 3907
rect 2033 3903 2037 3907
rect 2014 3888 2018 3892
rect 1998 3878 2002 3882
rect 2014 3868 2018 3872
rect 2030 3868 2034 3872
rect 1990 3848 1994 3852
rect 1998 3838 2002 3842
rect 1958 3828 1962 3832
rect 1974 3828 1978 3832
rect 1982 3828 1986 3832
rect 1926 3788 1930 3792
rect 1918 3768 1922 3772
rect 1902 3748 1906 3752
rect 1926 3748 1930 3752
rect 1894 3728 1898 3732
rect 1886 3678 1890 3682
rect 1726 3668 1730 3672
rect 1742 3668 1746 3672
rect 1798 3668 1802 3672
rect 1966 3768 1970 3772
rect 1982 3758 1986 3762
rect 2006 3758 2010 3762
rect 1950 3748 1954 3752
rect 1990 3748 1994 3752
rect 1934 3738 1938 3742
rect 1982 3738 1986 3742
rect 1934 3708 1938 3712
rect 1934 3698 1938 3702
rect 1934 3678 1938 3682
rect 1990 3698 1994 3702
rect 1590 3648 1594 3652
rect 1886 3658 1890 3662
rect 1918 3658 1922 3662
rect 2046 3858 2050 3862
rect 2054 3848 2058 3852
rect 2054 3798 2058 3802
rect 2078 3928 2082 3932
rect 2086 3928 2090 3932
rect 2086 3878 2090 3882
rect 2118 3878 2122 3882
rect 2102 3868 2106 3872
rect 2150 3898 2154 3902
rect 2150 3868 2154 3872
rect 2126 3858 2130 3862
rect 2142 3858 2146 3862
rect 2086 3838 2090 3842
rect 2118 3838 2122 3842
rect 2214 3978 2218 3982
rect 2190 3958 2194 3962
rect 2206 3958 2210 3962
rect 2238 3958 2242 3962
rect 2278 3958 2282 3962
rect 2190 3948 2194 3952
rect 2174 3928 2178 3932
rect 2190 3928 2194 3932
rect 2182 3878 2186 3882
rect 2174 3858 2178 3862
rect 2158 3848 2162 3852
rect 2166 3838 2170 3842
rect 2126 3808 2130 3812
rect 2150 3808 2154 3812
rect 2230 3908 2234 3912
rect 2214 3868 2218 3872
rect 2246 3868 2250 3872
rect 2278 3858 2282 3862
rect 2214 3848 2218 3852
rect 2246 3848 2250 3852
rect 2230 3838 2234 3842
rect 2334 4158 2338 4162
rect 2414 4258 2418 4262
rect 2374 4248 2378 4252
rect 2390 4228 2394 4232
rect 2414 4228 2418 4232
rect 2382 4188 2386 4192
rect 2398 4178 2402 4182
rect 2406 4158 2410 4162
rect 2350 4148 2354 4152
rect 2366 4138 2370 4142
rect 2350 4128 2354 4132
rect 2358 4118 2362 4122
rect 2398 4108 2402 4112
rect 2350 4098 2354 4102
rect 2382 4098 2386 4102
rect 2342 4078 2346 4082
rect 2334 4068 2338 4072
rect 2342 4058 2346 4062
rect 2358 4068 2362 4072
rect 2398 4058 2402 4062
rect 2438 4288 2442 4292
rect 2662 4328 2666 4332
rect 2886 4338 2890 4342
rect 2942 4338 2946 4342
rect 2974 4338 2978 4342
rect 2670 4318 2674 4322
rect 2462 4298 2466 4302
rect 2454 4288 2458 4292
rect 2494 4278 2498 4282
rect 2478 4268 2482 4272
rect 2446 4258 2450 4262
rect 2438 4248 2442 4252
rect 2526 4268 2530 4272
rect 2518 4248 2522 4252
rect 2966 4328 2970 4332
rect 2814 4318 2818 4322
rect 2710 4308 2714 4312
rect 2774 4298 2778 4302
rect 2702 4288 2706 4292
rect 2718 4278 2722 4282
rect 2574 4248 2578 4252
rect 2598 4248 2602 4252
rect 2454 4238 2458 4242
rect 2486 4238 2490 4242
rect 2526 4238 2530 4242
rect 2542 4238 2546 4242
rect 2598 4238 2602 4242
rect 2638 4268 2642 4272
rect 2686 4268 2690 4272
rect 2766 4268 2770 4272
rect 2662 4258 2666 4262
rect 2702 4258 2706 4262
rect 2630 4248 2634 4252
rect 2654 4248 2658 4252
rect 2670 4248 2674 4252
rect 2750 4248 2754 4252
rect 2486 4228 2490 4232
rect 2614 4228 2618 4232
rect 2494 4218 2498 4222
rect 2590 4218 2594 4222
rect 2546 4203 2550 4207
rect 2553 4203 2557 4207
rect 2462 4188 2466 4192
rect 2430 4168 2434 4172
rect 2422 4158 2426 4162
rect 2454 4168 2458 4172
rect 2502 4178 2506 4182
rect 2486 4168 2490 4172
rect 2486 4158 2490 4162
rect 2534 4158 2538 4162
rect 2438 4148 2442 4152
rect 2462 4148 2466 4152
rect 2502 4148 2506 4152
rect 2422 4108 2426 4112
rect 2446 4068 2450 4072
rect 2478 4108 2482 4112
rect 2502 4108 2506 4112
rect 2462 4078 2466 4082
rect 2438 4058 2442 4062
rect 2454 4058 2458 4062
rect 2326 4048 2330 4052
rect 2414 4048 2418 4052
rect 2430 4048 2434 4052
rect 2294 4028 2298 4032
rect 2358 4038 2362 4042
rect 2374 4038 2378 4042
rect 2414 4038 2418 4042
rect 2430 4038 2434 4042
rect 2486 4058 2490 4062
rect 2318 3968 2322 3972
rect 2350 3968 2354 3972
rect 2470 4018 2474 4022
rect 2358 3948 2362 3952
rect 2326 3938 2330 3942
rect 2342 3938 2346 3942
rect 2422 3978 2426 3982
rect 2454 3978 2458 3982
rect 2382 3948 2386 3952
rect 2374 3928 2378 3932
rect 2494 3928 2498 3932
rect 2382 3918 2386 3922
rect 2302 3898 2306 3902
rect 2286 3828 2290 3832
rect 2230 3818 2234 3822
rect 2126 3788 2130 3792
rect 2158 3788 2162 3792
rect 2102 3778 2106 3782
rect 2134 3778 2138 3782
rect 2158 3768 2162 3772
rect 2070 3758 2074 3762
rect 2126 3758 2130 3762
rect 1822 3648 1826 3652
rect 1942 3648 1946 3652
rect 1862 3638 1866 3642
rect 1886 3628 1890 3632
rect 1654 3618 1658 3622
rect 1918 3588 1922 3592
rect 1966 3658 1970 3662
rect 1982 3658 1986 3662
rect 1950 3638 1954 3642
rect 1646 3568 1650 3572
rect 1742 3568 1746 3572
rect 1574 3548 1578 3552
rect 1622 3548 1626 3552
rect 974 3538 978 3542
rect 990 3538 994 3542
rect 1030 3538 1034 3542
rect 1350 3538 1354 3542
rect 1382 3538 1386 3542
rect 1446 3538 1450 3542
rect 806 3488 810 3492
rect 830 3488 834 3492
rect 1062 3528 1066 3532
rect 1158 3528 1162 3532
rect 1002 3503 1006 3507
rect 1009 3503 1013 3507
rect 1030 3488 1034 3492
rect 942 3478 946 3482
rect 1142 3488 1146 3492
rect 1206 3518 1210 3522
rect 894 3468 898 3472
rect 822 3428 826 3432
rect 782 3418 786 3422
rect 822 3418 826 3422
rect 790 3348 794 3352
rect 694 3298 698 3302
rect 774 3308 778 3312
rect 750 3288 754 3292
rect 662 3218 666 3222
rect 710 3238 714 3242
rect 758 3228 762 3232
rect 726 3208 730 3212
rect 694 3178 698 3182
rect 766 3168 770 3172
rect 678 3128 682 3132
rect 670 3118 674 3122
rect 766 3118 770 3122
rect 702 3098 706 3102
rect 694 3078 698 3082
rect 574 3068 578 3072
rect 590 3058 594 3062
rect 486 3048 490 3052
rect 518 3048 522 3052
rect 598 3048 602 3052
rect 630 3048 634 3052
rect 622 3038 626 3042
rect 430 3028 434 3032
rect 498 3003 502 3007
rect 505 3003 509 3007
rect 374 2998 378 3002
rect 518 2998 522 3002
rect 494 2978 498 2982
rect 342 2968 346 2972
rect 438 2968 442 2972
rect 406 2958 410 2962
rect 462 2908 466 2912
rect 334 2888 338 2892
rect 438 2888 442 2892
rect 366 2848 370 2852
rect 350 2768 354 2772
rect 254 2748 258 2752
rect 430 2848 434 2852
rect 398 2838 402 2842
rect 438 2838 442 2842
rect 446 2828 450 2832
rect 478 2898 482 2902
rect 526 2968 530 2972
rect 534 2968 538 2972
rect 606 2968 610 2972
rect 542 2958 546 2962
rect 534 2898 538 2902
rect 566 2928 570 2932
rect 566 2908 570 2912
rect 550 2898 554 2902
rect 534 2878 538 2882
rect 646 2998 650 3002
rect 798 3308 802 3312
rect 782 3258 786 3262
rect 926 3448 930 3452
rect 870 3428 874 3432
rect 1270 3528 1274 3532
rect 1246 3488 1250 3492
rect 1342 3478 1346 3482
rect 1310 3468 1314 3472
rect 958 3448 962 3452
rect 1198 3458 1202 3462
rect 1150 3418 1154 3422
rect 1198 3418 1202 3422
rect 1038 3388 1042 3392
rect 1070 3388 1074 3392
rect 1102 3388 1106 3392
rect 886 3338 890 3342
rect 926 3338 930 3342
rect 942 3338 946 3342
rect 1014 3328 1018 3332
rect 990 3318 994 3322
rect 1030 3318 1034 3322
rect 1002 3303 1006 3307
rect 1009 3303 1013 3307
rect 1206 3378 1210 3382
rect 1142 3348 1146 3352
rect 1190 3348 1194 3352
rect 1222 3368 1226 3372
rect 1254 3448 1258 3452
rect 1246 3388 1250 3392
rect 1358 3458 1362 3462
rect 1398 3458 1402 3462
rect 1270 3378 1274 3382
rect 1326 3358 1330 3362
rect 1062 3338 1066 3342
rect 1110 3328 1114 3332
rect 1270 3348 1274 3352
rect 1294 3348 1298 3352
rect 1382 3448 1386 3452
rect 1422 3528 1426 3532
rect 1446 3528 1450 3532
rect 1414 3488 1418 3492
rect 1438 3478 1442 3482
rect 1230 3328 1234 3332
rect 1358 3328 1362 3332
rect 1206 3318 1210 3322
rect 1222 3318 1226 3322
rect 1318 3318 1322 3322
rect 1126 3308 1130 3312
rect 814 3268 818 3272
rect 854 3268 858 3272
rect 1190 3268 1194 3272
rect 814 3258 818 3262
rect 790 3248 794 3252
rect 790 3228 794 3232
rect 790 3218 794 3222
rect 798 3148 802 3152
rect 782 3108 786 3112
rect 774 3088 778 3092
rect 766 3078 770 3082
rect 662 3048 666 3052
rect 702 3048 706 3052
rect 710 3048 714 3052
rect 678 3038 682 3042
rect 702 2988 706 2992
rect 638 2978 642 2982
rect 654 2978 658 2982
rect 678 2978 682 2982
rect 670 2958 674 2962
rect 662 2948 666 2952
rect 598 2928 602 2932
rect 614 2928 618 2932
rect 582 2908 586 2912
rect 614 2898 618 2902
rect 630 2898 634 2902
rect 582 2888 586 2892
rect 590 2888 594 2892
rect 758 3058 762 3062
rect 774 3058 778 3062
rect 838 3248 842 3252
rect 814 3108 818 3112
rect 830 3098 834 3102
rect 830 3068 834 3072
rect 790 3058 794 3062
rect 750 3048 754 3052
rect 766 3048 770 3052
rect 750 3018 754 3022
rect 758 3018 762 3022
rect 742 2988 746 2992
rect 726 2978 730 2982
rect 710 2958 714 2962
rect 734 2948 738 2952
rect 646 2938 650 2942
rect 678 2938 682 2942
rect 638 2888 642 2892
rect 662 2928 666 2932
rect 718 2928 722 2932
rect 702 2918 706 2922
rect 670 2908 674 2912
rect 686 2908 690 2912
rect 654 2888 658 2892
rect 694 2898 698 2902
rect 686 2888 690 2892
rect 590 2878 594 2882
rect 598 2878 602 2882
rect 646 2878 650 2882
rect 542 2868 546 2872
rect 478 2858 482 2862
rect 526 2858 530 2862
rect 550 2858 554 2862
rect 590 2858 594 2862
rect 494 2838 498 2842
rect 542 2818 546 2822
rect 498 2803 502 2807
rect 505 2803 509 2807
rect 470 2788 474 2792
rect 462 2758 466 2762
rect 558 2838 562 2842
rect 662 2858 666 2862
rect 750 2958 754 2962
rect 710 2868 714 2872
rect 702 2858 706 2862
rect 694 2838 698 2842
rect 574 2828 578 2832
rect 598 2828 602 2832
rect 414 2688 418 2692
rect 254 2668 258 2672
rect 350 2668 354 2672
rect 246 2658 250 2662
rect 302 2658 306 2662
rect 190 2558 194 2562
rect 30 2528 34 2532
rect 46 2528 50 2532
rect 142 2528 146 2532
rect 70 2478 74 2482
rect 30 2468 34 2472
rect 54 2468 58 2472
rect 62 2458 66 2462
rect 6 2448 10 2452
rect 30 2448 34 2452
rect 46 2388 50 2392
rect 158 2478 162 2482
rect 398 2658 402 2662
rect 582 2688 586 2692
rect 558 2668 562 2672
rect 318 2648 322 2652
rect 366 2648 370 2652
rect 294 2618 298 2622
rect 366 2618 370 2622
rect 286 2538 290 2542
rect 262 2518 266 2522
rect 294 2518 298 2522
rect 246 2498 250 2502
rect 270 2478 274 2482
rect 206 2468 210 2472
rect 142 2458 146 2462
rect 118 2448 122 2452
rect 94 2378 98 2382
rect 110 2378 114 2382
rect 22 2358 26 2362
rect 6 2338 10 2342
rect 14 2338 18 2342
rect 30 2348 34 2352
rect 278 2428 282 2432
rect 190 2378 194 2382
rect 262 2378 266 2382
rect 174 2368 178 2372
rect 142 2358 146 2362
rect 190 2358 194 2362
rect 206 2358 210 2362
rect 158 2348 162 2352
rect 150 2328 154 2332
rect 174 2328 178 2332
rect 118 2308 122 2312
rect 126 2268 130 2272
rect 150 2268 154 2272
rect 174 2268 178 2272
rect 206 2338 210 2342
rect 270 2338 274 2342
rect 206 2328 210 2332
rect 222 2318 226 2322
rect 382 2568 386 2572
rect 542 2648 546 2652
rect 486 2638 490 2642
rect 486 2618 490 2622
rect 542 2608 546 2612
rect 498 2603 502 2607
rect 505 2603 509 2607
rect 638 2818 642 2822
rect 686 2818 690 2822
rect 614 2768 618 2772
rect 622 2758 626 2762
rect 694 2768 698 2772
rect 614 2748 618 2752
rect 630 2748 634 2752
rect 654 2748 658 2752
rect 622 2738 626 2742
rect 670 2738 674 2742
rect 654 2728 658 2732
rect 598 2688 602 2692
rect 654 2688 658 2692
rect 622 2678 626 2682
rect 638 2678 642 2682
rect 590 2658 594 2662
rect 598 2648 602 2652
rect 622 2648 626 2652
rect 646 2648 650 2652
rect 566 2638 570 2642
rect 614 2638 618 2642
rect 462 2548 466 2552
rect 510 2548 514 2552
rect 374 2538 378 2542
rect 422 2538 426 2542
rect 398 2528 402 2532
rect 358 2498 362 2502
rect 334 2478 338 2482
rect 326 2458 330 2462
rect 342 2438 346 2442
rect 342 2358 346 2362
rect 414 2448 418 2452
rect 390 2378 394 2382
rect 406 2378 410 2382
rect 326 2348 330 2352
rect 318 2308 322 2312
rect 526 2538 530 2542
rect 470 2528 474 2532
rect 494 2528 498 2532
rect 470 2518 474 2522
rect 486 2518 490 2522
rect 486 2508 490 2512
rect 478 2468 482 2472
rect 478 2448 482 2452
rect 454 2328 458 2332
rect 398 2318 402 2322
rect 454 2308 458 2312
rect 310 2288 314 2292
rect 334 2288 338 2292
rect 358 2288 362 2292
rect 238 2278 242 2282
rect 302 2278 306 2282
rect 350 2278 354 2282
rect 6 2248 10 2252
rect 78 2228 82 2232
rect 54 2208 58 2212
rect 166 2258 170 2262
rect 38 2188 42 2192
rect 94 2188 98 2192
rect 6 2178 10 2182
rect 22 2178 26 2182
rect 326 2268 330 2272
rect 342 2268 346 2272
rect 382 2258 386 2262
rect 230 2248 234 2252
rect 302 2228 306 2232
rect 318 2178 322 2182
rect 70 2168 74 2172
rect 110 2168 114 2172
rect 198 2168 202 2172
rect 118 2158 122 2162
rect 238 2158 242 2162
rect 310 2158 314 2162
rect 110 2148 114 2152
rect 30 2078 34 2082
rect 6 2048 10 2052
rect 22 2038 26 2042
rect 46 1998 50 2002
rect 102 2138 106 2142
rect 294 2148 298 2152
rect 182 2138 186 2142
rect 318 2148 322 2152
rect 310 2118 314 2122
rect 326 2118 330 2122
rect 262 2078 266 2082
rect 286 2078 290 2082
rect 310 2078 314 2082
rect 214 2068 218 2072
rect 118 2008 122 2012
rect 94 1988 98 1992
rect 30 1978 34 1982
rect 22 1958 26 1962
rect 54 1958 58 1962
rect 118 1958 122 1962
rect 6 1948 10 1952
rect 142 2038 146 2042
rect 166 2028 170 2032
rect 150 1998 154 2002
rect 46 1918 50 1922
rect 22 1888 26 1892
rect 6 1878 10 1882
rect 30 1848 34 1852
rect 38 1788 42 1792
rect 6 1778 10 1782
rect 54 1758 58 1762
rect 54 1748 58 1752
rect 110 1747 114 1751
rect 70 1738 74 1742
rect 22 1688 26 1692
rect 30 1678 34 1682
rect 46 1668 50 1672
rect 134 1858 138 1862
rect 150 1858 154 1862
rect 214 1968 218 1972
rect 246 2038 250 2042
rect 254 2038 258 2042
rect 254 1978 258 1982
rect 206 1938 210 1942
rect 214 1878 218 1882
rect 246 1928 250 1932
rect 270 2068 274 2072
rect 286 2068 290 2072
rect 318 2068 322 2072
rect 366 2168 370 2172
rect 334 2088 338 2092
rect 342 2088 346 2092
rect 294 2058 298 2062
rect 310 2058 314 2062
rect 342 2058 346 2062
rect 382 2158 386 2162
rect 430 2168 434 2172
rect 470 2278 474 2282
rect 470 2228 474 2232
rect 558 2518 562 2522
rect 550 2478 554 2482
rect 518 2448 522 2452
rect 510 2438 514 2442
rect 498 2403 502 2407
rect 505 2403 509 2407
rect 742 2838 746 2842
rect 710 2758 714 2762
rect 782 2998 786 3002
rect 790 2988 794 2992
rect 782 2978 786 2982
rect 798 2978 802 2982
rect 822 2978 826 2982
rect 798 2948 802 2952
rect 958 3238 962 3242
rect 958 3228 962 3232
rect 918 3198 922 3202
rect 1038 3208 1042 3212
rect 982 3188 986 3192
rect 1014 3178 1018 3182
rect 1014 3148 1018 3152
rect 886 3118 890 3122
rect 854 3108 858 3112
rect 862 3068 866 3072
rect 838 3028 842 3032
rect 790 2938 794 2942
rect 774 2908 778 2912
rect 814 2908 818 2912
rect 806 2868 810 2872
rect 806 2858 810 2862
rect 838 2858 842 2862
rect 958 3138 962 3142
rect 1022 3138 1026 3142
rect 950 3128 954 3132
rect 934 3108 938 3112
rect 1002 3103 1006 3107
rect 1009 3103 1013 3107
rect 958 3098 962 3102
rect 998 3088 1002 3092
rect 910 3058 914 3062
rect 926 2968 930 2972
rect 894 2948 898 2952
rect 910 2948 914 2952
rect 990 3048 994 3052
rect 982 2958 986 2962
rect 934 2918 938 2922
rect 990 2948 994 2952
rect 1022 3058 1026 3062
rect 1014 3028 1018 3032
rect 990 2938 994 2942
rect 886 2888 890 2892
rect 870 2878 874 2882
rect 918 2878 922 2882
rect 958 2878 962 2882
rect 854 2868 858 2872
rect 910 2868 914 2872
rect 814 2828 818 2832
rect 846 2828 850 2832
rect 814 2808 818 2812
rect 886 2858 890 2862
rect 950 2858 954 2862
rect 878 2848 882 2852
rect 942 2838 946 2842
rect 966 2848 970 2852
rect 950 2798 954 2802
rect 1002 2903 1006 2907
rect 1009 2903 1013 2907
rect 1046 3038 1050 3042
rect 1118 3208 1122 3212
rect 1158 3208 1162 3212
rect 1102 3178 1106 3182
rect 1230 3288 1234 3292
rect 1286 3278 1290 3282
rect 1262 3268 1266 3272
rect 1238 3258 1242 3262
rect 1150 3158 1154 3162
rect 1102 3078 1106 3082
rect 1070 2958 1074 2962
rect 1086 2958 1090 2962
rect 1070 2928 1074 2932
rect 1078 2928 1082 2932
rect 1078 2908 1082 2912
rect 1062 2898 1066 2902
rect 1038 2858 1042 2862
rect 894 2788 898 2792
rect 766 2758 770 2762
rect 814 2758 818 2762
rect 830 2758 834 2762
rect 1022 2758 1026 2762
rect 846 2748 850 2752
rect 862 2748 866 2752
rect 870 2738 874 2742
rect 910 2738 914 2742
rect 934 2738 938 2742
rect 1030 2738 1034 2742
rect 702 2728 706 2732
rect 718 2728 722 2732
rect 694 2708 698 2712
rect 718 2708 722 2712
rect 702 2698 706 2702
rect 686 2678 690 2682
rect 726 2678 730 2682
rect 822 2718 826 2722
rect 742 2708 746 2712
rect 846 2708 850 2712
rect 854 2708 858 2712
rect 878 2708 882 2712
rect 814 2678 818 2682
rect 838 2678 842 2682
rect 734 2668 738 2672
rect 742 2668 746 2672
rect 766 2668 770 2672
rect 670 2648 674 2652
rect 654 2598 658 2602
rect 702 2658 706 2662
rect 726 2658 730 2662
rect 694 2638 698 2642
rect 710 2648 714 2652
rect 702 2578 706 2582
rect 686 2568 690 2572
rect 710 2568 714 2572
rect 638 2558 642 2562
rect 630 2548 634 2552
rect 654 2548 658 2552
rect 598 2528 602 2532
rect 582 2498 586 2502
rect 566 2478 570 2482
rect 574 2468 578 2472
rect 694 2538 698 2542
rect 646 2528 650 2532
rect 686 2528 690 2532
rect 638 2508 642 2512
rect 638 2498 642 2502
rect 702 2458 706 2462
rect 606 2448 610 2452
rect 614 2448 618 2452
rect 582 2368 586 2372
rect 574 2348 578 2352
rect 510 2318 514 2322
rect 510 2298 514 2302
rect 478 2168 482 2172
rect 422 2148 426 2152
rect 446 2148 450 2152
rect 462 2148 466 2152
rect 390 2098 394 2102
rect 438 2078 442 2082
rect 398 2068 402 2072
rect 382 2058 386 2062
rect 358 2048 362 2052
rect 318 2038 322 2042
rect 350 2038 354 2042
rect 294 1978 298 1982
rect 270 1958 274 1962
rect 342 1988 346 1992
rect 326 1958 330 1962
rect 318 1948 322 1952
rect 278 1938 282 1942
rect 302 1928 306 1932
rect 262 1908 266 1912
rect 326 1888 330 1892
rect 230 1858 234 1862
rect 254 1859 258 1863
rect 222 1838 226 1842
rect 366 1978 370 1982
rect 398 1978 402 1982
rect 374 1968 378 1972
rect 398 1958 402 1962
rect 382 1938 386 1942
rect 350 1858 354 1862
rect 366 1858 370 1862
rect 382 1908 386 1912
rect 414 1998 418 2002
rect 454 2098 458 2102
rect 422 1958 426 1962
rect 470 2088 474 2092
rect 478 2058 482 2062
rect 462 2048 466 2052
rect 470 2038 474 2042
rect 582 2338 586 2342
rect 542 2248 546 2252
rect 542 2238 546 2242
rect 534 2228 538 2232
rect 498 2203 502 2207
rect 505 2203 509 2207
rect 518 2178 522 2182
rect 654 2448 658 2452
rect 614 2438 618 2442
rect 630 2438 634 2442
rect 718 2548 722 2552
rect 750 2658 754 2662
rect 766 2648 770 2652
rect 750 2638 754 2642
rect 758 2588 762 2592
rect 758 2558 762 2562
rect 798 2598 802 2602
rect 790 2578 794 2582
rect 766 2548 770 2552
rect 742 2518 746 2522
rect 742 2508 746 2512
rect 726 2468 730 2472
rect 718 2368 722 2372
rect 726 2358 730 2362
rect 846 2558 850 2562
rect 838 2548 842 2552
rect 878 2688 882 2692
rect 886 2678 890 2682
rect 902 2668 906 2672
rect 966 2648 970 2652
rect 886 2608 890 2612
rect 862 2578 866 2582
rect 870 2548 874 2552
rect 790 2538 794 2542
rect 822 2538 826 2542
rect 854 2538 858 2542
rect 758 2498 762 2502
rect 758 2478 762 2482
rect 798 2478 802 2482
rect 774 2458 778 2462
rect 646 2348 650 2352
rect 686 2348 690 2352
rect 710 2348 714 2352
rect 742 2348 746 2352
rect 678 2338 682 2342
rect 742 2338 746 2342
rect 646 2278 650 2282
rect 710 2268 714 2272
rect 734 2268 738 2272
rect 726 2258 730 2262
rect 686 2248 690 2252
rect 734 2238 738 2242
rect 598 2188 602 2192
rect 678 2188 682 2192
rect 606 2178 610 2182
rect 574 2168 578 2172
rect 566 2158 570 2162
rect 510 2138 514 2142
rect 726 2138 730 2142
rect 534 2128 538 2132
rect 542 2098 546 2102
rect 558 2098 562 2102
rect 526 2058 530 2062
rect 494 2048 498 2052
rect 526 2048 530 2052
rect 502 2038 506 2042
rect 494 2028 498 2032
rect 486 2018 490 2022
rect 406 1878 410 1882
rect 446 1878 450 1882
rect 498 2003 502 2007
rect 505 2003 509 2007
rect 558 1988 562 1992
rect 526 1968 530 1972
rect 558 1958 562 1962
rect 798 2338 802 2342
rect 838 2518 842 2522
rect 926 2558 930 2562
rect 902 2548 906 2552
rect 918 2548 922 2552
rect 870 2528 874 2532
rect 838 2488 842 2492
rect 862 2488 866 2492
rect 814 2328 818 2332
rect 758 2208 762 2212
rect 846 2478 850 2482
rect 838 2458 842 2462
rect 918 2538 922 2542
rect 942 2538 946 2542
rect 894 2528 898 2532
rect 910 2528 914 2532
rect 886 2488 890 2492
rect 878 2478 882 2482
rect 886 2478 890 2482
rect 878 2468 882 2472
rect 918 2478 922 2482
rect 958 2518 962 2522
rect 1002 2703 1006 2707
rect 1009 2703 1013 2707
rect 1086 2898 1090 2902
rect 1102 2888 1106 2892
rect 1254 3148 1258 3152
rect 1182 2998 1186 3002
rect 1230 2998 1234 3002
rect 1278 2998 1282 3002
rect 1334 3258 1338 3262
rect 1414 3358 1418 3362
rect 1422 3328 1426 3332
rect 1398 3288 1402 3292
rect 1438 3448 1442 3452
rect 1502 3488 1506 3492
rect 1918 3558 1922 3562
rect 1686 3538 1690 3542
rect 1622 3508 1626 3512
rect 1478 3468 1482 3472
rect 1494 3458 1498 3462
rect 1454 3448 1458 3452
rect 1574 3448 1578 3452
rect 1558 3418 1562 3422
rect 1598 3418 1602 3422
rect 1522 3403 1526 3407
rect 1529 3403 1533 3407
rect 1446 3388 1450 3392
rect 1550 3388 1554 3392
rect 1542 3358 1546 3362
rect 1478 3338 1482 3342
rect 1606 3408 1610 3412
rect 1590 3348 1594 3352
rect 1558 3338 1562 3342
rect 1598 3338 1602 3342
rect 1526 3328 1530 3332
rect 1566 3328 1570 3332
rect 1502 3318 1506 3322
rect 1446 3298 1450 3302
rect 1574 3308 1578 3312
rect 1438 3288 1442 3292
rect 1494 3288 1498 3292
rect 1430 3278 1434 3282
rect 1478 3278 1482 3282
rect 1518 3278 1522 3282
rect 1486 3268 1490 3272
rect 1510 3268 1514 3272
rect 1374 3258 1378 3262
rect 1422 3258 1426 3262
rect 1438 3258 1442 3262
rect 1470 3258 1474 3262
rect 1550 3258 1554 3262
rect 1374 3248 1378 3252
rect 1430 3248 1434 3252
rect 1334 3168 1338 3172
rect 1438 3238 1442 3242
rect 1406 3228 1410 3232
rect 1414 3208 1418 3212
rect 1414 3168 1418 3172
rect 1522 3203 1526 3207
rect 1529 3203 1533 3207
rect 1478 3198 1482 3202
rect 1462 3178 1466 3182
rect 1574 3208 1578 3212
rect 1550 3188 1554 3192
rect 1550 3168 1554 3172
rect 1606 3208 1610 3212
rect 1654 3508 1658 3512
rect 1862 3548 1866 3552
rect 1782 3538 1786 3542
rect 1814 3538 1818 3542
rect 1886 3538 1890 3542
rect 1718 3528 1722 3532
rect 1766 3478 1770 3482
rect 1638 3468 1642 3472
rect 1862 3528 1866 3532
rect 1918 3538 1922 3542
rect 1846 3518 1850 3522
rect 1942 3508 1946 3512
rect 1950 3498 1954 3502
rect 1790 3488 1794 3492
rect 1942 3488 1946 3492
rect 1902 3478 1906 3482
rect 1934 3478 1938 3482
rect 1902 3468 1906 3472
rect 1670 3448 1674 3452
rect 1702 3408 1706 3412
rect 1694 3368 1698 3372
rect 1630 3358 1634 3362
rect 1662 3358 1666 3362
rect 1798 3358 1802 3362
rect 1670 3348 1674 3352
rect 1662 3338 1666 3342
rect 1686 3338 1690 3342
rect 1678 3318 1682 3322
rect 1662 3288 1666 3292
rect 1702 3308 1706 3312
rect 1654 3258 1658 3262
rect 1758 3347 1762 3351
rect 1782 3348 1786 3352
rect 1822 3298 1826 3302
rect 1982 3648 1986 3652
rect 2006 3648 2010 3652
rect 2054 3738 2058 3742
rect 2026 3703 2030 3707
rect 2033 3703 2037 3707
rect 2022 3688 2026 3692
rect 2086 3698 2090 3702
rect 2078 3678 2082 3682
rect 2022 3648 2026 3652
rect 2014 3588 2018 3592
rect 2070 3588 2074 3592
rect 2022 3558 2026 3562
rect 1974 3548 1978 3552
rect 1982 3538 1986 3542
rect 1974 3528 1978 3532
rect 1998 3528 2002 3532
rect 2062 3548 2066 3552
rect 2038 3538 2042 3542
rect 2054 3538 2058 3542
rect 2038 3528 2042 3532
rect 2014 3518 2018 3522
rect 2006 3498 2010 3502
rect 1998 3478 2002 3482
rect 1958 3468 1962 3472
rect 1990 3468 1994 3472
rect 1926 3438 1930 3442
rect 1934 3428 1938 3432
rect 1910 3408 1914 3412
rect 1862 3398 1866 3402
rect 1910 3378 1914 3382
rect 1918 3368 1922 3372
rect 1846 3338 1850 3342
rect 1806 3288 1810 3292
rect 1830 3288 1834 3292
rect 1734 3258 1738 3262
rect 1774 3258 1778 3262
rect 1710 3238 1714 3242
rect 1630 3228 1634 3232
rect 1582 3188 1586 3192
rect 1598 3158 1602 3162
rect 1630 3178 1634 3182
rect 1510 3148 1514 3152
rect 1526 3148 1530 3152
rect 1590 3148 1594 3152
rect 1334 3128 1338 3132
rect 1318 3118 1322 3122
rect 1294 3098 1298 3102
rect 1326 3078 1330 3082
rect 1406 3128 1410 3132
rect 1390 3118 1394 3122
rect 1374 3068 1378 3072
rect 1390 3068 1394 3072
rect 1398 3068 1402 3072
rect 1486 3108 1490 3112
rect 1438 3088 1442 3092
rect 1486 3088 1490 3092
rect 1454 3078 1458 3082
rect 1350 3058 1354 3062
rect 1326 3038 1330 3042
rect 1166 2988 1170 2992
rect 1366 2978 1370 2982
rect 1454 3048 1458 3052
rect 1414 3038 1418 3042
rect 1382 3028 1386 3032
rect 1518 3088 1522 3092
rect 1446 2998 1450 3002
rect 1494 2998 1498 3002
rect 1414 2968 1418 2972
rect 1230 2948 1234 2952
rect 1422 2948 1426 2952
rect 1166 2908 1170 2912
rect 1142 2888 1146 2892
rect 1278 2908 1282 2912
rect 1462 2968 1466 2972
rect 1398 2938 1402 2942
rect 1406 2928 1410 2932
rect 1382 2908 1386 2912
rect 1350 2898 1354 2902
rect 1382 2898 1386 2902
rect 1446 2898 1450 2902
rect 1366 2888 1370 2892
rect 1462 2888 1466 2892
rect 1486 2888 1490 2892
rect 1294 2878 1298 2882
rect 1342 2878 1346 2882
rect 1462 2878 1466 2882
rect 1222 2868 1226 2872
rect 1158 2848 1162 2852
rect 1126 2788 1130 2792
rect 1190 2788 1194 2792
rect 1126 2748 1130 2752
rect 1102 2728 1106 2732
rect 1086 2708 1090 2712
rect 1118 2708 1122 2712
rect 1022 2658 1026 2662
rect 1022 2598 1026 2602
rect 1230 2858 1234 2862
rect 1182 2688 1186 2692
rect 1214 2688 1218 2692
rect 1142 2668 1146 2672
rect 1222 2658 1226 2662
rect 1078 2558 1082 2562
rect 1078 2548 1082 2552
rect 990 2538 994 2542
rect 1030 2538 1034 2542
rect 1102 2538 1106 2542
rect 1214 2638 1218 2642
rect 1142 2568 1146 2572
rect 1150 2548 1154 2552
rect 1206 2538 1210 2542
rect 1118 2518 1122 2522
rect 1002 2503 1006 2507
rect 1009 2503 1013 2507
rect 982 2488 986 2492
rect 1046 2488 1050 2492
rect 1102 2488 1106 2492
rect 974 2478 978 2482
rect 1030 2478 1034 2482
rect 1014 2468 1018 2472
rect 926 2458 930 2462
rect 1086 2478 1090 2482
rect 1142 2478 1146 2482
rect 1070 2458 1074 2462
rect 894 2448 898 2452
rect 982 2448 986 2452
rect 862 2428 866 2432
rect 870 2418 874 2422
rect 974 2418 978 2422
rect 870 2388 874 2392
rect 966 2378 970 2382
rect 934 2368 938 2372
rect 918 2358 922 2362
rect 894 2348 898 2352
rect 926 2348 930 2352
rect 950 2348 954 2352
rect 862 2328 866 2332
rect 942 2328 946 2332
rect 958 2328 962 2332
rect 1110 2468 1114 2472
rect 1126 2468 1130 2472
rect 1182 2468 1186 2472
rect 1118 2458 1122 2462
rect 1150 2458 1154 2462
rect 1094 2438 1098 2442
rect 1078 2428 1082 2432
rect 1126 2428 1130 2432
rect 998 2398 1002 2402
rect 998 2378 1002 2382
rect 990 2358 994 2362
rect 998 2358 1002 2362
rect 1014 2358 1018 2362
rect 1014 2338 1018 2342
rect 878 2318 882 2322
rect 830 2308 834 2312
rect 974 2318 978 2322
rect 982 2318 986 2322
rect 886 2298 890 2302
rect 966 2288 970 2292
rect 1002 2303 1006 2307
rect 1009 2303 1013 2307
rect 1062 2358 1066 2362
rect 1062 2338 1066 2342
rect 1158 2368 1162 2372
rect 1094 2338 1098 2342
rect 1142 2338 1146 2342
rect 1190 2338 1194 2342
rect 1078 2318 1082 2322
rect 1086 2288 1090 2292
rect 1102 2288 1106 2292
rect 798 2278 802 2282
rect 958 2278 962 2282
rect 974 2278 978 2282
rect 990 2278 994 2282
rect 1030 2278 1034 2282
rect 878 2268 882 2272
rect 894 2268 898 2272
rect 790 2248 794 2252
rect 822 2178 826 2182
rect 790 2158 794 2162
rect 790 2148 794 2152
rect 678 2128 682 2132
rect 686 2128 690 2132
rect 750 2128 754 2132
rect 686 2108 690 2112
rect 662 2098 666 2102
rect 590 2078 594 2082
rect 694 2078 698 2082
rect 750 2098 754 2102
rect 774 2098 778 2102
rect 782 2088 786 2092
rect 798 2088 802 2092
rect 670 2068 674 2072
rect 814 2068 818 2072
rect 638 2058 642 2062
rect 622 2048 626 2052
rect 654 2048 658 2052
rect 806 2058 810 2062
rect 870 2158 874 2162
rect 878 2158 882 2162
rect 926 2268 930 2272
rect 910 2238 914 2242
rect 950 2238 954 2242
rect 966 2228 970 2232
rect 966 2178 970 2182
rect 846 2148 850 2152
rect 878 2148 882 2152
rect 902 2148 906 2152
rect 838 2138 842 2142
rect 1262 2818 1266 2822
rect 1238 2718 1242 2722
rect 1230 2388 1234 2392
rect 1222 2358 1226 2362
rect 1206 2308 1210 2312
rect 1022 2268 1026 2272
rect 1070 2258 1074 2262
rect 1134 2248 1138 2252
rect 998 2238 1002 2242
rect 1038 2238 1042 2242
rect 1206 2238 1210 2242
rect 1062 2198 1066 2202
rect 1078 2198 1082 2202
rect 1086 2148 1090 2152
rect 1150 2158 1154 2162
rect 1158 2158 1162 2162
rect 1182 2158 1186 2162
rect 1214 2158 1218 2162
rect 1110 2148 1114 2152
rect 1142 2148 1146 2152
rect 1134 2138 1138 2142
rect 830 2128 834 2132
rect 910 2128 914 2132
rect 974 2128 978 2132
rect 990 2128 994 2132
rect 1002 2103 1006 2107
rect 1009 2103 1013 2107
rect 1094 2128 1098 2132
rect 1110 2128 1114 2132
rect 846 2088 850 2092
rect 918 2088 922 2092
rect 982 2088 986 2092
rect 1078 2088 1082 2092
rect 910 2078 914 2082
rect 966 2078 970 2082
rect 1014 2078 1018 2082
rect 1054 2078 1058 2082
rect 1070 2078 1074 2082
rect 1094 2078 1098 2082
rect 838 2068 842 2072
rect 886 2068 890 2072
rect 1038 2068 1042 2072
rect 878 2058 882 2062
rect 990 2058 994 2062
rect 1030 2058 1034 2062
rect 1046 2058 1050 2062
rect 1054 2058 1058 2062
rect 1094 2058 1098 2062
rect 710 2038 714 2042
rect 790 2038 794 2042
rect 798 2038 802 2042
rect 678 2028 682 2032
rect 638 1988 642 1992
rect 694 1988 698 1992
rect 606 1978 610 1982
rect 646 1968 650 1972
rect 630 1958 634 1962
rect 662 1958 666 1962
rect 678 1958 682 1962
rect 510 1948 514 1952
rect 518 1948 522 1952
rect 534 1948 538 1952
rect 590 1948 594 1952
rect 614 1948 618 1952
rect 478 1938 482 1942
rect 534 1938 538 1942
rect 550 1938 554 1942
rect 566 1938 570 1942
rect 582 1938 586 1942
rect 478 1908 482 1912
rect 406 1858 410 1862
rect 398 1848 402 1852
rect 342 1838 346 1842
rect 382 1838 386 1842
rect 310 1828 314 1832
rect 334 1828 338 1832
rect 350 1828 354 1832
rect 302 1788 306 1792
rect 254 1758 258 1762
rect 390 1778 394 1782
rect 318 1768 322 1772
rect 334 1768 338 1772
rect 366 1758 370 1762
rect 246 1748 250 1752
rect 278 1748 282 1752
rect 238 1738 242 1742
rect 254 1738 258 1742
rect 118 1698 122 1702
rect 206 1688 210 1692
rect 198 1678 202 1682
rect 158 1668 162 1672
rect 30 1658 34 1662
rect 54 1658 58 1662
rect 6 1648 10 1652
rect 6 1548 10 1552
rect 22 1538 26 1542
rect 166 1658 170 1662
rect 198 1658 202 1662
rect 118 1648 122 1652
rect 182 1638 186 1642
rect 94 1628 98 1632
rect 166 1618 170 1622
rect 126 1578 130 1582
rect 30 1478 34 1482
rect 126 1468 130 1472
rect 6 1448 10 1452
rect 38 1378 42 1382
rect 22 1368 26 1372
rect 62 1408 66 1412
rect 70 1398 74 1402
rect 54 1378 58 1382
rect 46 1358 50 1362
rect 190 1608 194 1612
rect 174 1548 178 1552
rect 230 1678 234 1682
rect 238 1678 242 1682
rect 214 1668 218 1672
rect 374 1748 378 1752
rect 310 1738 314 1742
rect 262 1728 266 1732
rect 310 1728 314 1732
rect 366 1728 370 1732
rect 254 1718 258 1722
rect 286 1718 290 1722
rect 246 1638 250 1642
rect 238 1608 242 1612
rect 286 1688 290 1692
rect 278 1678 282 1682
rect 286 1678 290 1682
rect 270 1658 274 1662
rect 302 1658 306 1662
rect 318 1708 322 1712
rect 286 1638 290 1642
rect 310 1638 314 1642
rect 294 1608 298 1612
rect 246 1588 250 1592
rect 230 1578 234 1582
rect 230 1558 234 1562
rect 238 1558 242 1562
rect 214 1548 218 1552
rect 206 1498 210 1502
rect 206 1488 210 1492
rect 222 1488 226 1492
rect 230 1488 234 1492
rect 182 1478 186 1482
rect 158 1448 162 1452
rect 150 1388 154 1392
rect 254 1578 258 1582
rect 262 1548 266 1552
rect 302 1548 306 1552
rect 246 1508 250 1512
rect 270 1508 274 1512
rect 254 1488 258 1492
rect 238 1468 242 1472
rect 190 1388 194 1392
rect 142 1378 146 1382
rect 86 1368 90 1372
rect 6 1348 10 1352
rect 54 1348 58 1352
rect 22 1298 26 1302
rect 30 1278 34 1282
rect 174 1358 178 1362
rect 302 1478 306 1482
rect 278 1468 282 1472
rect 350 1688 354 1692
rect 334 1658 338 1662
rect 334 1638 338 1642
rect 390 1678 394 1682
rect 382 1668 386 1672
rect 550 1918 554 1922
rect 438 1848 442 1852
rect 526 1858 530 1862
rect 422 1788 426 1792
rect 430 1747 434 1751
rect 454 1748 458 1752
rect 614 1878 618 1882
rect 582 1868 586 1872
rect 598 1868 602 1872
rect 622 1868 626 1872
rect 638 1868 642 1872
rect 646 1868 650 1872
rect 670 1908 674 1912
rect 702 1968 706 1972
rect 894 2048 898 2052
rect 974 2048 978 2052
rect 982 2048 986 2052
rect 838 2038 842 2042
rect 886 2038 890 2042
rect 822 2008 826 2012
rect 902 1988 906 1992
rect 934 1978 938 1982
rect 1094 1978 1098 1982
rect 790 1968 794 1972
rect 990 1968 994 1972
rect 798 1958 802 1962
rect 1446 2818 1450 2822
rect 1270 2768 1274 2772
rect 1310 2768 1314 2772
rect 1478 2768 1482 2772
rect 1278 2758 1282 2762
rect 1310 2758 1314 2762
rect 1422 2748 1426 2752
rect 1374 2728 1378 2732
rect 1462 2708 1466 2712
rect 1334 2668 1338 2672
rect 1318 2658 1322 2662
rect 1382 2658 1386 2662
rect 1478 2658 1482 2662
rect 1366 2648 1370 2652
rect 1398 2648 1402 2652
rect 1350 2638 1354 2642
rect 1262 2568 1266 2572
rect 1270 2538 1274 2542
rect 1446 2598 1450 2602
rect 1494 2598 1498 2602
rect 1542 3138 1546 3142
rect 1622 3138 1626 3142
rect 1550 3128 1554 3132
rect 1550 3118 1554 3122
rect 1566 3118 1570 3122
rect 1558 3098 1562 3102
rect 1542 3068 1546 3072
rect 1614 3128 1618 3132
rect 1606 3118 1610 3122
rect 1590 3108 1594 3112
rect 1606 3088 1610 3092
rect 1518 3058 1522 3062
rect 1582 3058 1586 3062
rect 1542 3048 1546 3052
rect 1558 3048 1562 3052
rect 1694 3168 1698 3172
rect 1718 3168 1722 3172
rect 1654 3158 1658 3162
rect 1790 3248 1794 3252
rect 1894 3328 1898 3332
rect 1926 3298 1930 3302
rect 1902 3288 1906 3292
rect 1918 3278 1922 3282
rect 1974 3458 1978 3462
rect 2006 3458 2010 3462
rect 1950 3438 1954 3442
rect 1958 3438 1962 3442
rect 1958 3358 1962 3362
rect 1950 3348 1954 3352
rect 1958 3338 1962 3342
rect 1926 3268 1930 3272
rect 1950 3258 1954 3262
rect 1886 3238 1890 3242
rect 1878 3228 1882 3232
rect 1990 3328 1994 3332
rect 2026 3503 2030 3507
rect 2033 3503 2037 3507
rect 2030 3468 2034 3472
rect 2046 3468 2050 3472
rect 2166 3758 2170 3762
rect 2142 3708 2146 3712
rect 2134 3678 2138 3682
rect 2150 3678 2154 3682
rect 2134 3668 2138 3672
rect 2142 3658 2146 3662
rect 2166 3638 2170 3642
rect 2182 3698 2186 3702
rect 2222 3738 2226 3742
rect 2214 3728 2218 3732
rect 2238 3708 2242 3712
rect 2198 3668 2202 3672
rect 2198 3658 2202 3662
rect 2222 3658 2226 3662
rect 2206 3638 2210 3642
rect 2126 3628 2130 3632
rect 2142 3618 2146 3622
rect 2198 3618 2202 3622
rect 2110 3608 2114 3612
rect 2094 3598 2098 3602
rect 2190 3588 2194 3592
rect 2142 3568 2146 3572
rect 2134 3558 2138 3562
rect 2158 3558 2162 3562
rect 2174 3558 2178 3562
rect 2102 3548 2106 3552
rect 2094 3538 2098 3542
rect 2070 3458 2074 3462
rect 2094 3458 2098 3462
rect 2086 3448 2090 3452
rect 2102 3448 2106 3452
rect 2118 3388 2122 3392
rect 2118 3368 2122 3372
rect 2102 3358 2106 3362
rect 2094 3348 2098 3352
rect 2110 3348 2114 3352
rect 2142 3538 2146 3542
rect 2166 3538 2170 3542
rect 2134 3488 2138 3492
rect 2166 3528 2170 3532
rect 2142 3478 2146 3482
rect 2142 3468 2146 3472
rect 2142 3458 2146 3462
rect 2158 3448 2162 3452
rect 2190 3518 2194 3522
rect 2230 3638 2234 3642
rect 2238 3528 2242 3532
rect 2270 3768 2274 3772
rect 2278 3758 2282 3762
rect 2262 3748 2266 3752
rect 2270 3748 2274 3752
rect 2262 3698 2266 3702
rect 2262 3678 2266 3682
rect 2286 3708 2290 3712
rect 2294 3678 2298 3682
rect 2406 3908 2410 3912
rect 2494 3898 2498 3902
rect 2438 3888 2442 3892
rect 2614 4178 2618 4182
rect 2606 4158 2610 4162
rect 2582 4148 2586 4152
rect 2574 4138 2578 4142
rect 2598 4138 2602 4142
rect 2694 4238 2698 4242
rect 2678 4228 2682 4232
rect 2630 4128 2634 4132
rect 2582 4118 2586 4122
rect 2598 4118 2602 4122
rect 2518 4108 2522 4112
rect 2558 4098 2562 4102
rect 2526 4078 2530 4082
rect 2598 4058 2602 4062
rect 2518 4048 2522 4052
rect 2590 4048 2594 4052
rect 2662 4208 2666 4212
rect 2918 4308 2922 4312
rect 2870 4288 2874 4292
rect 2910 4288 2914 4292
rect 2830 4268 2834 4272
rect 2838 4268 2842 4272
rect 2854 4268 2858 4272
rect 2782 4258 2786 4262
rect 2814 4248 2818 4252
rect 2846 4248 2850 4252
rect 2790 4238 2794 4242
rect 2742 4228 2746 4232
rect 2790 4228 2794 4232
rect 2718 4208 2722 4212
rect 2710 4198 2714 4202
rect 2678 4168 2682 4172
rect 2686 4158 2690 4162
rect 2678 4128 2682 4132
rect 2654 4098 2658 4102
rect 2638 4068 2642 4072
rect 2662 4068 2666 4072
rect 2622 4048 2626 4052
rect 2630 4048 2634 4052
rect 2582 4018 2586 4022
rect 2622 4008 2626 4012
rect 2546 4003 2550 4007
rect 2553 4003 2557 4007
rect 2534 3998 2538 4002
rect 2598 3968 2602 3972
rect 2622 3968 2626 3972
rect 2526 3948 2530 3952
rect 2534 3948 2538 3952
rect 2550 3948 2554 3952
rect 2550 3938 2554 3942
rect 2382 3878 2386 3882
rect 2430 3878 2434 3882
rect 2486 3878 2490 3882
rect 2510 3878 2514 3882
rect 2446 3868 2450 3872
rect 2366 3858 2370 3862
rect 2454 3858 2458 3862
rect 2462 3858 2466 3862
rect 2318 3838 2322 3842
rect 2326 3838 2330 3842
rect 2310 3798 2314 3802
rect 2326 3778 2330 3782
rect 2414 3848 2418 3852
rect 2374 3838 2378 3842
rect 2422 3838 2426 3842
rect 2398 3828 2402 3832
rect 2358 3818 2362 3822
rect 2350 3808 2354 3812
rect 2374 3788 2378 3792
rect 2310 3768 2314 3772
rect 2342 3768 2346 3772
rect 2310 3748 2314 3752
rect 2318 3718 2322 3722
rect 2334 3718 2338 3722
rect 2326 3688 2330 3692
rect 2414 3808 2418 3812
rect 2422 3788 2426 3792
rect 2382 3748 2386 3752
rect 2422 3748 2426 3752
rect 2398 3738 2402 3742
rect 2342 3708 2346 3712
rect 2350 3708 2354 3712
rect 2342 3688 2346 3692
rect 2374 3678 2378 3682
rect 2390 3678 2394 3682
rect 2310 3668 2314 3672
rect 2270 3658 2274 3662
rect 2286 3648 2290 3652
rect 2470 3848 2474 3852
rect 2510 3848 2514 3852
rect 2470 3838 2474 3842
rect 2486 3838 2490 3842
rect 2582 3898 2586 3902
rect 2846 4238 2850 4242
rect 2910 4268 2914 4272
rect 2878 4258 2882 4262
rect 2838 4228 2842 4232
rect 2806 4218 2810 4222
rect 2798 4208 2802 4212
rect 2774 4188 2778 4192
rect 2790 4188 2794 4192
rect 2806 4178 2810 4182
rect 2798 4158 2802 4162
rect 2766 4148 2770 4152
rect 2830 4168 2834 4172
rect 2846 4218 2850 4222
rect 2846 4158 2850 4162
rect 2862 4158 2866 4162
rect 2870 4158 2874 4162
rect 2878 4148 2882 4152
rect 2846 4128 2850 4132
rect 2806 4118 2810 4122
rect 2686 4108 2690 4112
rect 2718 4108 2722 4112
rect 2750 4108 2754 4112
rect 2734 4078 2738 4082
rect 2750 4068 2754 4072
rect 2878 4118 2882 4122
rect 2934 4308 2938 4312
rect 2950 4298 2954 4302
rect 2926 4278 2930 4282
rect 2934 4268 2938 4272
rect 2918 4228 2922 4232
rect 2894 4208 2898 4212
rect 2926 4208 2930 4212
rect 2982 4298 2986 4302
rect 2990 4288 2994 4292
rect 2958 4278 2962 4282
rect 2950 4258 2954 4262
rect 3038 4308 3042 4312
rect 3050 4303 3054 4307
rect 3057 4303 3061 4307
rect 3230 4338 3234 4342
rect 3086 4298 3090 4302
rect 3278 4348 3282 4352
rect 3422 4348 3426 4352
rect 3438 4348 3442 4352
rect 3478 4348 3482 4352
rect 3494 4348 3498 4352
rect 3518 4348 3522 4352
rect 3558 4348 3562 4352
rect 3670 4368 3674 4372
rect 3638 4358 3642 4362
rect 3790 4398 3794 4402
rect 3806 4398 3810 4402
rect 3830 4398 3834 4402
rect 3766 4378 3770 4382
rect 3718 4358 3722 4362
rect 3750 4358 3754 4362
rect 3862 4388 3866 4392
rect 3814 4358 3818 4362
rect 3742 4348 3746 4352
rect 3758 4348 3762 4352
rect 3790 4348 3794 4352
rect 3822 4348 3826 4352
rect 3870 4348 3874 4352
rect 3262 4338 3266 4342
rect 3246 4318 3250 4322
rect 3238 4308 3242 4312
rect 3302 4318 3306 4322
rect 3358 4338 3362 4342
rect 3366 4328 3370 4332
rect 3262 4298 3266 4302
rect 3270 4298 3274 4302
rect 3334 4298 3338 4302
rect 3094 4288 3098 4292
rect 3230 4288 3234 4292
rect 3358 4288 3362 4292
rect 3390 4288 3394 4292
rect 3126 4278 3130 4282
rect 3142 4278 3146 4282
rect 3326 4278 3330 4282
rect 3014 4268 3018 4272
rect 3078 4268 3082 4272
rect 2950 4248 2954 4252
rect 2982 4248 2986 4252
rect 3046 4248 3050 4252
rect 2966 4238 2970 4242
rect 2942 4228 2946 4232
rect 3054 4218 3058 4222
rect 2950 4198 2954 4202
rect 2934 4158 2938 4162
rect 2942 4158 2946 4162
rect 2902 4148 2906 4152
rect 2942 4148 2946 4152
rect 2894 4128 2898 4132
rect 2910 4128 2914 4132
rect 2942 4098 2946 4102
rect 2910 4088 2914 4092
rect 2886 4078 2890 4082
rect 2774 4058 2778 4062
rect 2814 4058 2818 4062
rect 2822 4058 2826 4062
rect 2886 4058 2890 4062
rect 2918 4058 2922 4062
rect 2694 4048 2698 4052
rect 2710 4048 2714 4052
rect 2758 4048 2762 4052
rect 2782 4048 2786 4052
rect 2742 4038 2746 4042
rect 2782 4038 2786 4042
rect 2678 4028 2682 4032
rect 2718 4028 2722 4032
rect 2750 4028 2754 4032
rect 2806 4038 2810 4042
rect 2838 4038 2842 4042
rect 2702 4018 2706 4022
rect 2670 3998 2674 4002
rect 2686 3968 2690 3972
rect 2646 3958 2650 3962
rect 2614 3938 2618 3942
rect 2662 3928 2666 3932
rect 2694 3948 2698 3952
rect 2630 3918 2634 3922
rect 2670 3918 2674 3922
rect 2574 3888 2578 3892
rect 2606 3888 2610 3892
rect 2598 3858 2602 3862
rect 2558 3848 2562 3852
rect 2518 3828 2522 3832
rect 2542 3828 2546 3832
rect 2486 3808 2490 3812
rect 2446 3728 2450 3732
rect 2462 3678 2466 3682
rect 2430 3668 2434 3672
rect 2390 3658 2394 3662
rect 2406 3658 2410 3662
rect 2438 3658 2442 3662
rect 2302 3648 2306 3652
rect 2326 3648 2330 3652
rect 2350 3648 2354 3652
rect 2262 3638 2266 3642
rect 2286 3628 2290 3632
rect 2286 3608 2290 3612
rect 2246 3508 2250 3512
rect 2246 3498 2250 3502
rect 2190 3478 2194 3482
rect 2198 3478 2202 3482
rect 2214 3478 2218 3482
rect 2174 3468 2178 3472
rect 2150 3378 2154 3382
rect 2142 3368 2146 3372
rect 2190 3438 2194 3442
rect 2310 3588 2314 3592
rect 2302 3538 2306 3542
rect 2318 3538 2322 3542
rect 2278 3528 2282 3532
rect 2262 3488 2266 3492
rect 2334 3638 2338 3642
rect 2262 3468 2266 3472
rect 2302 3468 2306 3472
rect 2206 3448 2210 3452
rect 2230 3448 2234 3452
rect 2254 3448 2258 3452
rect 2238 3438 2242 3442
rect 2198 3428 2202 3432
rect 2206 3428 2210 3432
rect 2238 3428 2242 3432
rect 2294 3458 2298 3462
rect 2294 3448 2298 3452
rect 2278 3388 2282 3392
rect 2254 3368 2258 3372
rect 2262 3368 2266 3372
rect 2318 3448 2322 3452
rect 2382 3638 2386 3642
rect 2406 3638 2410 3642
rect 2366 3628 2370 3632
rect 2430 3588 2434 3592
rect 2454 3658 2458 3662
rect 2546 3803 2550 3807
rect 2553 3803 2557 3807
rect 2518 3768 2522 3772
rect 2534 3758 2538 3762
rect 2510 3748 2514 3752
rect 2534 3748 2538 3752
rect 2646 3888 2650 3892
rect 2686 3908 2690 3912
rect 2702 3908 2706 3912
rect 2662 3858 2666 3862
rect 2678 3858 2682 3862
rect 2638 3848 2642 3852
rect 2598 3838 2602 3842
rect 2678 3838 2682 3842
rect 2614 3828 2618 3832
rect 2646 3828 2650 3832
rect 2622 3808 2626 3812
rect 2670 3798 2674 3802
rect 2598 3768 2602 3772
rect 2606 3768 2610 3772
rect 2590 3748 2594 3752
rect 2494 3738 2498 3742
rect 2518 3738 2522 3742
rect 2542 3738 2546 3742
rect 2574 3738 2578 3742
rect 2494 3668 2498 3672
rect 2478 3648 2482 3652
rect 2478 3638 2482 3642
rect 2470 3628 2474 3632
rect 2470 3608 2474 3612
rect 2446 3578 2450 3582
rect 2462 3578 2466 3582
rect 2462 3568 2466 3572
rect 2446 3558 2450 3562
rect 2374 3547 2378 3551
rect 2422 3538 2426 3542
rect 2430 3538 2434 3542
rect 2382 3528 2386 3532
rect 2414 3528 2418 3532
rect 2366 3498 2370 3502
rect 2350 3478 2354 3482
rect 2366 3478 2370 3482
rect 2342 3458 2346 3462
rect 2374 3468 2378 3472
rect 2382 3448 2386 3452
rect 2334 3438 2338 3442
rect 2366 3368 2370 3372
rect 2134 3358 2138 3362
rect 2166 3358 2170 3362
rect 2174 3358 2178 3362
rect 2230 3358 2234 3362
rect 2310 3358 2314 3362
rect 2102 3338 2106 3342
rect 2118 3338 2122 3342
rect 2182 3348 2186 3352
rect 2198 3348 2202 3352
rect 2190 3338 2194 3342
rect 2022 3328 2026 3332
rect 2054 3328 2058 3332
rect 2110 3328 2114 3332
rect 2026 3303 2030 3307
rect 2033 3303 2037 3307
rect 2054 3298 2058 3302
rect 2022 3288 2026 3292
rect 2094 3288 2098 3292
rect 2062 3268 2066 3272
rect 2094 3248 2098 3252
rect 1982 3208 1986 3212
rect 1950 3198 1954 3202
rect 1974 3198 1978 3202
rect 1838 3168 1842 3172
rect 1806 3158 1810 3162
rect 1918 3158 1922 3162
rect 1654 3148 1658 3152
rect 1694 3148 1698 3152
rect 1726 3148 1730 3152
rect 1646 3118 1650 3122
rect 1686 3108 1690 3112
rect 1718 3108 1722 3112
rect 1694 3098 1698 3102
rect 1678 3078 1682 3082
rect 2070 3168 2074 3172
rect 2086 3158 2090 3162
rect 2126 3298 2130 3302
rect 2166 3298 2170 3302
rect 2142 3208 2146 3212
rect 2190 3288 2194 3292
rect 2174 3278 2178 3282
rect 2142 3178 2146 3182
rect 2006 3147 2010 3151
rect 2086 3138 2090 3142
rect 2102 3138 2106 3142
rect 1990 3128 1994 3132
rect 2094 3128 2098 3132
rect 1790 3098 1794 3102
rect 1878 3088 1882 3092
rect 1990 3088 1994 3092
rect 2026 3103 2030 3107
rect 2033 3103 2037 3107
rect 1726 3068 1730 3072
rect 1758 3068 1762 3072
rect 1846 3059 1850 3063
rect 1638 3048 1642 3052
rect 1846 3048 1850 3052
rect 1758 3028 1762 3032
rect 1662 3008 1666 3012
rect 1522 3003 1526 3007
rect 1529 3003 1533 3007
rect 1662 2978 1666 2982
rect 1526 2947 1530 2951
rect 1550 2948 1554 2952
rect 1814 2968 1818 2972
rect 1854 2998 1858 3002
rect 1902 2968 1906 2972
rect 1678 2938 1682 2942
rect 1734 2938 1738 2942
rect 1662 2928 1666 2932
rect 1574 2898 1578 2902
rect 1590 2898 1594 2902
rect 1630 2898 1634 2902
rect 1550 2868 1554 2872
rect 1522 2803 1526 2807
rect 1529 2803 1533 2807
rect 1518 2768 1522 2772
rect 1558 2848 1562 2852
rect 1558 2698 1562 2702
rect 1670 2908 1674 2912
rect 1662 2888 1666 2892
rect 1590 2878 1594 2882
rect 1598 2868 1602 2872
rect 1654 2868 1658 2872
rect 1694 2908 1698 2912
rect 1790 2888 1794 2892
rect 1774 2878 1778 2882
rect 1766 2868 1770 2872
rect 1622 2858 1626 2862
rect 1646 2858 1650 2862
rect 1726 2858 1730 2862
rect 1622 2848 1626 2852
rect 1654 2848 1658 2852
rect 1678 2768 1682 2772
rect 1614 2758 1618 2762
rect 1598 2748 1602 2752
rect 1662 2748 1666 2752
rect 1582 2738 1586 2742
rect 1590 2728 1594 2732
rect 1590 2688 1594 2692
rect 1574 2668 1578 2672
rect 1614 2678 1618 2682
rect 1654 2678 1658 2682
rect 1622 2668 1626 2672
rect 1694 2758 1698 2762
rect 1678 2718 1682 2722
rect 1670 2698 1674 2702
rect 1646 2658 1650 2662
rect 1646 2648 1650 2652
rect 1522 2603 1526 2607
rect 1529 2603 1533 2607
rect 1462 2588 1466 2592
rect 1502 2588 1506 2592
rect 1558 2588 1562 2592
rect 1662 2578 1666 2582
rect 1542 2568 1546 2572
rect 1598 2568 1602 2572
rect 1294 2468 1298 2472
rect 1302 2468 1306 2472
rect 1254 2438 1258 2442
rect 1326 2368 1330 2372
rect 1254 2358 1258 2362
rect 1262 2348 1266 2352
rect 1262 2338 1266 2342
rect 1374 2478 1378 2482
rect 1390 2448 1394 2452
rect 1518 2508 1522 2512
rect 1518 2498 1522 2502
rect 1462 2488 1466 2492
rect 1486 2488 1490 2492
rect 1470 2478 1474 2482
rect 1406 2428 1410 2432
rect 1422 2418 1426 2422
rect 1406 2358 1410 2362
rect 1630 2528 1634 2532
rect 1646 2498 1650 2502
rect 1494 2458 1498 2462
rect 1510 2458 1514 2462
rect 1534 2458 1538 2462
rect 1542 2448 1546 2452
rect 1522 2403 1526 2407
rect 1529 2403 1533 2407
rect 1550 2408 1554 2412
rect 1446 2348 1450 2352
rect 1358 2338 1362 2342
rect 1382 2338 1386 2342
rect 1374 2298 1378 2302
rect 1350 2288 1354 2292
rect 1318 2278 1322 2282
rect 1382 2278 1386 2282
rect 1398 2268 1402 2272
rect 1238 2258 1242 2262
rect 1278 2228 1282 2232
rect 1246 2168 1250 2172
rect 1198 2138 1202 2142
rect 1222 2138 1226 2142
rect 1158 2128 1162 2132
rect 1206 2128 1210 2132
rect 1222 2078 1226 2082
rect 1230 2078 1234 2082
rect 1134 2048 1138 2052
rect 1174 2068 1178 2072
rect 1206 2068 1210 2072
rect 1438 2308 1442 2312
rect 1438 2298 1442 2302
rect 1470 2288 1474 2292
rect 1486 2298 1490 2302
rect 1630 2458 1634 2462
rect 1606 2438 1610 2442
rect 1734 2848 1738 2852
rect 1726 2748 1730 2752
rect 1734 2738 1738 2742
rect 1758 2848 1762 2852
rect 1758 2768 1762 2772
rect 1750 2758 1754 2762
rect 1846 2898 1850 2902
rect 1830 2888 1834 2892
rect 1838 2888 1842 2892
rect 1806 2878 1810 2882
rect 1822 2878 1826 2882
rect 1830 2868 1834 2872
rect 1846 2868 1850 2872
rect 1798 2858 1802 2862
rect 1798 2778 1802 2782
rect 1790 2758 1794 2762
rect 1774 2748 1778 2752
rect 1806 2758 1810 2762
rect 1950 3048 1954 3052
rect 2038 3059 2042 3063
rect 2238 3348 2242 3352
rect 2214 3308 2218 3312
rect 2222 3258 2226 3262
rect 2286 3348 2290 3352
rect 2302 3348 2306 3352
rect 2334 3348 2338 3352
rect 2342 3338 2346 3342
rect 2254 3318 2258 3322
rect 2278 3318 2282 3322
rect 2278 3308 2282 3312
rect 2294 3288 2298 3292
rect 2246 3268 2250 3272
rect 2254 3258 2258 3262
rect 2222 3248 2226 3252
rect 2206 3228 2210 3232
rect 2214 3228 2218 3232
rect 2206 3198 2210 3202
rect 2190 3188 2194 3192
rect 2166 3168 2170 3172
rect 2174 3168 2178 3172
rect 2206 3168 2210 3172
rect 2166 3138 2170 3142
rect 2174 3138 2178 3142
rect 2150 3128 2154 3132
rect 2158 3128 2162 3132
rect 2182 3128 2186 3132
rect 2142 3108 2146 3112
rect 2126 3098 2130 3102
rect 2078 3068 2082 3072
rect 2110 3058 2114 3062
rect 2062 3028 2066 3032
rect 2118 3018 2122 3022
rect 2190 3118 2194 3122
rect 2174 3108 2178 3112
rect 2150 3078 2154 3082
rect 2158 3068 2162 3072
rect 2246 3208 2250 3212
rect 2230 3178 2234 3182
rect 2230 3168 2234 3172
rect 2238 3088 2242 3092
rect 2182 3078 2186 3082
rect 2214 3078 2218 3082
rect 2174 3058 2178 3062
rect 2198 3058 2202 3062
rect 2134 2998 2138 3002
rect 2198 3048 2202 3052
rect 2214 3048 2218 3052
rect 2166 3038 2170 3042
rect 2158 3028 2162 3032
rect 2166 2998 2170 3002
rect 2190 2998 2194 3002
rect 2134 2948 2138 2952
rect 2014 2938 2018 2942
rect 2062 2938 2066 2942
rect 2118 2938 2122 2942
rect 2238 3028 2242 3032
rect 2254 3168 2258 3172
rect 2262 3148 2266 3152
rect 2262 3098 2266 3102
rect 2254 3088 2258 3092
rect 2254 3078 2258 3082
rect 2246 3018 2250 3022
rect 2262 2978 2266 2982
rect 2262 2968 2266 2972
rect 2222 2947 2226 2951
rect 2310 3198 2314 3202
rect 2358 3328 2362 3332
rect 2366 3328 2370 3332
rect 2414 3498 2418 3502
rect 2422 3488 2426 3492
rect 2566 3698 2570 3702
rect 2542 3668 2546 3672
rect 2590 3678 2594 3682
rect 2590 3658 2594 3662
rect 2550 3648 2554 3652
rect 2526 3638 2530 3642
rect 2518 3628 2522 3632
rect 2494 3608 2498 3612
rect 2546 3603 2550 3607
rect 2553 3603 2557 3607
rect 2518 3598 2522 3602
rect 2486 3588 2490 3592
rect 2486 3578 2490 3582
rect 2494 3568 2498 3572
rect 2510 3568 2514 3572
rect 2534 3568 2538 3572
rect 2446 3538 2450 3542
rect 2478 3538 2482 3542
rect 2526 3538 2530 3542
rect 2542 3538 2546 3542
rect 2558 3538 2562 3542
rect 2486 3528 2490 3532
rect 2478 3518 2482 3522
rect 2438 3478 2442 3482
rect 2502 3478 2506 3482
rect 2430 3468 2434 3472
rect 2454 3468 2458 3472
rect 2414 3428 2418 3432
rect 2398 3388 2402 3392
rect 2390 3348 2394 3352
rect 2374 3318 2378 3322
rect 2358 3298 2362 3302
rect 2390 3308 2394 3312
rect 2382 3288 2386 3292
rect 2406 3278 2410 3282
rect 2390 3248 2394 3252
rect 2446 3458 2450 3462
rect 2478 3448 2482 3452
rect 2798 4008 2802 4012
rect 2790 3978 2794 3982
rect 2830 3978 2834 3982
rect 2822 3968 2826 3972
rect 2734 3958 2738 3962
rect 2806 3958 2810 3962
rect 2718 3928 2722 3932
rect 2782 3948 2786 3952
rect 2838 3948 2842 3952
rect 2814 3938 2818 3942
rect 2742 3928 2746 3932
rect 2758 3928 2762 3932
rect 2774 3928 2778 3932
rect 2798 3928 2802 3932
rect 2830 3928 2834 3932
rect 2734 3918 2738 3922
rect 2710 3898 2714 3902
rect 2718 3898 2722 3902
rect 2702 3868 2706 3872
rect 2702 3858 2706 3862
rect 2702 3788 2706 3792
rect 2726 3878 2730 3882
rect 2718 3858 2722 3862
rect 2710 3778 2714 3782
rect 2718 3758 2722 3762
rect 2574 3648 2578 3652
rect 2598 3648 2602 3652
rect 2566 3478 2570 3482
rect 2526 3468 2530 3472
rect 2526 3458 2530 3462
rect 2470 3438 2474 3442
rect 2486 3438 2490 3442
rect 2494 3418 2498 3422
rect 2438 3368 2442 3372
rect 2438 3358 2442 3362
rect 2486 3358 2490 3362
rect 2422 3268 2426 3272
rect 2478 3348 2482 3352
rect 2446 3338 2450 3342
rect 2462 3298 2466 3302
rect 2518 3438 2522 3442
rect 2546 3403 2550 3407
rect 2553 3403 2557 3407
rect 2510 3398 2514 3402
rect 2550 3388 2554 3392
rect 2526 3368 2530 3372
rect 2622 3688 2626 3692
rect 2694 3748 2698 3752
rect 2686 3678 2690 3682
rect 2654 3668 2658 3672
rect 2678 3668 2682 3672
rect 2750 3868 2754 3872
rect 2742 3858 2746 3862
rect 2742 3788 2746 3792
rect 2774 3848 2778 3852
rect 2790 3838 2794 3842
rect 2862 4048 2866 4052
rect 2894 4048 2898 4052
rect 2910 4038 2914 4042
rect 2894 3998 2898 4002
rect 2862 3958 2866 3962
rect 2886 3958 2890 3962
rect 2854 3928 2858 3932
rect 2846 3908 2850 3912
rect 2822 3898 2826 3902
rect 2766 3788 2770 3792
rect 2758 3768 2762 3772
rect 2774 3758 2778 3762
rect 2726 3688 2730 3692
rect 2638 3658 2642 3662
rect 2662 3658 2666 3662
rect 2702 3658 2706 3662
rect 2630 3648 2634 3652
rect 2606 3628 2610 3632
rect 2646 3638 2650 3642
rect 2702 3638 2706 3642
rect 2686 3628 2690 3632
rect 2646 3568 2650 3572
rect 2662 3588 2666 3592
rect 2654 3548 2658 3552
rect 2606 3538 2610 3542
rect 2582 3478 2586 3482
rect 2574 3438 2578 3442
rect 2622 3468 2626 3472
rect 2598 3458 2602 3462
rect 2630 3458 2634 3462
rect 2622 3448 2626 3452
rect 2614 3438 2618 3442
rect 2622 3438 2626 3442
rect 2654 3508 2658 3512
rect 2670 3548 2674 3552
rect 2694 3598 2698 3602
rect 2726 3658 2730 3662
rect 2742 3708 2746 3712
rect 2750 3668 2754 3672
rect 2758 3668 2762 3672
rect 2774 3668 2778 3672
rect 2742 3658 2746 3662
rect 2774 3648 2778 3652
rect 2742 3638 2746 3642
rect 2734 3628 2738 3632
rect 2726 3618 2730 3622
rect 2710 3568 2714 3572
rect 2678 3538 2682 3542
rect 2686 3528 2690 3532
rect 2710 3518 2714 3522
rect 2694 3488 2698 3492
rect 2662 3478 2666 3482
rect 2686 3468 2690 3472
rect 2726 3468 2730 3472
rect 2662 3458 2666 3462
rect 2694 3458 2698 3462
rect 2798 3808 2802 3812
rect 2838 3868 2842 3872
rect 2846 3858 2850 3862
rect 2886 3898 2890 3902
rect 2878 3868 2882 3872
rect 2934 4038 2938 4042
rect 2926 4018 2930 4022
rect 2918 3988 2922 3992
rect 2934 3947 2938 3951
rect 2918 3908 2922 3912
rect 2910 3898 2914 3902
rect 2894 3858 2898 3862
rect 2910 3878 2914 3882
rect 2942 3868 2946 3872
rect 2854 3848 2858 3852
rect 2870 3848 2874 3852
rect 2902 3848 2906 3852
rect 2830 3838 2834 3842
rect 2846 3828 2850 3832
rect 2814 3788 2818 3792
rect 2806 3768 2810 3772
rect 2806 3758 2810 3762
rect 2854 3798 2858 3802
rect 2862 3788 2866 3792
rect 2878 3788 2882 3792
rect 2862 3778 2866 3782
rect 2990 4168 2994 4172
rect 3022 4148 3026 4152
rect 2998 4138 3002 4142
rect 2966 4098 2970 4102
rect 2990 4058 2994 4062
rect 3174 4268 3178 4272
rect 3102 4258 3106 4262
rect 3118 4178 3122 4182
rect 3142 4168 3146 4172
rect 3134 4148 3138 4152
rect 3150 4148 3154 4152
rect 3038 4138 3042 4142
rect 3190 4138 3194 4142
rect 3038 4128 3042 4132
rect 3078 4118 3082 4122
rect 3050 4103 3054 4107
rect 3057 4103 3061 4107
rect 3070 4098 3074 4102
rect 3086 4078 3090 4082
rect 3070 4058 3074 4062
rect 3046 4048 3050 4052
rect 3246 4198 3250 4202
rect 3246 4178 3250 4182
rect 3230 4168 3234 4172
rect 3470 4338 3474 4342
rect 3486 4338 3490 4342
rect 3446 4318 3450 4322
rect 3446 4298 3450 4302
rect 3398 4278 3402 4282
rect 3430 4278 3434 4282
rect 3438 4278 3442 4282
rect 3366 4268 3370 4272
rect 3286 4258 3290 4262
rect 3310 4258 3314 4262
rect 3358 4258 3362 4262
rect 3278 4228 3282 4232
rect 3262 4218 3266 4222
rect 3222 4148 3226 4152
rect 3214 4138 3218 4142
rect 3166 4128 3170 4132
rect 3198 4128 3202 4132
rect 3102 4098 3106 4102
rect 3174 4088 3178 4092
rect 3126 4058 3130 4062
rect 3182 4058 3186 4062
rect 3206 4058 3210 4062
rect 2998 3988 3002 3992
rect 3038 3988 3042 3992
rect 3086 3988 3090 3992
rect 3094 3988 3098 3992
rect 3022 3968 3026 3972
rect 3142 3968 3146 3972
rect 3126 3928 3130 3932
rect 3050 3903 3054 3907
rect 3057 3903 3061 3907
rect 3006 3898 3010 3902
rect 3126 3898 3130 3902
rect 3142 3898 3146 3902
rect 3006 3888 3010 3892
rect 3030 3888 3034 3892
rect 3110 3888 3114 3892
rect 3022 3868 3026 3872
rect 2982 3858 2986 3862
rect 3038 3868 3042 3872
rect 3102 3868 3106 3872
rect 3046 3848 3050 3852
rect 3070 3848 3074 3852
rect 3014 3838 3018 3842
rect 3062 3838 3066 3842
rect 3006 3828 3010 3832
rect 2958 3768 2962 3772
rect 2886 3758 2890 3762
rect 2934 3758 2938 3762
rect 2846 3748 2850 3752
rect 2878 3748 2882 3752
rect 2934 3748 2938 3752
rect 3014 3778 3018 3782
rect 3022 3768 3026 3772
rect 2982 3758 2986 3762
rect 3006 3758 3010 3762
rect 3014 3748 3018 3752
rect 2790 3738 2794 3742
rect 2830 3738 2834 3742
rect 2918 3738 2922 3742
rect 3014 3738 3018 3742
rect 2822 3728 2826 3732
rect 2886 3728 2890 3732
rect 2910 3728 2914 3732
rect 2926 3728 2930 3732
rect 2942 3728 2946 3732
rect 2798 3718 2802 3722
rect 2862 3708 2866 3712
rect 2902 3708 2906 3712
rect 2926 3708 2930 3712
rect 2806 3698 2810 3702
rect 2806 3678 2810 3682
rect 2854 3678 2858 3682
rect 2798 3658 2802 3662
rect 2830 3668 2834 3672
rect 2846 3668 2850 3672
rect 2790 3638 2794 3642
rect 2814 3638 2818 3642
rect 2782 3568 2786 3572
rect 2766 3548 2770 3552
rect 2782 3548 2786 3552
rect 2830 3638 2834 3642
rect 2822 3628 2826 3632
rect 2838 3618 2842 3622
rect 2902 3688 2906 3692
rect 2886 3678 2890 3682
rect 2910 3668 2914 3672
rect 2870 3648 2874 3652
rect 2942 3698 2946 3702
rect 3038 3728 3042 3732
rect 2998 3718 3002 3722
rect 2966 3678 2970 3682
rect 3050 3703 3054 3707
rect 3057 3703 3061 3707
rect 3014 3688 3018 3692
rect 3062 3678 3066 3682
rect 2990 3668 2994 3672
rect 2950 3658 2954 3662
rect 2942 3648 2946 3652
rect 2966 3638 2970 3642
rect 2862 3578 2866 3582
rect 2854 3568 2858 3572
rect 2806 3558 2810 3562
rect 2838 3548 2842 3552
rect 2806 3518 2810 3522
rect 2670 3448 2674 3452
rect 2734 3448 2738 3452
rect 2654 3438 2658 3442
rect 2694 3438 2698 3442
rect 2606 3388 2610 3392
rect 2646 3388 2650 3392
rect 2630 3378 2634 3382
rect 2566 3368 2570 3372
rect 2606 3368 2610 3372
rect 2614 3368 2618 3372
rect 2582 3358 2586 3362
rect 2510 3298 2514 3302
rect 2558 3328 2562 3332
rect 2550 3308 2554 3312
rect 2470 3288 2474 3292
rect 2462 3268 2466 3272
rect 2470 3268 2474 3272
rect 2566 3268 2570 3272
rect 2414 3248 2418 3252
rect 2470 3248 2474 3252
rect 2414 3238 2418 3242
rect 2454 3238 2458 3242
rect 2678 3408 2682 3412
rect 2670 3388 2674 3392
rect 2654 3378 2658 3382
rect 2598 3348 2602 3352
rect 2606 3348 2610 3352
rect 2726 3438 2730 3442
rect 2734 3398 2738 3402
rect 2782 3498 2786 3502
rect 2798 3458 2802 3462
rect 2822 3508 2826 3512
rect 2862 3508 2866 3512
rect 2830 3478 2834 3482
rect 2822 3468 2826 3472
rect 2838 3468 2842 3472
rect 2782 3448 2786 3452
rect 2814 3448 2818 3452
rect 2846 3448 2850 3452
rect 2854 3448 2858 3452
rect 2806 3438 2810 3442
rect 2758 3408 2762 3412
rect 2822 3398 2826 3402
rect 2782 3388 2786 3392
rect 2750 3378 2754 3382
rect 2742 3368 2746 3372
rect 2774 3368 2778 3372
rect 2782 3358 2786 3362
rect 2734 3348 2738 3352
rect 2886 3568 2890 3572
rect 2886 3548 2890 3552
rect 2918 3538 2922 3542
rect 2918 3508 2922 3512
rect 2926 3498 2930 3502
rect 2910 3488 2914 3492
rect 2894 3478 2898 3482
rect 2878 3468 2882 3472
rect 2870 3458 2874 3462
rect 2902 3468 2906 3472
rect 2990 3598 2994 3602
rect 2950 3578 2954 3582
rect 2974 3578 2978 3582
rect 2982 3578 2986 3582
rect 2998 3578 3002 3582
rect 2966 3538 2970 3542
rect 2942 3518 2946 3522
rect 2966 3518 2970 3522
rect 2934 3468 2938 3472
rect 2910 3458 2914 3462
rect 2926 3458 2930 3462
rect 2966 3458 2970 3462
rect 2894 3448 2898 3452
rect 2918 3448 2922 3452
rect 2878 3438 2882 3442
rect 2942 3448 2946 3452
rect 3014 3628 3018 3632
rect 3022 3608 3026 3612
rect 3038 3648 3042 3652
rect 3118 3868 3122 3872
rect 3230 4128 3234 4132
rect 3278 4178 3282 4182
rect 3270 4158 3274 4162
rect 3294 4248 3298 4252
rect 3334 4248 3338 4252
rect 3302 4238 3306 4242
rect 3326 4238 3330 4242
rect 3358 4238 3362 4242
rect 3310 4218 3314 4222
rect 3302 4178 3306 4182
rect 3286 4168 3290 4172
rect 3302 4148 3306 4152
rect 3270 4138 3274 4142
rect 3286 4138 3290 4142
rect 3302 4138 3306 4142
rect 3230 4078 3234 4082
rect 3238 4068 3242 4072
rect 3222 4048 3226 4052
rect 3198 4038 3202 4042
rect 3222 4038 3226 4042
rect 3214 3998 3218 4002
rect 3206 3938 3210 3942
rect 3142 3888 3146 3892
rect 3086 3828 3090 3832
rect 3126 3758 3130 3762
rect 3094 3748 3098 3752
rect 3118 3748 3122 3752
rect 3142 3748 3146 3752
rect 3150 3748 3154 3752
rect 3166 3748 3170 3752
rect 3198 3748 3202 3752
rect 3262 4068 3266 4072
rect 3254 4058 3258 4062
rect 3262 4048 3266 4052
rect 3310 4128 3314 4132
rect 3302 4108 3306 4112
rect 3358 4188 3362 4192
rect 3454 4268 3458 4272
rect 3406 4258 3410 4262
rect 3374 4248 3378 4252
rect 3382 4238 3386 4242
rect 3398 4238 3402 4242
rect 3374 4218 3378 4222
rect 3350 4158 3354 4162
rect 3326 4148 3330 4152
rect 3350 4148 3354 4152
rect 3334 4108 3338 4112
rect 3374 4138 3378 4142
rect 3366 4088 3370 4092
rect 3302 4068 3306 4072
rect 3278 4058 3282 4062
rect 3222 3938 3226 3942
rect 3270 3948 3274 3952
rect 3286 3948 3290 3952
rect 3326 4058 3330 4062
rect 3318 4048 3322 4052
rect 3310 4038 3314 4042
rect 3334 3968 3338 3972
rect 3422 4228 3426 4232
rect 3462 4228 3466 4232
rect 3446 4208 3450 4212
rect 3502 4328 3506 4332
rect 3478 4308 3482 4312
rect 3486 4298 3490 4302
rect 3518 4298 3522 4302
rect 3542 4308 3546 4312
rect 3486 4268 3490 4272
rect 3502 4258 3506 4262
rect 3478 4248 3482 4252
rect 3502 4248 3506 4252
rect 3478 4238 3482 4242
rect 3510 4218 3514 4222
rect 3510 4208 3514 4212
rect 3494 4178 3498 4182
rect 3414 4158 3418 4162
rect 3446 4158 3450 4162
rect 3638 4338 3642 4342
rect 3646 4328 3650 4332
rect 3614 4318 3618 4322
rect 3630 4318 3634 4322
rect 3598 4298 3602 4302
rect 3598 4288 3602 4292
rect 3630 4288 3634 4292
rect 3702 4338 3706 4342
rect 3662 4328 3666 4332
rect 3726 4328 3730 4332
rect 3710 4308 3714 4312
rect 3686 4298 3690 4302
rect 3670 4288 3674 4292
rect 3678 4288 3682 4292
rect 3654 4278 3658 4282
rect 3622 4268 3626 4272
rect 3654 4268 3658 4272
rect 3638 4258 3642 4262
rect 3534 4248 3538 4252
rect 3606 4248 3610 4252
rect 3526 4158 3530 4162
rect 3570 4203 3574 4207
rect 3577 4203 3581 4207
rect 3638 4168 3642 4172
rect 3494 4148 3498 4152
rect 3558 4148 3562 4152
rect 3438 4138 3442 4142
rect 3422 4128 3426 4132
rect 3438 4118 3442 4122
rect 3454 4138 3458 4142
rect 3470 4138 3474 4142
rect 3486 4118 3490 4122
rect 3446 4078 3450 4082
rect 3478 4078 3482 4082
rect 3454 4068 3458 4072
rect 3390 4058 3394 4062
rect 3446 4058 3450 4062
rect 3414 3988 3418 3992
rect 3406 3968 3410 3972
rect 3422 3968 3426 3972
rect 3446 3968 3450 3972
rect 3358 3958 3362 3962
rect 3318 3948 3322 3952
rect 3334 3948 3338 3952
rect 3318 3928 3322 3932
rect 3254 3878 3258 3882
rect 3086 3738 3090 3742
rect 3118 3738 3122 3742
rect 3094 3698 3098 3702
rect 3102 3678 3106 3682
rect 3110 3668 3114 3672
rect 3078 3658 3082 3662
rect 3126 3728 3130 3732
rect 3222 3718 3226 3722
rect 3174 3688 3178 3692
rect 3206 3678 3210 3682
rect 3134 3668 3138 3672
rect 3190 3668 3194 3672
rect 3118 3658 3122 3662
rect 3150 3658 3154 3662
rect 3166 3658 3170 3662
rect 3086 3648 3090 3652
rect 3150 3648 3154 3652
rect 3054 3638 3058 3642
rect 3070 3638 3074 3642
rect 3118 3638 3122 3642
rect 3030 3588 3034 3592
rect 2990 3568 2994 3572
rect 3006 3568 3010 3572
rect 3006 3558 3010 3562
rect 2982 3548 2986 3552
rect 3014 3548 3018 3552
rect 3294 3848 3298 3852
rect 3278 3758 3282 3762
rect 3246 3748 3250 3752
rect 3262 3748 3266 3752
rect 3382 3948 3386 3952
rect 3374 3938 3378 3942
rect 3358 3928 3362 3932
rect 3406 3948 3410 3952
rect 3430 3938 3434 3942
rect 3438 3938 3442 3942
rect 3462 3978 3466 3982
rect 3502 4138 3506 4142
rect 3502 4118 3506 4122
rect 3510 4078 3514 4082
rect 3550 4108 3554 4112
rect 3558 4098 3562 4102
rect 3574 4128 3578 4132
rect 3582 4118 3586 4122
rect 3574 4098 3578 4102
rect 3566 4078 3570 4082
rect 3526 4068 3530 4072
rect 3502 4058 3506 4062
rect 3542 4048 3546 4052
rect 3510 3988 3514 3992
rect 3662 4258 3666 4262
rect 3654 4248 3658 4252
rect 3678 4248 3682 4252
rect 3678 4168 3682 4172
rect 3670 4148 3674 4152
rect 3678 4118 3682 4122
rect 3686 4108 3690 4112
rect 3662 4098 3666 4102
rect 3598 4088 3602 4092
rect 3630 4088 3634 4092
rect 3646 4088 3650 4092
rect 3566 4058 3570 4062
rect 3582 4058 3586 4062
rect 3614 4058 3618 4062
rect 3598 4048 3602 4052
rect 3646 4068 3650 4072
rect 3686 4088 3690 4092
rect 3678 4078 3682 4082
rect 3670 4058 3674 4062
rect 3646 4048 3650 4052
rect 3662 4048 3666 4052
rect 3574 4038 3578 4042
rect 3590 4038 3594 4042
rect 3630 4038 3634 4042
rect 3570 4003 3574 4007
rect 3577 4003 3581 4007
rect 3550 3978 3554 3982
rect 3566 3978 3570 3982
rect 3614 3978 3618 3982
rect 3590 3968 3594 3972
rect 3550 3958 3554 3962
rect 3470 3938 3474 3942
rect 3526 3928 3530 3932
rect 3550 3928 3554 3932
rect 3454 3918 3458 3922
rect 3518 3918 3522 3922
rect 3390 3898 3394 3902
rect 3430 3878 3434 3882
rect 3438 3878 3442 3882
rect 3382 3868 3386 3872
rect 3422 3868 3426 3872
rect 3494 3868 3498 3872
rect 3414 3858 3418 3862
rect 3462 3858 3466 3862
rect 3510 3858 3514 3862
rect 3350 3838 3354 3842
rect 3382 3818 3386 3822
rect 3414 3768 3418 3772
rect 3326 3758 3330 3762
rect 3398 3758 3402 3762
rect 3438 3758 3442 3762
rect 3518 3758 3522 3762
rect 3406 3748 3410 3752
rect 3454 3748 3458 3752
rect 3606 3958 3610 3962
rect 3582 3948 3586 3952
rect 3622 3958 3626 3962
rect 3622 3948 3626 3952
rect 3590 3938 3594 3942
rect 3654 3948 3658 3952
rect 3742 4268 3746 4272
rect 3710 4258 3714 4262
rect 3742 4258 3746 4262
rect 3710 4218 3714 4222
rect 3798 4338 3802 4342
rect 3758 4308 3762 4312
rect 3806 4328 3810 4332
rect 3838 4328 3842 4332
rect 3822 4318 3826 4322
rect 3902 4398 3906 4402
rect 3918 4398 3922 4402
rect 3942 4398 3946 4402
rect 3950 4398 3954 4402
rect 3966 4398 3970 4402
rect 3886 4348 3890 4352
rect 3894 4338 3898 4342
rect 3782 4298 3786 4302
rect 3830 4298 3834 4302
rect 3774 4288 3778 4292
rect 3878 4298 3882 4302
rect 3878 4288 3882 4292
rect 3886 4288 3890 4292
rect 3838 4278 3842 4282
rect 3758 4258 3762 4262
rect 3774 4258 3778 4262
rect 3750 4228 3754 4232
rect 3798 4258 3802 4262
rect 3822 4258 3826 4262
rect 3790 4248 3794 4252
rect 3822 4228 3826 4232
rect 3814 4208 3818 4212
rect 3758 4198 3762 4202
rect 3758 4158 3762 4162
rect 3766 4148 3770 4152
rect 3734 4138 3738 4142
rect 3758 4138 3762 4142
rect 3710 4128 3714 4132
rect 3734 4078 3738 4082
rect 3710 4038 3714 4042
rect 3750 4068 3754 4072
rect 3750 4048 3754 4052
rect 3702 4028 3706 4032
rect 3726 4028 3730 4032
rect 3766 4128 3770 4132
rect 3782 4098 3786 4102
rect 3814 4148 3818 4152
rect 3830 4158 3834 4162
rect 3814 4118 3818 4122
rect 3822 4108 3826 4112
rect 3798 4088 3802 4092
rect 3782 4078 3786 4082
rect 3814 4078 3818 4082
rect 3766 4068 3770 4072
rect 3798 4068 3802 4072
rect 3870 4258 3874 4262
rect 3846 4228 3850 4232
rect 3854 4208 3858 4212
rect 3934 4378 3938 4382
rect 3918 4368 3922 4372
rect 3926 4358 3930 4362
rect 3942 4368 3946 4372
rect 3942 4338 3946 4342
rect 3990 4398 3994 4402
rect 4006 4398 4010 4402
rect 4022 4398 4026 4402
rect 3982 4388 3986 4392
rect 3974 4368 3978 4372
rect 4062 4398 4066 4402
rect 4046 4388 4050 4392
rect 4022 4368 4026 4372
rect 4038 4368 4042 4372
rect 3966 4358 3970 4362
rect 3966 4348 3970 4352
rect 3998 4348 4002 4352
rect 4062 4348 4066 4352
rect 3966 4338 3970 4342
rect 3990 4338 3994 4342
rect 4006 4338 4010 4342
rect 3918 4298 3922 4302
rect 3918 4268 3922 4272
rect 3878 4208 3882 4212
rect 3878 4198 3882 4202
rect 3870 4178 3874 4182
rect 3870 4168 3874 4172
rect 3854 4138 3858 4142
rect 3846 4088 3850 4092
rect 3862 4118 3866 4122
rect 3870 4078 3874 4082
rect 3838 4058 3842 4062
rect 3910 4258 3914 4262
rect 3894 4228 3898 4232
rect 3886 4188 3890 4192
rect 3910 4168 3914 4172
rect 3958 4268 3962 4272
rect 3982 4328 3986 4332
rect 3974 4298 3978 4302
rect 4054 4328 4058 4332
rect 4086 4328 4090 4332
rect 4126 4398 4130 4402
rect 4118 4378 4122 4382
rect 4198 4378 4202 4382
rect 4318 4398 4322 4402
rect 4342 4398 4346 4402
rect 4230 4378 4234 4382
rect 4150 4358 4154 4362
rect 4222 4358 4226 4362
rect 4110 4348 4114 4352
rect 4142 4348 4146 4352
rect 4182 4348 4186 4352
rect 4222 4348 4226 4352
rect 4198 4338 4202 4342
rect 4126 4328 4130 4332
rect 4142 4328 4146 4332
rect 4046 4318 4050 4322
rect 4062 4318 4066 4322
rect 4078 4318 4082 4322
rect 4102 4318 4106 4322
rect 4166 4318 4170 4322
rect 4182 4318 4186 4322
rect 4054 4308 4058 4312
rect 4046 4298 4050 4302
rect 3998 4288 4002 4292
rect 4038 4288 4042 4292
rect 3998 4258 4002 4262
rect 4014 4258 4018 4262
rect 3966 4238 3970 4242
rect 3974 4228 3978 4232
rect 3942 4198 3946 4202
rect 3974 4198 3978 4202
rect 3974 4178 3978 4182
rect 3998 4178 4002 4182
rect 3950 4168 3954 4172
rect 3966 4158 3970 4162
rect 4022 4248 4026 4252
rect 4014 4208 4018 4212
rect 4006 4148 4010 4152
rect 3918 4138 3922 4142
rect 3950 4138 3954 4142
rect 3894 4128 3898 4132
rect 3926 4128 3930 4132
rect 3918 4108 3922 4112
rect 3926 4108 3930 4112
rect 3918 4078 3922 4082
rect 3886 4068 3890 4072
rect 3894 4058 3898 4062
rect 3934 4058 3938 4062
rect 3774 4048 3778 4052
rect 3790 4048 3794 4052
rect 3806 4048 3810 4052
rect 3870 4048 3874 4052
rect 3734 4018 3738 4022
rect 3694 3978 3698 3982
rect 3750 3988 3754 3992
rect 3726 3958 3730 3962
rect 3686 3938 3690 3942
rect 3662 3928 3666 3932
rect 3630 3918 3634 3922
rect 3646 3918 3650 3922
rect 3582 3908 3586 3912
rect 3582 3898 3586 3902
rect 3566 3878 3570 3882
rect 3566 3868 3570 3872
rect 3590 3858 3594 3862
rect 3590 3848 3594 3852
rect 3558 3828 3562 3832
rect 3606 3818 3610 3822
rect 3570 3803 3574 3807
rect 3577 3803 3581 3807
rect 3606 3778 3610 3782
rect 3270 3738 3274 3742
rect 3406 3738 3410 3742
rect 3430 3738 3434 3742
rect 3462 3738 3466 3742
rect 3254 3728 3258 3732
rect 3358 3728 3362 3732
rect 3438 3718 3442 3722
rect 3262 3708 3266 3712
rect 3390 3708 3394 3712
rect 3238 3698 3242 3702
rect 3214 3668 3218 3672
rect 3230 3668 3234 3672
rect 3222 3658 3226 3662
rect 3182 3638 3186 3642
rect 3214 3638 3218 3642
rect 3078 3628 3082 3632
rect 3174 3628 3178 3632
rect 3430 3678 3434 3682
rect 3310 3658 3314 3662
rect 3342 3658 3346 3662
rect 3294 3648 3298 3652
rect 3366 3638 3370 3642
rect 3254 3628 3258 3632
rect 3222 3618 3226 3622
rect 3102 3588 3106 3592
rect 3110 3578 3114 3582
rect 3078 3558 3082 3562
rect 3046 3528 3050 3532
rect 3054 3528 3058 3532
rect 3062 3518 3066 3522
rect 3050 3503 3054 3507
rect 3057 3503 3061 3507
rect 3014 3498 3018 3502
rect 3110 3548 3114 3552
rect 3126 3548 3130 3552
rect 3086 3528 3090 3532
rect 3094 3518 3098 3522
rect 3006 3468 3010 3472
rect 3038 3468 3042 3472
rect 3102 3468 3106 3472
rect 2990 3458 2994 3462
rect 3030 3458 3034 3462
rect 2998 3448 3002 3452
rect 2958 3438 2962 3442
rect 2974 3438 2978 3442
rect 2886 3428 2890 3432
rect 2934 3428 2938 3432
rect 2966 3428 2970 3432
rect 3022 3438 3026 3442
rect 3014 3428 3018 3432
rect 2862 3418 2866 3422
rect 2990 3418 2994 3422
rect 2886 3398 2890 3402
rect 2846 3388 2850 3392
rect 2846 3378 2850 3382
rect 2830 3368 2834 3372
rect 2926 3378 2930 3382
rect 2910 3368 2914 3372
rect 2974 3408 2978 3412
rect 2998 3378 3002 3382
rect 2958 3358 2962 3362
rect 2998 3358 3002 3362
rect 2806 3348 2810 3352
rect 2822 3348 2826 3352
rect 2846 3348 2850 3352
rect 2902 3348 2906 3352
rect 2998 3348 3002 3352
rect 2686 3338 2690 3342
rect 2574 3258 2578 3262
rect 2510 3248 2514 3252
rect 2542 3248 2546 3252
rect 2630 3308 2634 3312
rect 2694 3328 2698 3332
rect 2790 3338 2794 3342
rect 2854 3338 2858 3342
rect 2918 3338 2922 3342
rect 2966 3338 2970 3342
rect 2710 3308 2714 3312
rect 2782 3318 2786 3322
rect 2838 3318 2842 3322
rect 2846 3308 2850 3312
rect 2870 3328 2874 3332
rect 2878 3318 2882 3322
rect 2886 3308 2890 3312
rect 2894 3308 2898 3312
rect 2910 3328 2914 3332
rect 2902 3298 2906 3302
rect 2934 3308 2938 3312
rect 2926 3298 2930 3302
rect 2958 3328 2962 3332
rect 2998 3318 3002 3322
rect 3022 3328 3026 3332
rect 3030 3318 3034 3322
rect 3086 3458 3090 3462
rect 3094 3458 3098 3462
rect 3270 3618 3274 3622
rect 3278 3618 3282 3622
rect 3246 3608 3250 3612
rect 3238 3598 3242 3602
rect 3190 3578 3194 3582
rect 3150 3568 3154 3572
rect 3230 3568 3234 3572
rect 3150 3538 3154 3542
rect 3182 3538 3186 3542
rect 3150 3498 3154 3502
rect 3142 3468 3146 3472
rect 3126 3458 3130 3462
rect 3158 3458 3162 3462
rect 3222 3518 3226 3522
rect 3222 3488 3226 3492
rect 3214 3468 3218 3472
rect 3118 3448 3122 3452
rect 3150 3448 3154 3452
rect 3174 3448 3178 3452
rect 3198 3448 3202 3452
rect 3222 3448 3226 3452
rect 3254 3518 3258 3522
rect 3254 3468 3258 3472
rect 3326 3588 3330 3592
rect 3286 3568 3290 3572
rect 3310 3568 3314 3572
rect 3278 3538 3282 3542
rect 3318 3518 3322 3522
rect 3294 3498 3298 3502
rect 3286 3468 3290 3472
rect 3278 3458 3282 3462
rect 3278 3448 3282 3452
rect 3318 3468 3322 3472
rect 3334 3578 3338 3582
rect 3334 3568 3338 3572
rect 3374 3558 3378 3562
rect 3342 3538 3346 3542
rect 3358 3528 3362 3532
rect 3342 3518 3346 3522
rect 3446 3668 3450 3672
rect 3534 3728 3538 3732
rect 3494 3698 3498 3702
rect 3414 3658 3418 3662
rect 3542 3658 3546 3662
rect 3406 3648 3410 3652
rect 3406 3578 3410 3582
rect 3390 3568 3394 3572
rect 3398 3558 3402 3562
rect 3438 3648 3442 3652
rect 3438 3608 3442 3612
rect 3422 3558 3426 3562
rect 3398 3538 3402 3542
rect 3414 3538 3418 3542
rect 3358 3468 3362 3472
rect 3390 3468 3394 3472
rect 3414 3468 3418 3472
rect 3430 3468 3434 3472
rect 3342 3458 3346 3462
rect 3374 3458 3378 3462
rect 3326 3448 3330 3452
rect 3150 3438 3154 3442
rect 3198 3438 3202 3442
rect 3310 3438 3314 3442
rect 3350 3438 3354 3442
rect 3230 3428 3234 3432
rect 3070 3358 3074 3362
rect 3054 3318 3058 3322
rect 3062 3318 3066 3322
rect 3050 3303 3054 3307
rect 3057 3303 3061 3307
rect 2974 3288 2978 3292
rect 2630 3278 2634 3282
rect 2934 3278 2938 3282
rect 2614 3268 2618 3272
rect 2638 3268 2642 3272
rect 2662 3268 2666 3272
rect 2718 3268 2722 3272
rect 2910 3268 2914 3272
rect 2606 3258 2610 3262
rect 2590 3238 2594 3242
rect 2398 3208 2402 3212
rect 2494 3208 2498 3212
rect 2574 3208 2578 3212
rect 2546 3203 2550 3207
rect 2553 3203 2557 3207
rect 2358 3198 2362 3202
rect 2366 3198 2370 3202
rect 2438 3168 2442 3172
rect 2462 3168 2466 3172
rect 2486 3168 2490 3172
rect 2510 3168 2514 3172
rect 2398 3158 2402 3162
rect 2542 3158 2546 3162
rect 2294 3148 2298 3152
rect 2318 3148 2322 3152
rect 2334 3148 2338 3152
rect 2302 3138 2306 3142
rect 2278 3108 2282 3112
rect 2294 3098 2298 3102
rect 2318 3098 2322 3102
rect 2294 3088 2298 3092
rect 2318 3088 2322 3092
rect 2310 3068 2314 3072
rect 2294 3058 2298 3062
rect 2286 3048 2290 3052
rect 2294 3038 2298 3042
rect 2318 3028 2322 3032
rect 2310 2998 2314 3002
rect 2358 3148 2362 3152
rect 2382 3148 2386 3152
rect 2342 3128 2346 3132
rect 2342 3108 2346 3112
rect 2398 3118 2402 3122
rect 2382 3098 2386 3102
rect 2374 3088 2378 3092
rect 2358 3058 2362 3062
rect 2358 3048 2362 3052
rect 2334 2978 2338 2982
rect 2310 2968 2314 2972
rect 2158 2938 2162 2942
rect 2198 2938 2202 2942
rect 2270 2938 2274 2942
rect 2286 2938 2290 2942
rect 2030 2928 2034 2932
rect 2118 2928 2122 2932
rect 1910 2918 1914 2922
rect 1942 2898 1946 2902
rect 2046 2908 2050 2912
rect 2026 2903 2030 2907
rect 2033 2903 2037 2907
rect 1950 2868 1954 2872
rect 1910 2848 1914 2852
rect 1902 2778 1906 2782
rect 2022 2858 2026 2862
rect 2006 2828 2010 2832
rect 2006 2808 2010 2812
rect 1974 2778 1978 2782
rect 1910 2768 1914 2772
rect 1862 2758 1866 2762
rect 1814 2748 1818 2752
rect 1886 2748 1890 2752
rect 1822 2738 1826 2742
rect 1742 2728 1746 2732
rect 1742 2718 1746 2722
rect 1790 2718 1794 2722
rect 1758 2708 1762 2712
rect 1702 2678 1706 2682
rect 1798 2678 1802 2682
rect 1766 2668 1770 2672
rect 1702 2658 1706 2662
rect 1734 2658 1738 2662
rect 1782 2598 1786 2602
rect 1798 2588 1802 2592
rect 1734 2568 1738 2572
rect 1734 2548 1738 2552
rect 1726 2538 1730 2542
rect 1670 2498 1674 2502
rect 1678 2468 1682 2472
rect 1686 2448 1690 2452
rect 1662 2418 1666 2422
rect 1662 2398 1666 2402
rect 1654 2358 1658 2362
rect 1702 2358 1706 2362
rect 1574 2298 1578 2302
rect 1590 2298 1594 2302
rect 1550 2278 1554 2282
rect 1574 2268 1578 2272
rect 1478 2228 1482 2232
rect 1422 2218 1426 2222
rect 1470 2218 1474 2222
rect 1286 2178 1290 2182
rect 1310 2178 1314 2182
rect 1318 2168 1322 2172
rect 1422 2168 1426 2172
rect 1294 2078 1298 2082
rect 1246 2058 1250 2062
rect 1262 2058 1266 2062
rect 1414 2158 1418 2162
rect 1430 2158 1434 2162
rect 1438 2158 1442 2162
rect 1470 2158 1474 2162
rect 1334 2138 1338 2142
rect 1522 2203 1526 2207
rect 1529 2203 1533 2207
rect 1502 2158 1506 2162
rect 1446 2138 1450 2142
rect 1454 2138 1458 2142
rect 1398 2128 1402 2132
rect 1462 2128 1466 2132
rect 1494 2128 1498 2132
rect 1326 2058 1330 2062
rect 1278 2048 1282 2052
rect 1302 2048 1306 2052
rect 1158 2038 1162 2042
rect 1310 2038 1314 2042
rect 1326 2038 1330 2042
rect 1118 1968 1122 1972
rect 814 1948 818 1952
rect 1046 1948 1050 1952
rect 1126 1948 1130 1952
rect 1134 1948 1138 1952
rect 758 1938 762 1942
rect 910 1938 914 1942
rect 830 1928 834 1932
rect 974 1928 978 1932
rect 734 1918 738 1922
rect 782 1908 786 1912
rect 686 1888 690 1892
rect 726 1888 730 1892
rect 734 1888 738 1892
rect 766 1888 770 1892
rect 710 1868 714 1872
rect 606 1858 610 1862
rect 630 1858 634 1862
rect 662 1858 666 1862
rect 558 1828 562 1832
rect 498 1803 502 1807
rect 505 1803 509 1807
rect 582 1798 586 1802
rect 550 1768 554 1772
rect 486 1758 490 1762
rect 606 1848 610 1852
rect 622 1848 626 1852
rect 638 1848 642 1852
rect 678 1818 682 1822
rect 590 1768 594 1772
rect 638 1758 642 1762
rect 438 1668 442 1672
rect 366 1638 370 1642
rect 390 1628 394 1632
rect 398 1608 402 1612
rect 398 1588 402 1592
rect 350 1578 354 1582
rect 374 1578 378 1582
rect 374 1568 378 1572
rect 382 1558 386 1562
rect 390 1548 394 1552
rect 374 1538 378 1542
rect 398 1538 402 1542
rect 342 1528 346 1532
rect 366 1528 370 1532
rect 382 1518 386 1522
rect 334 1508 338 1512
rect 366 1508 370 1512
rect 350 1498 354 1502
rect 334 1488 338 1492
rect 350 1488 354 1492
rect 390 1488 394 1492
rect 326 1478 330 1482
rect 278 1458 282 1462
rect 286 1448 290 1452
rect 262 1438 266 1442
rect 294 1438 298 1442
rect 222 1428 226 1432
rect 262 1408 266 1412
rect 278 1358 282 1362
rect 230 1348 234 1352
rect 214 1318 218 1322
rect 246 1318 250 1322
rect 190 1278 194 1282
rect 206 1278 210 1282
rect 230 1278 234 1282
rect 158 1268 162 1272
rect 182 1268 186 1272
rect 6 1248 10 1252
rect 30 1178 34 1182
rect 54 1178 58 1182
rect 70 1178 74 1182
rect 46 1158 50 1162
rect 78 1158 82 1162
rect 166 1258 170 1262
rect 190 1258 194 1262
rect 214 1258 218 1262
rect 230 1258 234 1262
rect 318 1368 322 1372
rect 422 1648 426 1652
rect 414 1578 418 1582
rect 422 1558 426 1562
rect 438 1558 442 1562
rect 462 1558 466 1562
rect 438 1538 442 1542
rect 454 1538 458 1542
rect 422 1528 426 1532
rect 454 1528 458 1532
rect 470 1518 474 1522
rect 598 1748 602 1752
rect 742 1878 746 1882
rect 766 1878 770 1882
rect 758 1778 762 1782
rect 734 1768 738 1772
rect 718 1758 722 1762
rect 710 1748 714 1752
rect 726 1748 730 1752
rect 494 1659 498 1663
rect 534 1658 538 1662
rect 670 1728 674 1732
rect 670 1718 674 1722
rect 606 1668 610 1672
rect 902 1898 906 1902
rect 934 1898 938 1902
rect 822 1878 826 1882
rect 806 1868 810 1872
rect 838 1868 842 1872
rect 870 1868 874 1872
rect 1002 1903 1006 1907
rect 1009 1903 1013 1907
rect 1070 1938 1074 1942
rect 1078 1928 1082 1932
rect 1054 1918 1058 1922
rect 1382 2098 1386 2102
rect 1406 2098 1410 2102
rect 1358 2088 1362 2092
rect 1406 2088 1410 2092
rect 1438 2108 1442 2112
rect 1422 2078 1426 2082
rect 1350 2068 1354 2072
rect 1366 2068 1370 2072
rect 1382 2068 1386 2072
rect 1406 2068 1410 2072
rect 1518 2098 1522 2102
rect 1462 2088 1466 2092
rect 1510 2088 1514 2092
rect 1342 2048 1346 2052
rect 1374 2048 1378 2052
rect 1390 2048 1394 2052
rect 1398 2038 1402 2042
rect 1334 2018 1338 2022
rect 1366 2018 1370 2022
rect 1190 1998 1194 2002
rect 1222 1998 1226 2002
rect 1174 1968 1178 1972
rect 1166 1948 1170 1952
rect 1134 1938 1138 1942
rect 1134 1928 1138 1932
rect 1150 1928 1154 1932
rect 1094 1908 1098 1912
rect 1158 1908 1162 1912
rect 1022 1888 1026 1892
rect 1030 1878 1034 1882
rect 958 1868 962 1872
rect 918 1858 922 1862
rect 790 1848 794 1852
rect 838 1848 842 1852
rect 790 1838 794 1842
rect 910 1838 914 1842
rect 862 1818 866 1822
rect 838 1768 842 1772
rect 894 1758 898 1762
rect 830 1748 834 1752
rect 846 1748 850 1752
rect 766 1728 770 1732
rect 742 1688 746 1692
rect 806 1738 810 1742
rect 798 1698 802 1702
rect 694 1658 698 1662
rect 718 1658 722 1662
rect 566 1638 570 1642
rect 686 1638 690 1642
rect 702 1638 706 1642
rect 498 1603 502 1607
rect 505 1603 509 1607
rect 734 1658 738 1662
rect 750 1658 754 1662
rect 1110 1898 1114 1902
rect 1118 1888 1122 1892
rect 1118 1868 1122 1872
rect 1094 1828 1098 1832
rect 990 1818 994 1822
rect 1046 1818 1050 1822
rect 958 1808 962 1812
rect 1022 1768 1026 1772
rect 1054 1768 1058 1772
rect 998 1748 1002 1752
rect 1006 1748 1010 1752
rect 1046 1758 1050 1762
rect 1030 1748 1034 1752
rect 1158 1798 1162 1802
rect 1094 1758 1098 1762
rect 1126 1758 1130 1762
rect 1134 1758 1138 1762
rect 1086 1748 1090 1752
rect 1078 1738 1082 1742
rect 1094 1738 1098 1742
rect 1110 1738 1114 1742
rect 974 1728 978 1732
rect 1118 1728 1122 1732
rect 862 1688 866 1692
rect 1002 1703 1006 1707
rect 1009 1703 1013 1707
rect 1014 1688 1018 1692
rect 1206 1948 1210 1952
rect 1230 1948 1234 1952
rect 1262 1948 1266 1952
rect 1430 1998 1434 2002
rect 1334 1958 1338 1962
rect 1366 1958 1370 1962
rect 1470 2068 1474 2072
rect 1550 2068 1554 2072
rect 1534 2058 1538 2062
rect 1502 2028 1506 2032
rect 1522 2003 1526 2007
rect 1529 2003 1533 2007
rect 1518 1958 1522 1962
rect 1454 1948 1458 1952
rect 1486 1948 1490 1952
rect 1510 1948 1514 1952
rect 1214 1938 1218 1942
rect 1238 1938 1242 1942
rect 1254 1938 1258 1942
rect 1270 1938 1274 1942
rect 1286 1938 1290 1942
rect 1294 1938 1298 1942
rect 1262 1928 1266 1932
rect 1286 1928 1290 1932
rect 1406 1928 1410 1932
rect 1198 1918 1202 1922
rect 1222 1918 1226 1922
rect 1182 1878 1186 1882
rect 1174 1848 1178 1852
rect 1166 1768 1170 1772
rect 1142 1708 1146 1712
rect 1158 1708 1162 1712
rect 1134 1698 1138 1702
rect 1182 1838 1186 1842
rect 1206 1908 1210 1912
rect 1254 1908 1258 1912
rect 1334 1918 1338 1922
rect 1278 1868 1282 1872
rect 1198 1858 1202 1862
rect 1230 1858 1234 1862
rect 1246 1848 1250 1852
rect 1222 1828 1226 1832
rect 1198 1798 1202 1802
rect 1190 1788 1194 1792
rect 1262 1858 1266 1862
rect 1278 1858 1282 1862
rect 1254 1768 1258 1772
rect 1182 1758 1186 1762
rect 1294 1848 1298 1852
rect 1278 1768 1282 1772
rect 1270 1758 1274 1762
rect 1310 1878 1314 1882
rect 1326 1868 1330 1872
rect 1382 1888 1386 1892
rect 1406 1888 1410 1892
rect 1350 1878 1354 1882
rect 1366 1878 1370 1882
rect 1374 1868 1378 1872
rect 1502 1938 1506 1942
rect 1534 1938 1538 1942
rect 1742 2508 1746 2512
rect 1830 2718 1834 2722
rect 1830 2668 1834 2672
rect 1862 2718 1866 2722
rect 1894 2718 1898 2722
rect 1894 2678 1898 2682
rect 1846 2598 1850 2602
rect 1926 2758 1930 2762
rect 1990 2748 1994 2752
rect 1974 2688 1978 2692
rect 1990 2678 1994 2682
rect 2054 2898 2058 2902
rect 2086 2868 2090 2872
rect 2150 2878 2154 2882
rect 2182 2868 2186 2872
rect 2134 2858 2138 2862
rect 2046 2778 2050 2782
rect 2086 2778 2090 2782
rect 2174 2798 2178 2802
rect 2150 2747 2154 2751
rect 2022 2738 2026 2742
rect 2014 2728 2018 2732
rect 2086 2728 2090 2732
rect 1966 2558 1970 2562
rect 1886 2548 1890 2552
rect 1910 2548 1914 2552
rect 1950 2548 1954 2552
rect 1982 2548 1986 2552
rect 1830 2538 1834 2542
rect 1942 2538 1946 2542
rect 1838 2528 1842 2532
rect 1854 2528 1858 2532
rect 1758 2478 1762 2482
rect 1806 2478 1810 2482
rect 1774 2468 1778 2472
rect 1870 2468 1874 2472
rect 1798 2459 1802 2463
rect 1798 2418 1802 2422
rect 2158 2718 2162 2722
rect 2026 2703 2030 2707
rect 2033 2703 2037 2707
rect 2054 2698 2058 2702
rect 2030 2688 2034 2692
rect 2110 2688 2114 2692
rect 2102 2678 2106 2682
rect 2086 2618 2090 2622
rect 2110 2608 2114 2612
rect 2142 2588 2146 2592
rect 2054 2558 2058 2562
rect 2086 2558 2090 2562
rect 1966 2538 1970 2542
rect 1990 2538 1994 2542
rect 1998 2538 2002 2542
rect 2126 2538 2130 2542
rect 2142 2538 2146 2542
rect 1902 2448 1906 2452
rect 1798 2368 1802 2372
rect 1894 2368 1898 2372
rect 1950 2368 1954 2372
rect 1646 2338 1650 2342
rect 1694 2338 1698 2342
rect 1790 2338 1794 2342
rect 1750 2318 1754 2322
rect 1670 2278 1674 2282
rect 1606 2258 1610 2262
rect 1918 2358 1922 2362
rect 1822 2298 1826 2302
rect 1846 2298 1850 2302
rect 1886 2288 1890 2292
rect 1886 2278 1890 2282
rect 1918 2268 1922 2272
rect 1854 2178 1858 2182
rect 1686 2168 1690 2172
rect 1774 2168 1778 2172
rect 1726 2158 1730 2162
rect 1854 2158 1858 2162
rect 1694 2148 1698 2152
rect 1742 2148 1746 2152
rect 1774 2148 1778 2152
rect 1950 2328 1954 2332
rect 2026 2503 2030 2507
rect 2033 2503 2037 2507
rect 2094 2498 2098 2502
rect 2022 2488 2026 2492
rect 2038 2488 2042 2492
rect 2046 2488 2050 2492
rect 2078 2468 2082 2472
rect 1974 2358 1978 2362
rect 1670 2138 1674 2142
rect 1686 2138 1690 2142
rect 1702 2138 1706 2142
rect 1654 2088 1658 2092
rect 1678 2128 1682 2132
rect 1574 2078 1578 2082
rect 1606 2078 1610 2082
rect 1622 2078 1626 2082
rect 1670 2078 1674 2082
rect 1566 2058 1570 2062
rect 1590 2058 1594 2062
rect 1574 2028 1578 2032
rect 1726 2138 1730 2142
rect 1718 2128 1722 2132
rect 1710 2118 1714 2122
rect 1782 2138 1786 2142
rect 1758 2128 1762 2132
rect 1750 2108 1754 2112
rect 1710 2098 1714 2102
rect 1742 2098 1746 2102
rect 1702 2068 1706 2072
rect 1638 2058 1642 2062
rect 1630 2028 1634 2032
rect 1686 2058 1690 2062
rect 1766 2088 1770 2092
rect 1734 2078 1738 2082
rect 1670 2048 1674 2052
rect 1710 2038 1714 2042
rect 1646 2018 1650 2022
rect 1662 2018 1666 2022
rect 1702 2018 1706 2022
rect 1718 2018 1722 2022
rect 1646 1978 1650 1982
rect 1598 1968 1602 1972
rect 1678 1968 1682 1972
rect 1614 1958 1618 1962
rect 1638 1958 1642 1962
rect 1622 1948 1626 1952
rect 1654 1948 1658 1952
rect 1558 1938 1562 1942
rect 1566 1938 1570 1942
rect 1638 1938 1642 1942
rect 1662 1938 1666 1942
rect 1550 1928 1554 1932
rect 1590 1928 1594 1932
rect 1614 1928 1618 1932
rect 1470 1918 1474 1922
rect 1494 1918 1498 1922
rect 1566 1918 1570 1922
rect 1630 1918 1634 1922
rect 1422 1878 1426 1882
rect 1350 1858 1354 1862
rect 1414 1848 1418 1852
rect 1454 1848 1458 1852
rect 1342 1838 1346 1842
rect 1246 1748 1250 1752
rect 1254 1748 1258 1752
rect 1278 1748 1282 1752
rect 1302 1748 1306 1752
rect 1326 1748 1330 1752
rect 1182 1728 1186 1732
rect 1198 1728 1202 1732
rect 1254 1728 1258 1732
rect 1222 1708 1226 1712
rect 1374 1788 1378 1792
rect 1366 1768 1370 1772
rect 1310 1738 1314 1742
rect 1342 1738 1346 1742
rect 1342 1728 1346 1732
rect 1358 1728 1362 1732
rect 1174 1688 1178 1692
rect 1222 1688 1226 1692
rect 1286 1688 1290 1692
rect 1310 1688 1314 1692
rect 1326 1688 1330 1692
rect 974 1678 978 1682
rect 1054 1678 1058 1682
rect 1126 1678 1130 1682
rect 1206 1678 1210 1682
rect 1246 1678 1250 1682
rect 1310 1678 1314 1682
rect 926 1668 930 1672
rect 966 1668 970 1672
rect 1158 1668 1162 1672
rect 1174 1668 1178 1672
rect 1254 1668 1258 1672
rect 726 1638 730 1642
rect 726 1618 730 1622
rect 510 1578 514 1582
rect 598 1578 602 1582
rect 622 1578 626 1582
rect 534 1568 538 1572
rect 502 1548 506 1552
rect 630 1558 634 1562
rect 542 1548 546 1552
rect 558 1548 562 1552
rect 566 1538 570 1542
rect 558 1518 562 1522
rect 486 1508 490 1512
rect 406 1478 410 1482
rect 414 1478 418 1482
rect 430 1478 434 1482
rect 406 1468 410 1472
rect 350 1458 354 1462
rect 358 1448 362 1452
rect 390 1378 394 1382
rect 390 1368 394 1372
rect 310 1348 314 1352
rect 326 1328 330 1332
rect 294 1318 298 1322
rect 302 1308 306 1312
rect 270 1278 274 1282
rect 278 1278 282 1282
rect 318 1278 322 1282
rect 254 1268 258 1272
rect 334 1268 338 1272
rect 286 1258 290 1262
rect 302 1258 306 1262
rect 326 1258 330 1262
rect 270 1248 274 1252
rect 342 1248 346 1252
rect 238 1228 242 1232
rect 118 1188 122 1192
rect 166 1178 170 1182
rect 142 1158 146 1162
rect 6 1148 10 1152
rect 22 1118 26 1122
rect 30 1078 34 1082
rect 46 1068 50 1072
rect 158 1148 162 1152
rect 206 1138 210 1142
rect 230 1138 234 1142
rect 134 1118 138 1122
rect 118 1088 122 1092
rect 30 1058 34 1062
rect 54 1058 58 1062
rect 6 1048 10 1052
rect 94 988 98 992
rect 6 948 10 952
rect 334 1218 338 1222
rect 342 1198 346 1202
rect 334 1188 338 1192
rect 286 1178 290 1182
rect 326 1168 330 1172
rect 302 1158 306 1162
rect 318 1128 322 1132
rect 302 1108 306 1112
rect 294 1098 298 1102
rect 270 1078 274 1082
rect 150 1068 154 1072
rect 270 1068 274 1072
rect 158 1058 162 1062
rect 246 1048 250 1052
rect 214 1008 218 1012
rect 206 998 210 1002
rect 246 968 250 972
rect 142 958 146 962
rect 198 948 202 952
rect 214 948 218 952
rect 222 938 226 942
rect 22 928 26 932
rect 126 928 130 932
rect 182 928 186 932
rect 6 878 10 882
rect 30 848 34 852
rect 134 858 138 862
rect 150 858 154 862
rect 118 818 122 822
rect 70 798 74 802
rect 134 768 138 772
rect 142 758 146 762
rect 182 878 186 882
rect 222 878 226 882
rect 246 878 250 882
rect 206 868 210 872
rect 310 1068 314 1072
rect 270 1058 274 1062
rect 310 1058 314 1062
rect 382 1348 386 1352
rect 358 1318 362 1322
rect 366 1308 370 1312
rect 446 1438 450 1442
rect 462 1428 466 1432
rect 438 1398 442 1402
rect 462 1388 466 1392
rect 438 1358 442 1362
rect 582 1548 586 1552
rect 614 1548 618 1552
rect 590 1538 594 1542
rect 574 1528 578 1532
rect 582 1528 586 1532
rect 566 1498 570 1502
rect 550 1478 554 1482
rect 606 1458 610 1462
rect 622 1468 626 1472
rect 534 1448 538 1452
rect 566 1448 570 1452
rect 598 1448 602 1452
rect 558 1438 562 1442
rect 566 1438 570 1442
rect 478 1418 482 1422
rect 498 1403 502 1407
rect 505 1403 509 1407
rect 478 1358 482 1362
rect 574 1348 578 1352
rect 470 1338 474 1342
rect 494 1338 498 1342
rect 542 1338 546 1342
rect 438 1318 442 1322
rect 358 1278 362 1282
rect 422 1278 426 1282
rect 366 1268 370 1272
rect 374 1268 378 1272
rect 414 1258 418 1262
rect 558 1328 562 1332
rect 550 1288 554 1292
rect 478 1278 482 1282
rect 470 1268 474 1272
rect 582 1318 586 1322
rect 614 1438 618 1442
rect 606 1378 610 1382
rect 598 1338 602 1342
rect 590 1288 594 1292
rect 590 1278 594 1282
rect 558 1268 562 1272
rect 606 1328 610 1332
rect 670 1538 674 1542
rect 718 1528 722 1532
rect 718 1518 722 1522
rect 662 1428 666 1432
rect 854 1658 858 1662
rect 878 1658 882 1662
rect 766 1648 770 1652
rect 838 1638 842 1642
rect 870 1638 874 1642
rect 774 1608 778 1612
rect 758 1598 762 1602
rect 742 1578 746 1582
rect 870 1608 874 1612
rect 894 1608 898 1612
rect 838 1598 842 1602
rect 910 1598 914 1602
rect 830 1588 834 1592
rect 958 1588 962 1592
rect 782 1578 786 1582
rect 1286 1668 1290 1672
rect 1318 1668 1322 1672
rect 982 1608 986 1612
rect 1062 1598 1066 1602
rect 982 1578 986 1582
rect 878 1568 882 1572
rect 918 1568 922 1572
rect 926 1568 930 1572
rect 790 1558 794 1562
rect 822 1558 826 1562
rect 766 1548 770 1552
rect 806 1528 810 1532
rect 902 1528 906 1532
rect 878 1488 882 1492
rect 918 1488 922 1492
rect 758 1478 762 1482
rect 814 1468 818 1472
rect 862 1468 866 1472
rect 806 1458 810 1462
rect 718 1378 722 1382
rect 678 1358 682 1362
rect 710 1358 714 1362
rect 694 1328 698 1332
rect 614 1308 618 1312
rect 654 1308 658 1312
rect 622 1298 626 1302
rect 782 1368 786 1372
rect 774 1358 778 1362
rect 782 1358 786 1362
rect 758 1348 762 1352
rect 734 1288 738 1292
rect 702 1258 706 1262
rect 718 1258 722 1262
rect 446 1248 450 1252
rect 542 1248 546 1252
rect 510 1228 514 1232
rect 498 1203 502 1207
rect 505 1203 509 1207
rect 446 1198 450 1202
rect 350 1168 354 1172
rect 406 1168 410 1172
rect 406 1158 410 1162
rect 598 1248 602 1252
rect 582 1238 586 1242
rect 574 1208 578 1212
rect 566 1188 570 1192
rect 454 1168 458 1172
rect 478 1168 482 1172
rect 606 1238 610 1242
rect 678 1228 682 1232
rect 654 1168 658 1172
rect 470 1158 474 1162
rect 566 1158 570 1162
rect 582 1158 586 1162
rect 614 1158 618 1162
rect 638 1158 642 1162
rect 438 1148 442 1152
rect 470 1148 474 1152
rect 558 1148 562 1152
rect 398 1138 402 1142
rect 446 1138 450 1142
rect 350 1118 354 1122
rect 398 1118 402 1122
rect 414 1108 418 1112
rect 542 1138 546 1142
rect 574 1138 578 1142
rect 486 1118 490 1122
rect 478 1098 482 1102
rect 454 1078 458 1082
rect 414 1068 418 1072
rect 438 1068 442 1072
rect 350 1058 354 1062
rect 342 1038 346 1042
rect 358 1018 362 1022
rect 278 998 282 1002
rect 326 998 330 1002
rect 310 968 314 972
rect 278 958 282 962
rect 262 948 266 952
rect 286 948 290 952
rect 310 948 314 952
rect 358 948 362 952
rect 326 938 330 942
rect 438 1058 442 1062
rect 382 1028 386 1032
rect 390 1028 394 1032
rect 390 1018 394 1022
rect 374 1008 378 1012
rect 390 988 394 992
rect 406 978 410 982
rect 422 978 426 982
rect 398 958 402 962
rect 390 948 394 952
rect 270 928 274 932
rect 286 928 290 932
rect 366 928 370 932
rect 382 928 386 932
rect 270 898 274 902
rect 222 828 226 832
rect 230 788 234 792
rect 142 748 146 752
rect 174 748 178 752
rect 150 738 154 742
rect 182 738 186 742
rect 206 738 210 742
rect 222 738 226 742
rect 286 858 290 862
rect 374 858 378 862
rect 358 848 362 852
rect 374 838 378 842
rect 334 828 338 832
rect 318 798 322 802
rect 302 788 306 792
rect 302 778 306 782
rect 318 768 322 772
rect 286 758 290 762
rect 142 728 146 732
rect 166 728 170 732
rect 198 728 202 732
rect 6 688 10 692
rect 22 688 26 692
rect 102 718 106 722
rect 134 718 138 722
rect 126 688 130 692
rect 86 659 90 663
rect 6 648 10 652
rect 30 648 34 652
rect 30 578 34 582
rect 182 718 186 722
rect 174 708 178 712
rect 150 698 154 702
rect 142 658 146 662
rect 134 648 138 652
rect 158 648 162 652
rect 182 688 186 692
rect 230 718 234 722
rect 214 698 218 702
rect 206 678 210 682
rect 222 688 226 692
rect 246 668 250 672
rect 182 658 186 662
rect 238 658 242 662
rect 190 648 194 652
rect 166 618 170 622
rect 142 578 146 582
rect 174 578 178 582
rect 6 548 10 552
rect 110 548 114 552
rect 246 648 250 652
rect 262 738 266 742
rect 318 738 322 742
rect 302 728 306 732
rect 366 748 370 752
rect 358 738 362 742
rect 342 708 346 712
rect 294 688 298 692
rect 270 678 274 682
rect 286 648 290 652
rect 254 638 258 642
rect 262 638 266 642
rect 254 618 258 622
rect 278 618 282 622
rect 254 558 258 562
rect 278 548 282 552
rect 206 538 210 542
rect 198 498 202 502
rect 22 458 26 462
rect 6 448 10 452
rect 86 458 90 462
rect 54 448 58 452
rect 78 368 82 372
rect 22 358 26 362
rect 46 358 50 362
rect 38 348 42 352
rect 70 348 74 352
rect 22 328 26 332
rect 6 318 10 322
rect 30 318 34 322
rect 54 318 58 322
rect 6 248 10 252
rect 22 188 26 192
rect 222 468 226 472
rect 166 458 170 462
rect 310 658 314 662
rect 326 648 330 652
rect 326 558 330 562
rect 310 548 314 552
rect 270 498 274 502
rect 262 488 266 492
rect 254 458 258 462
rect 126 448 130 452
rect 190 448 194 452
rect 230 448 234 452
rect 238 448 242 452
rect 126 438 130 442
rect 238 428 242 432
rect 246 388 250 392
rect 222 378 226 382
rect 118 368 122 372
rect 126 368 130 372
rect 142 368 146 372
rect 102 338 106 342
rect 126 338 130 342
rect 126 318 130 322
rect 174 348 178 352
rect 190 348 194 352
rect 230 348 234 352
rect 278 478 282 482
rect 366 658 370 662
rect 342 648 346 652
rect 342 638 346 642
rect 358 638 362 642
rect 334 498 338 502
rect 294 488 298 492
rect 318 468 322 472
rect 302 458 306 462
rect 270 418 274 422
rect 262 408 266 412
rect 294 448 298 452
rect 302 448 306 452
rect 286 438 290 442
rect 406 938 410 942
rect 438 1048 442 1052
rect 498 1003 502 1007
rect 505 1003 509 1007
rect 454 978 458 982
rect 478 968 482 972
rect 494 968 498 972
rect 510 958 514 962
rect 446 948 450 952
rect 470 948 474 952
rect 446 928 450 932
rect 438 908 442 912
rect 446 898 450 902
rect 430 878 434 882
rect 438 868 442 872
rect 430 758 434 762
rect 406 718 410 722
rect 422 718 426 722
rect 414 708 418 712
rect 406 698 410 702
rect 446 758 450 762
rect 494 938 498 942
rect 534 1128 538 1132
rect 526 1078 530 1082
rect 550 1048 554 1052
rect 646 1148 650 1152
rect 670 1148 674 1152
rect 606 1138 610 1142
rect 622 1118 626 1122
rect 614 1108 618 1112
rect 710 1208 714 1212
rect 718 1178 722 1182
rect 702 1158 706 1162
rect 694 1148 698 1152
rect 718 1148 722 1152
rect 670 1108 674 1112
rect 678 1108 682 1112
rect 598 1088 602 1092
rect 582 1068 586 1072
rect 598 1058 602 1062
rect 574 988 578 992
rect 614 1038 618 1042
rect 622 988 626 992
rect 558 958 562 962
rect 550 938 554 942
rect 518 928 522 932
rect 462 908 466 912
rect 486 858 490 862
rect 502 859 506 863
rect 550 858 554 862
rect 498 803 502 807
rect 505 803 509 807
rect 470 758 474 762
rect 526 748 530 752
rect 454 738 458 742
rect 454 708 458 712
rect 438 698 442 702
rect 414 688 418 692
rect 502 738 506 742
rect 478 678 482 682
rect 534 678 538 682
rect 518 668 522 672
rect 390 638 394 642
rect 398 638 402 642
rect 366 628 370 632
rect 390 598 394 602
rect 390 578 394 582
rect 358 558 362 562
rect 478 658 482 662
rect 526 648 530 652
rect 686 1088 690 1092
rect 662 1078 666 1082
rect 654 978 658 982
rect 702 1088 706 1092
rect 702 1078 706 1082
rect 678 1058 682 1062
rect 670 1048 674 1052
rect 694 1048 698 1052
rect 630 948 634 952
rect 614 938 618 942
rect 598 908 602 912
rect 574 848 578 852
rect 566 838 570 842
rect 566 788 570 792
rect 558 768 562 772
rect 574 748 578 752
rect 558 708 562 712
rect 574 708 578 712
rect 582 708 586 712
rect 550 678 554 682
rect 526 638 530 642
rect 542 638 546 642
rect 422 598 426 602
rect 498 603 502 607
rect 505 603 509 607
rect 622 898 626 902
rect 646 878 650 882
rect 734 1198 738 1202
rect 966 1528 970 1532
rect 886 1478 890 1482
rect 902 1478 906 1482
rect 902 1458 906 1462
rect 998 1558 1002 1562
rect 1006 1548 1010 1552
rect 1046 1548 1050 1552
rect 1054 1548 1058 1552
rect 990 1538 994 1542
rect 1006 1528 1010 1532
rect 1002 1503 1006 1507
rect 1009 1503 1013 1507
rect 998 1478 1002 1482
rect 1022 1468 1026 1472
rect 998 1458 1002 1462
rect 902 1448 906 1452
rect 926 1448 930 1452
rect 958 1448 962 1452
rect 990 1448 994 1452
rect 934 1438 938 1442
rect 830 1418 834 1422
rect 894 1388 898 1392
rect 838 1348 842 1352
rect 846 1348 850 1352
rect 926 1378 930 1382
rect 910 1368 914 1372
rect 982 1438 986 1442
rect 966 1388 970 1392
rect 1014 1388 1018 1392
rect 950 1378 954 1382
rect 950 1358 954 1362
rect 974 1368 978 1372
rect 1022 1358 1026 1362
rect 1054 1508 1058 1512
rect 1206 1658 1210 1662
rect 1126 1648 1130 1652
rect 1118 1588 1122 1592
rect 1078 1578 1082 1582
rect 1078 1548 1082 1552
rect 1118 1548 1122 1552
rect 1086 1538 1090 1542
rect 1070 1518 1074 1522
rect 1038 1458 1042 1462
rect 1046 1448 1050 1452
rect 1038 1438 1042 1442
rect 1038 1368 1042 1372
rect 942 1338 946 1342
rect 998 1338 1002 1342
rect 1038 1338 1042 1342
rect 838 1328 842 1332
rect 926 1328 930 1332
rect 942 1328 946 1332
rect 814 1308 818 1312
rect 790 1278 794 1282
rect 862 1318 866 1322
rect 862 1308 866 1312
rect 846 1298 850 1302
rect 894 1298 898 1302
rect 870 1288 874 1292
rect 854 1278 858 1282
rect 942 1318 946 1322
rect 958 1298 962 1302
rect 1534 1908 1538 1912
rect 1742 2058 1746 2062
rect 1726 1988 1730 1992
rect 1710 1978 1714 1982
rect 1702 1938 1706 1942
rect 1550 1878 1554 1882
rect 1638 1878 1642 1882
rect 1502 1868 1506 1872
rect 1566 1868 1570 1872
rect 1630 1858 1634 1862
rect 1686 1858 1690 1862
rect 1686 1848 1690 1852
rect 1478 1788 1482 1792
rect 1422 1758 1426 1762
rect 1446 1748 1450 1752
rect 1390 1738 1394 1742
rect 1630 1828 1634 1832
rect 1566 1808 1570 1812
rect 1522 1803 1526 1807
rect 1529 1803 1533 1807
rect 1574 1778 1578 1782
rect 1502 1748 1506 1752
rect 1454 1718 1458 1722
rect 1358 1668 1362 1672
rect 1254 1648 1258 1652
rect 1142 1598 1146 1602
rect 1134 1588 1138 1592
rect 1150 1558 1154 1562
rect 1158 1558 1162 1562
rect 1206 1558 1210 1562
rect 1270 1558 1274 1562
rect 1214 1548 1218 1552
rect 1222 1548 1226 1552
rect 1190 1538 1194 1542
rect 1294 1538 1298 1542
rect 1158 1528 1162 1532
rect 1206 1528 1210 1532
rect 1238 1518 1242 1522
rect 1110 1468 1114 1472
rect 1134 1468 1138 1472
rect 1078 1458 1082 1462
rect 1102 1458 1106 1462
rect 1094 1448 1098 1452
rect 1070 1438 1074 1442
rect 1102 1368 1106 1372
rect 1078 1358 1082 1362
rect 1110 1358 1114 1362
rect 1062 1348 1066 1352
rect 1002 1303 1006 1307
rect 1009 1303 1013 1307
rect 1022 1298 1026 1302
rect 1046 1298 1050 1302
rect 990 1288 994 1292
rect 910 1278 914 1282
rect 910 1268 914 1272
rect 950 1258 954 1262
rect 878 1248 882 1252
rect 918 1248 922 1252
rect 1038 1248 1042 1252
rect 1054 1248 1058 1252
rect 1022 1238 1026 1242
rect 806 1218 810 1222
rect 982 1218 986 1222
rect 806 1208 810 1212
rect 742 1168 746 1172
rect 758 1168 762 1172
rect 758 1148 762 1152
rect 766 1148 770 1152
rect 782 1148 786 1152
rect 878 1168 882 1172
rect 918 1168 922 1172
rect 902 1148 906 1152
rect 990 1168 994 1172
rect 974 1158 978 1162
rect 854 1138 858 1142
rect 830 1128 834 1132
rect 838 1088 842 1092
rect 742 1078 746 1082
rect 902 1128 906 1132
rect 942 1118 946 1122
rect 918 1068 922 1072
rect 950 1068 954 1072
rect 750 1059 754 1063
rect 694 1028 698 1032
rect 702 948 706 952
rect 958 1048 962 1052
rect 926 1038 930 1042
rect 910 1028 914 1032
rect 870 978 874 982
rect 806 958 810 962
rect 742 938 746 942
rect 798 908 802 912
rect 678 878 682 882
rect 902 958 906 962
rect 918 958 922 962
rect 1014 1168 1018 1172
rect 1002 1103 1006 1107
rect 1009 1103 1013 1107
rect 1030 1158 1034 1162
rect 1134 1428 1138 1432
rect 1326 1568 1330 1572
rect 1318 1558 1322 1562
rect 1326 1538 1330 1542
rect 1150 1478 1154 1482
rect 1230 1478 1234 1482
rect 1246 1478 1250 1482
rect 1270 1478 1274 1482
rect 1310 1478 1314 1482
rect 1150 1458 1154 1462
rect 1174 1458 1178 1462
rect 1190 1458 1194 1462
rect 1206 1458 1210 1462
rect 1174 1448 1178 1452
rect 1190 1448 1194 1452
rect 1198 1438 1202 1442
rect 1142 1388 1146 1392
rect 1342 1598 1346 1602
rect 1414 1658 1418 1662
rect 1382 1628 1386 1632
rect 1478 1638 1482 1642
rect 1446 1618 1450 1622
rect 1454 1618 1458 1622
rect 1366 1598 1370 1602
rect 1366 1578 1370 1582
rect 1358 1568 1362 1572
rect 1374 1568 1378 1572
rect 1406 1568 1410 1572
rect 1358 1548 1362 1552
rect 1414 1558 1418 1562
rect 1398 1548 1402 1552
rect 1398 1538 1402 1542
rect 1350 1528 1354 1532
rect 1334 1488 1338 1492
rect 1326 1478 1330 1482
rect 1430 1498 1434 1502
rect 1382 1488 1386 1492
rect 1438 1488 1442 1492
rect 1430 1478 1434 1482
rect 1278 1468 1282 1472
rect 1262 1438 1266 1442
rect 1214 1408 1218 1412
rect 1222 1408 1226 1412
rect 1166 1368 1170 1372
rect 1158 1358 1162 1362
rect 1174 1358 1178 1362
rect 1206 1358 1210 1362
rect 1134 1348 1138 1352
rect 1158 1348 1162 1352
rect 1174 1348 1178 1352
rect 1206 1348 1210 1352
rect 1086 1338 1090 1342
rect 1126 1338 1130 1342
rect 1070 1328 1074 1332
rect 1094 1328 1098 1332
rect 1118 1328 1122 1332
rect 1158 1328 1162 1332
rect 1190 1328 1194 1332
rect 1086 1318 1090 1322
rect 1102 1318 1106 1322
rect 1086 1278 1090 1282
rect 1086 1268 1090 1272
rect 1062 1238 1066 1242
rect 1110 1288 1114 1292
rect 1118 1288 1122 1292
rect 1126 1288 1130 1292
rect 1214 1298 1218 1302
rect 1198 1278 1202 1282
rect 1182 1268 1186 1272
rect 1142 1258 1146 1262
rect 1094 1198 1098 1202
rect 1118 1198 1122 1202
rect 1150 1238 1154 1242
rect 1182 1238 1186 1242
rect 1206 1258 1210 1262
rect 1270 1408 1274 1412
rect 1302 1458 1306 1462
rect 1318 1458 1322 1462
rect 1374 1458 1378 1462
rect 1302 1448 1306 1452
rect 1326 1448 1330 1452
rect 1310 1418 1314 1422
rect 1286 1388 1290 1392
rect 1230 1368 1234 1372
rect 1246 1368 1250 1372
rect 1246 1358 1250 1362
rect 1254 1358 1258 1362
rect 1262 1358 1266 1362
rect 1238 1348 1242 1352
rect 1254 1318 1258 1322
rect 1238 1298 1242 1302
rect 1254 1298 1258 1302
rect 1286 1338 1290 1342
rect 1334 1358 1338 1362
rect 1358 1348 1362 1352
rect 1310 1338 1314 1342
rect 1382 1368 1386 1372
rect 1390 1368 1394 1372
rect 1582 1768 1586 1772
rect 1590 1768 1594 1772
rect 1606 1758 1610 1762
rect 1598 1748 1602 1752
rect 1638 1778 1642 1782
rect 1694 1818 1698 1822
rect 1686 1768 1690 1772
rect 1582 1738 1586 1742
rect 1534 1688 1538 1692
rect 1550 1678 1554 1682
rect 1598 1678 1602 1682
rect 1598 1668 1602 1672
rect 1606 1668 1610 1672
rect 1574 1658 1578 1662
rect 1622 1658 1626 1662
rect 1526 1648 1530 1652
rect 1494 1608 1498 1612
rect 1522 1603 1526 1607
rect 1529 1603 1533 1607
rect 1614 1638 1618 1642
rect 1614 1628 1618 1632
rect 1662 1728 1666 1732
rect 1678 1718 1682 1722
rect 1686 1708 1690 1712
rect 1654 1698 1658 1702
rect 1790 2059 1794 2063
rect 1758 2038 1762 2042
rect 1934 2148 1938 2152
rect 1854 2088 1858 2092
rect 1886 2078 1890 2082
rect 1918 2078 1922 2082
rect 1886 2068 1890 2072
rect 2094 2408 2098 2412
rect 1998 2348 2002 2352
rect 2070 2347 2074 2351
rect 1982 2278 1986 2282
rect 2026 2303 2030 2307
rect 2033 2303 2037 2307
rect 2046 2298 2050 2302
rect 2014 2248 2018 2252
rect 1998 2198 2002 2202
rect 2126 2508 2130 2512
rect 2142 2478 2146 2482
rect 2110 2468 2114 2472
rect 2118 2348 2122 2352
rect 2134 2348 2138 2352
rect 2350 2928 2354 2932
rect 2230 2898 2234 2902
rect 2238 2888 2242 2892
rect 2214 2868 2218 2872
rect 2198 2778 2202 2782
rect 2254 2778 2258 2782
rect 2182 2688 2186 2692
rect 2182 2648 2186 2652
rect 2302 2908 2306 2912
rect 2326 2858 2330 2862
rect 2310 2848 2314 2852
rect 2294 2778 2298 2782
rect 2286 2748 2290 2752
rect 2254 2728 2258 2732
rect 2222 2678 2226 2682
rect 2246 2678 2250 2682
rect 2286 2678 2290 2682
rect 2238 2668 2242 2672
rect 2230 2628 2234 2632
rect 2238 2598 2242 2602
rect 2214 2568 2218 2572
rect 2238 2568 2242 2572
rect 2174 2498 2178 2502
rect 2174 2468 2178 2472
rect 2174 2358 2178 2362
rect 2150 2338 2154 2342
rect 2286 2668 2290 2672
rect 2262 2648 2266 2652
rect 2246 2518 2250 2522
rect 2206 2498 2210 2502
rect 2206 2448 2210 2452
rect 2222 2448 2226 2452
rect 2222 2348 2226 2352
rect 2230 2348 2234 2352
rect 2198 2338 2202 2342
rect 2182 2318 2186 2322
rect 2166 2308 2170 2312
rect 2158 2298 2162 2302
rect 2158 2278 2162 2282
rect 2158 2228 2162 2232
rect 2198 2298 2202 2302
rect 2206 2278 2210 2282
rect 2214 2278 2218 2282
rect 2246 2488 2250 2492
rect 2270 2488 2274 2492
rect 2262 2468 2266 2472
rect 2254 2458 2258 2462
rect 2246 2438 2250 2442
rect 2246 2368 2250 2372
rect 2382 2938 2386 2942
rect 2414 3148 2418 3152
rect 2478 3148 2482 3152
rect 2598 3178 2602 3182
rect 2614 3238 2618 3242
rect 2670 3258 2674 3262
rect 2710 3258 2714 3262
rect 2750 3258 2754 3262
rect 2646 3248 2650 3252
rect 2678 3248 2682 3252
rect 2638 3238 2642 3242
rect 2622 3208 2626 3212
rect 2630 3158 2634 3162
rect 2622 3148 2626 3152
rect 2462 3138 2466 3142
rect 2510 3138 2514 3142
rect 2598 3138 2602 3142
rect 2614 3138 2618 3142
rect 2430 3128 2434 3132
rect 2494 3128 2498 3132
rect 2526 3128 2530 3132
rect 2470 3118 2474 3122
rect 2478 3118 2482 3122
rect 2414 3108 2418 3112
rect 2542 3118 2546 3122
rect 2414 3068 2418 3072
rect 2438 3068 2442 3072
rect 2478 3068 2482 3072
rect 2422 3058 2426 3062
rect 2406 3008 2410 3012
rect 2414 2968 2418 2972
rect 2454 3058 2458 3062
rect 2438 3038 2442 3042
rect 2470 3048 2474 3052
rect 2510 3108 2514 3112
rect 2526 3078 2530 3082
rect 2518 3068 2522 3072
rect 2518 3048 2522 3052
rect 2430 2948 2434 2952
rect 2462 2948 2466 2952
rect 2486 2938 2490 2942
rect 2382 2928 2386 2932
rect 2398 2928 2402 2932
rect 2366 2898 2370 2902
rect 2374 2868 2378 2872
rect 2438 2918 2442 2922
rect 2446 2918 2450 2922
rect 2398 2908 2402 2912
rect 2414 2908 2418 2912
rect 2430 2908 2434 2912
rect 2430 2888 2434 2892
rect 2438 2868 2442 2872
rect 2422 2858 2426 2862
rect 2406 2848 2410 2852
rect 2478 2928 2482 2932
rect 2470 2858 2474 2862
rect 2454 2838 2458 2842
rect 2310 2748 2314 2752
rect 2334 2748 2338 2752
rect 2446 2748 2450 2752
rect 2334 2738 2338 2742
rect 2350 2738 2354 2742
rect 2366 2738 2370 2742
rect 2382 2738 2386 2742
rect 2406 2738 2410 2742
rect 2318 2708 2322 2712
rect 2302 2658 2306 2662
rect 2302 2628 2306 2632
rect 2334 2668 2338 2672
rect 2406 2718 2410 2722
rect 2374 2698 2378 2702
rect 2382 2688 2386 2692
rect 2350 2658 2354 2662
rect 2318 2568 2322 2572
rect 2310 2548 2314 2552
rect 2318 2548 2322 2552
rect 2294 2508 2298 2512
rect 2286 2498 2290 2502
rect 2318 2418 2322 2422
rect 2302 2398 2306 2402
rect 2358 2648 2362 2652
rect 2382 2628 2386 2632
rect 2446 2708 2450 2712
rect 2430 2648 2434 2652
rect 2358 2608 2362 2612
rect 2422 2608 2426 2612
rect 2390 2588 2394 2592
rect 2358 2558 2362 2562
rect 2430 2558 2434 2562
rect 2478 2828 2482 2832
rect 2502 2948 2506 2952
rect 2518 2948 2522 2952
rect 2510 2928 2514 2932
rect 2582 3098 2586 3102
rect 2558 3068 2562 3072
rect 2598 3068 2602 3072
rect 2606 3068 2610 3072
rect 2550 3058 2554 3062
rect 2566 3058 2570 3062
rect 2534 3028 2538 3032
rect 2546 3003 2550 3007
rect 2553 3003 2557 3007
rect 2534 2948 2538 2952
rect 2606 3048 2610 3052
rect 2590 3038 2594 3042
rect 2590 2978 2594 2982
rect 2566 2938 2570 2942
rect 2526 2888 2530 2892
rect 2630 3048 2634 3052
rect 2710 3238 2714 3242
rect 2678 3208 2682 3212
rect 2694 3208 2698 3212
rect 2654 3158 2658 3162
rect 2670 3158 2674 3162
rect 2646 3148 2650 3152
rect 2662 3138 2666 3142
rect 2646 3108 2650 3112
rect 2646 3068 2650 3072
rect 2646 3058 2650 3062
rect 2678 3128 2682 3132
rect 2694 3108 2698 3112
rect 2702 3098 2706 3102
rect 2678 3078 2682 3082
rect 2662 3048 2666 3052
rect 2678 3048 2682 3052
rect 2766 3248 2770 3252
rect 2742 3218 2746 3222
rect 2750 3218 2754 3222
rect 2734 3208 2738 3212
rect 2726 3198 2730 3202
rect 2822 3238 2826 3242
rect 2806 3218 2810 3222
rect 2822 3208 2826 3212
rect 2798 3198 2802 3202
rect 2814 3188 2818 3192
rect 2774 3168 2778 3172
rect 2782 3168 2786 3172
rect 2742 3138 2746 3142
rect 2806 3138 2810 3142
rect 2742 3118 2746 3122
rect 2734 3108 2738 3112
rect 2750 3108 2754 3112
rect 2734 3098 2738 3102
rect 2710 3048 2714 3052
rect 2702 3038 2706 3042
rect 2726 3038 2730 3042
rect 2798 3128 2802 3132
rect 2766 3118 2770 3122
rect 2774 3108 2778 3112
rect 2742 3048 2746 3052
rect 2758 3018 2762 3022
rect 2758 2988 2762 2992
rect 2750 2958 2754 2962
rect 2686 2948 2690 2952
rect 2606 2938 2610 2942
rect 2630 2938 2634 2942
rect 2670 2938 2674 2942
rect 2710 2938 2714 2942
rect 2630 2878 2634 2882
rect 2502 2868 2506 2872
rect 2614 2868 2618 2872
rect 2534 2858 2538 2862
rect 2566 2858 2570 2862
rect 2606 2858 2610 2862
rect 2622 2858 2626 2862
rect 2546 2803 2550 2807
rect 2553 2803 2557 2807
rect 2614 2848 2618 2852
rect 2598 2838 2602 2842
rect 2574 2798 2578 2802
rect 2494 2778 2498 2782
rect 2518 2778 2522 2782
rect 2542 2768 2546 2772
rect 2614 2768 2618 2772
rect 2486 2758 2490 2762
rect 2670 2908 2674 2912
rect 2670 2898 2674 2902
rect 2646 2858 2650 2862
rect 2638 2828 2642 2832
rect 2678 2858 2682 2862
rect 2670 2838 2674 2842
rect 2702 2828 2706 2832
rect 2710 2808 2714 2812
rect 2694 2758 2698 2762
rect 2702 2758 2706 2762
rect 2622 2748 2626 2752
rect 2726 2868 2730 2872
rect 2758 2948 2762 2952
rect 2766 2948 2770 2952
rect 2758 2918 2762 2922
rect 2758 2868 2762 2872
rect 2734 2848 2738 2852
rect 2766 2848 2770 2852
rect 2774 2848 2778 2852
rect 2734 2838 2738 2842
rect 2870 3258 2874 3262
rect 2854 3248 2858 3252
rect 2846 3238 2850 3242
rect 2862 3218 2866 3222
rect 2854 3208 2858 3212
rect 2838 3168 2842 3172
rect 2918 3248 2922 3252
rect 2894 3238 2898 3242
rect 2878 3188 2882 3192
rect 2870 3148 2874 3152
rect 2886 3138 2890 3142
rect 2838 3128 2842 3132
rect 2830 3098 2834 3102
rect 2846 3118 2850 3122
rect 2878 3128 2882 3132
rect 2886 3118 2890 3122
rect 2902 3208 2906 3212
rect 2918 3168 2922 3172
rect 2982 3268 2986 3272
rect 3062 3268 3066 3272
rect 2942 3258 2946 3262
rect 2966 3258 2970 3262
rect 2990 3258 2994 3262
rect 2942 3248 2946 3252
rect 3006 3248 3010 3252
rect 2966 3208 2970 3212
rect 2990 3198 2994 3202
rect 3022 3248 3026 3252
rect 3014 3238 3018 3242
rect 3038 3208 3042 3212
rect 3022 3168 3026 3172
rect 3086 3348 3090 3352
rect 3118 3378 3122 3382
rect 3190 3388 3194 3392
rect 3166 3378 3170 3382
rect 3134 3358 3138 3362
rect 3150 3358 3154 3362
rect 3174 3358 3178 3362
rect 3110 3348 3114 3352
rect 3126 3318 3130 3322
rect 3102 3288 3106 3292
rect 3094 3278 3098 3282
rect 3102 3268 3106 3272
rect 3078 3258 3082 3262
rect 3126 3308 3130 3312
rect 3142 3308 3146 3312
rect 3206 3328 3210 3332
rect 3166 3308 3170 3312
rect 3182 3308 3186 3312
rect 3150 3278 3154 3282
rect 3134 3258 3138 3262
rect 3118 3248 3122 3252
rect 3086 3238 3090 3242
rect 3110 3208 3114 3212
rect 3102 3168 3106 3172
rect 2942 3138 2946 3142
rect 2974 3138 2978 3142
rect 3014 3138 3018 3142
rect 3054 3138 3058 3142
rect 2934 3128 2938 3132
rect 2846 3088 2850 3092
rect 2854 3088 2858 3092
rect 2790 3038 2794 3042
rect 2798 2958 2802 2962
rect 2806 2928 2810 2932
rect 2878 3058 2882 3062
rect 2894 3098 2898 3102
rect 2910 3078 2914 3082
rect 2894 3068 2898 3072
rect 2910 3058 2914 3062
rect 2918 3048 2922 3052
rect 2838 3038 2842 3042
rect 2862 3038 2866 3042
rect 2822 3028 2826 3032
rect 2838 3028 2842 3032
rect 2902 3028 2906 3032
rect 2886 2998 2890 3002
rect 2838 2938 2842 2942
rect 2814 2898 2818 2902
rect 2806 2828 2810 2832
rect 2838 2858 2842 2862
rect 2862 2868 2866 2872
rect 2838 2848 2842 2852
rect 2846 2768 2850 2772
rect 2766 2758 2770 2762
rect 2814 2758 2818 2762
rect 2462 2738 2466 2742
rect 2598 2738 2602 2742
rect 2646 2738 2650 2742
rect 2694 2738 2698 2742
rect 2726 2738 2730 2742
rect 2734 2738 2738 2742
rect 2478 2698 2482 2702
rect 2454 2688 2458 2692
rect 2478 2688 2482 2692
rect 2590 2718 2594 2722
rect 2542 2668 2546 2672
rect 2566 2658 2570 2662
rect 2550 2648 2554 2652
rect 2518 2608 2522 2612
rect 2546 2603 2550 2607
rect 2553 2603 2557 2607
rect 2582 2648 2586 2652
rect 2566 2598 2570 2602
rect 2542 2588 2546 2592
rect 2454 2568 2458 2572
rect 2462 2558 2466 2562
rect 2462 2548 2466 2552
rect 2614 2708 2618 2712
rect 2678 2708 2682 2712
rect 2630 2698 2634 2702
rect 2662 2698 2666 2702
rect 2606 2678 2610 2682
rect 2670 2648 2674 2652
rect 2606 2558 2610 2562
rect 2662 2558 2666 2562
rect 2438 2538 2442 2542
rect 2358 2518 2362 2522
rect 2350 2488 2354 2492
rect 2390 2448 2394 2452
rect 2558 2528 2562 2532
rect 2654 2528 2658 2532
rect 2510 2488 2514 2492
rect 2518 2478 2522 2482
rect 2574 2478 2578 2482
rect 2590 2478 2594 2482
rect 2454 2468 2458 2472
rect 2502 2468 2506 2472
rect 2510 2468 2514 2472
rect 2574 2468 2578 2472
rect 2630 2468 2634 2472
rect 2478 2448 2482 2452
rect 2422 2438 2426 2442
rect 2342 2408 2346 2412
rect 2318 2388 2322 2392
rect 2342 2388 2346 2392
rect 2278 2358 2282 2362
rect 2310 2358 2314 2362
rect 2254 2348 2258 2352
rect 2278 2348 2282 2352
rect 2334 2358 2338 2362
rect 2374 2368 2378 2372
rect 2406 2358 2410 2362
rect 2390 2338 2394 2342
rect 2302 2328 2306 2332
rect 2366 2328 2370 2332
rect 2246 2308 2250 2312
rect 2262 2288 2266 2292
rect 2278 2268 2282 2272
rect 2182 2248 2186 2252
rect 2230 2248 2234 2252
rect 2246 2248 2250 2252
rect 2214 2188 2218 2192
rect 2110 2168 2114 2172
rect 1998 2138 2002 2142
rect 2014 2118 2018 2122
rect 1966 2078 1970 2082
rect 1990 2078 1994 2082
rect 2026 2103 2030 2107
rect 2033 2103 2037 2107
rect 2094 2068 2098 2072
rect 1830 2058 1834 2062
rect 1990 2058 1994 2062
rect 2102 2058 2106 2062
rect 2046 2038 2050 2042
rect 1862 2028 1866 2032
rect 1806 2018 1810 2022
rect 1822 1998 1826 2002
rect 1854 1978 1858 1982
rect 1758 1968 1762 1972
rect 1854 1968 1858 1972
rect 1774 1958 1778 1962
rect 1798 1958 1802 1962
rect 1734 1948 1738 1952
rect 1750 1948 1754 1952
rect 1726 1878 1730 1882
rect 1718 1868 1722 1872
rect 1766 1878 1770 1882
rect 1798 1928 1802 1932
rect 1806 1878 1810 1882
rect 1742 1868 1746 1872
rect 1782 1868 1786 1872
rect 1798 1868 1802 1872
rect 1830 1938 1834 1942
rect 1822 1928 1826 1932
rect 1750 1858 1754 1862
rect 1734 1848 1738 1852
rect 1774 1848 1778 1852
rect 1814 1848 1818 1852
rect 1830 1848 1834 1852
rect 1894 2008 1898 2012
rect 1894 1968 1898 1972
rect 1934 1968 1938 1972
rect 1870 1938 1874 1942
rect 1870 1928 1874 1932
rect 1902 1938 1906 1942
rect 1934 1938 1938 1942
rect 1934 1928 1938 1932
rect 1886 1908 1890 1912
rect 1886 1888 1890 1892
rect 1862 1858 1866 1862
rect 1846 1828 1850 1832
rect 1782 1808 1786 1812
rect 1758 1798 1762 1802
rect 1726 1788 1730 1792
rect 1718 1768 1722 1772
rect 1742 1768 1746 1772
rect 1822 1768 1826 1772
rect 1854 1768 1858 1772
rect 1782 1748 1786 1752
rect 1774 1738 1778 1742
rect 1942 1918 1946 1922
rect 1918 1878 1922 1882
rect 1934 1878 1938 1882
rect 1894 1858 1898 1862
rect 1918 1858 1922 1862
rect 1894 1848 1898 1852
rect 1926 1808 1930 1812
rect 2054 2008 2058 2012
rect 2102 1998 2106 2002
rect 2086 1978 2090 1982
rect 1958 1968 1962 1972
rect 2006 1968 2010 1972
rect 2062 1968 2066 1972
rect 1950 1898 1954 1902
rect 2006 1948 2010 1952
rect 2054 1948 2058 1952
rect 2094 1948 2098 1952
rect 2070 1938 2074 1942
rect 2190 2178 2194 2182
rect 2222 2178 2226 2182
rect 2230 2178 2234 2182
rect 2246 2178 2250 2182
rect 2254 2178 2258 2182
rect 2270 2158 2274 2162
rect 2206 2148 2210 2152
rect 2230 2148 2234 2152
rect 2326 2288 2330 2292
rect 2454 2378 2458 2382
rect 2478 2358 2482 2362
rect 2446 2348 2450 2352
rect 2422 2338 2426 2342
rect 2454 2338 2458 2342
rect 2470 2328 2474 2332
rect 2406 2308 2410 2312
rect 2350 2298 2354 2302
rect 2398 2288 2402 2292
rect 2334 2268 2338 2272
rect 2358 2268 2362 2272
rect 2382 2268 2386 2272
rect 2398 2248 2402 2252
rect 2310 2238 2314 2242
rect 2582 2458 2586 2462
rect 2526 2448 2530 2452
rect 2598 2448 2602 2452
rect 2638 2438 2642 2442
rect 2546 2403 2550 2407
rect 2553 2403 2557 2407
rect 2582 2358 2586 2362
rect 2726 2708 2730 2712
rect 2726 2668 2730 2672
rect 2702 2658 2706 2662
rect 2718 2648 2722 2652
rect 2806 2738 2810 2742
rect 2830 2738 2834 2742
rect 2814 2718 2818 2722
rect 2766 2628 2770 2632
rect 2750 2578 2754 2582
rect 2758 2578 2762 2582
rect 2686 2568 2690 2572
rect 2742 2548 2746 2552
rect 2678 2538 2682 2542
rect 2742 2528 2746 2532
rect 2750 2528 2754 2532
rect 2830 2698 2834 2702
rect 2846 2678 2850 2682
rect 2886 2908 2890 2912
rect 2942 3118 2946 3122
rect 2910 2958 2914 2962
rect 2886 2778 2890 2782
rect 2934 3028 2938 3032
rect 2982 3128 2986 3132
rect 3030 3098 3034 3102
rect 3030 3078 3034 3082
rect 3086 3118 3090 3122
rect 3050 3103 3054 3107
rect 3057 3103 3061 3107
rect 3054 3088 3058 3092
rect 2990 3068 2994 3072
rect 2974 3048 2978 3052
rect 2974 3038 2978 3042
rect 2926 2958 2930 2962
rect 2982 2938 2986 2942
rect 2958 2918 2962 2922
rect 2958 2908 2962 2912
rect 2966 2878 2970 2882
rect 2950 2858 2954 2862
rect 2926 2848 2930 2852
rect 2950 2838 2954 2842
rect 2942 2828 2946 2832
rect 2982 2868 2986 2872
rect 2974 2848 2978 2852
rect 2982 2838 2986 2842
rect 2998 3058 3002 3062
rect 3022 3058 3026 3062
rect 3006 3048 3010 3052
rect 3030 3048 3034 3052
rect 3014 3038 3018 3042
rect 3030 3038 3034 3042
rect 3046 3038 3050 3042
rect 3022 2968 3026 2972
rect 3038 3028 3042 3032
rect 3094 3108 3098 3112
rect 3070 3078 3074 3082
rect 3094 3078 3098 3082
rect 3078 3068 3082 3072
rect 3062 3058 3066 3062
rect 3110 3058 3114 3062
rect 3110 3048 3114 3052
rect 3134 3208 3138 3212
rect 3158 3208 3162 3212
rect 3158 3178 3162 3182
rect 3150 3168 3154 3172
rect 3182 3268 3186 3272
rect 3310 3408 3314 3412
rect 3294 3358 3298 3362
rect 3430 3428 3434 3432
rect 3398 3398 3402 3402
rect 3406 3388 3410 3392
rect 3366 3368 3370 3372
rect 3358 3358 3362 3362
rect 3238 3348 3242 3352
rect 3262 3348 3266 3352
rect 3278 3348 3282 3352
rect 3310 3338 3314 3342
rect 3318 3338 3322 3342
rect 3246 3318 3250 3322
rect 3230 3308 3234 3312
rect 3222 3298 3226 3302
rect 3262 3328 3266 3332
rect 3246 3278 3250 3282
rect 3214 3258 3218 3262
rect 3214 3248 3218 3252
rect 3174 3238 3178 3242
rect 3198 3238 3202 3242
rect 3230 3258 3234 3262
rect 3254 3258 3258 3262
rect 3222 3218 3226 3222
rect 3230 3198 3234 3202
rect 3222 3188 3226 3192
rect 3182 3178 3186 3182
rect 3222 3178 3226 3182
rect 3166 3168 3170 3172
rect 3126 3088 3130 3092
rect 3118 3038 3122 3042
rect 3102 2988 3106 2992
rect 3166 3118 3170 3122
rect 3182 3128 3186 3132
rect 3254 3168 3258 3172
rect 3238 3148 3242 3152
rect 3254 3148 3258 3152
rect 3246 3138 3250 3142
rect 3230 3088 3234 3092
rect 3158 3078 3162 3082
rect 3174 3078 3178 3082
rect 3214 3078 3218 3082
rect 3198 3068 3202 3072
rect 3182 3058 3186 3062
rect 3214 3058 3218 3062
rect 3142 3048 3146 3052
rect 3182 3048 3186 3052
rect 3190 3048 3194 3052
rect 3142 2998 3146 3002
rect 3222 3048 3226 3052
rect 3254 3118 3258 3122
rect 3238 3058 3242 3062
rect 3238 3048 3242 3052
rect 3326 3328 3330 3332
rect 3310 3318 3314 3322
rect 3302 3298 3306 3302
rect 3366 3348 3370 3352
rect 3374 3348 3378 3352
rect 3398 3348 3402 3352
rect 3430 3348 3434 3352
rect 3342 3338 3346 3342
rect 3366 3338 3370 3342
rect 3406 3338 3410 3342
rect 3294 3268 3298 3272
rect 3278 3258 3282 3262
rect 3286 3248 3290 3252
rect 3310 3248 3314 3252
rect 3350 3328 3354 3332
rect 3342 3278 3346 3282
rect 3350 3278 3354 3282
rect 3366 3228 3370 3232
rect 3278 3158 3282 3162
rect 3382 3328 3386 3332
rect 3390 3288 3394 3292
rect 3286 3148 3290 3152
rect 3302 3148 3306 3152
rect 3350 3148 3354 3152
rect 3374 3148 3378 3152
rect 3358 3138 3362 3142
rect 3310 3128 3314 3132
rect 3294 3108 3298 3112
rect 3270 3088 3274 3092
rect 3326 3078 3330 3082
rect 3278 3068 3282 3072
rect 3294 3068 3298 3072
rect 3270 3048 3274 3052
rect 3286 2998 3290 3002
rect 3270 2988 3274 2992
rect 3230 2958 3234 2962
rect 3038 2938 3042 2942
rect 3094 2938 3098 2942
rect 3134 2938 3138 2942
rect 3174 2938 3178 2942
rect 2998 2928 3002 2932
rect 3006 2928 3010 2932
rect 3030 2928 3034 2932
rect 3006 2848 3010 2852
rect 2870 2768 2874 2772
rect 2934 2768 2938 2772
rect 2958 2768 2962 2772
rect 2966 2768 2970 2772
rect 2934 2748 2938 2752
rect 2862 2738 2866 2742
rect 2886 2738 2890 2742
rect 2886 2668 2890 2672
rect 2902 2668 2906 2672
rect 2910 2658 2914 2662
rect 2822 2648 2826 2652
rect 2838 2648 2842 2652
rect 2798 2548 2802 2552
rect 2790 2538 2794 2542
rect 2758 2478 2762 2482
rect 2774 2468 2778 2472
rect 2678 2418 2682 2422
rect 2598 2348 2602 2352
rect 2654 2348 2658 2352
rect 2710 2348 2714 2352
rect 2486 2338 2490 2342
rect 2526 2338 2530 2342
rect 2534 2298 2538 2302
rect 2518 2288 2522 2292
rect 2654 2328 2658 2332
rect 2614 2318 2618 2322
rect 2718 2318 2722 2322
rect 2566 2288 2570 2292
rect 2502 2268 2506 2272
rect 2430 2228 2434 2232
rect 2478 2228 2482 2232
rect 2366 2178 2370 2182
rect 2398 2178 2402 2182
rect 2310 2158 2314 2162
rect 2374 2158 2378 2162
rect 2422 2158 2426 2162
rect 2510 2218 2514 2222
rect 2438 2188 2442 2192
rect 2454 2158 2458 2162
rect 2286 2148 2290 2152
rect 2310 2148 2314 2152
rect 2326 2148 2330 2152
rect 2350 2148 2354 2152
rect 2438 2148 2442 2152
rect 2454 2148 2458 2152
rect 2462 2148 2466 2152
rect 2534 2208 2538 2212
rect 2546 2203 2550 2207
rect 2553 2203 2557 2207
rect 2686 2298 2690 2302
rect 2630 2288 2634 2292
rect 2678 2288 2682 2292
rect 2598 2258 2602 2262
rect 2630 2258 2634 2262
rect 2638 2258 2642 2262
rect 2574 2248 2578 2252
rect 2606 2248 2610 2252
rect 2614 2248 2618 2252
rect 2606 2228 2610 2232
rect 2606 2208 2610 2212
rect 2630 2208 2634 2212
rect 2598 2158 2602 2162
rect 2670 2268 2674 2272
rect 2758 2458 2762 2462
rect 2734 2448 2738 2452
rect 2790 2468 2794 2472
rect 2822 2568 2826 2572
rect 2854 2568 2858 2572
rect 2862 2558 2866 2562
rect 2870 2548 2874 2552
rect 2838 2508 2842 2512
rect 2854 2508 2858 2512
rect 2806 2478 2810 2482
rect 2878 2478 2882 2482
rect 2774 2388 2778 2392
rect 2798 2388 2802 2392
rect 2758 2368 2762 2372
rect 2758 2348 2762 2352
rect 2782 2348 2786 2352
rect 2854 2448 2858 2452
rect 2974 2758 2978 2762
rect 2918 2648 2922 2652
rect 2910 2548 2914 2552
rect 2902 2418 2906 2422
rect 2878 2398 2882 2402
rect 2870 2368 2874 2372
rect 2806 2358 2810 2362
rect 2862 2358 2866 2362
rect 2814 2348 2818 2352
rect 2838 2348 2842 2352
rect 2734 2338 2738 2342
rect 2742 2338 2746 2342
rect 2838 2318 2842 2322
rect 2742 2308 2746 2312
rect 2766 2308 2770 2312
rect 2774 2298 2778 2302
rect 2726 2288 2730 2292
rect 2758 2278 2762 2282
rect 2734 2258 2738 2262
rect 2686 2248 2690 2252
rect 2710 2248 2714 2252
rect 2782 2278 2786 2282
rect 2814 2278 2818 2282
rect 2902 2358 2906 2362
rect 2902 2348 2906 2352
rect 2854 2298 2858 2302
rect 2862 2298 2866 2302
rect 2894 2278 2898 2282
rect 2838 2258 2842 2262
rect 2774 2248 2778 2252
rect 2790 2248 2794 2252
rect 2878 2258 2882 2262
rect 2894 2258 2898 2262
rect 2878 2248 2882 2252
rect 2758 2238 2762 2242
rect 2806 2238 2810 2242
rect 2862 2238 2866 2242
rect 2886 2238 2890 2242
rect 2654 2228 2658 2232
rect 2750 2228 2754 2232
rect 2758 2228 2762 2232
rect 2838 2228 2842 2232
rect 2654 2158 2658 2162
rect 2670 2158 2674 2162
rect 2686 2158 2690 2162
rect 2734 2158 2738 2162
rect 2686 2148 2690 2152
rect 2198 2138 2202 2142
rect 2246 2138 2250 2142
rect 2286 2138 2290 2142
rect 2318 2138 2322 2142
rect 2406 2138 2410 2142
rect 2638 2138 2642 2142
rect 2654 2138 2658 2142
rect 2678 2138 2682 2142
rect 2710 2138 2714 2142
rect 2230 2118 2234 2122
rect 2230 2098 2234 2102
rect 2166 2078 2170 2082
rect 2222 2078 2226 2082
rect 2118 2059 2122 2063
rect 2166 2048 2170 2052
rect 2190 2048 2194 2052
rect 2198 2048 2202 2052
rect 2214 1998 2218 2002
rect 2198 1978 2202 1982
rect 2134 1948 2138 1952
rect 2150 1948 2154 1952
rect 2118 1938 2122 1942
rect 2014 1928 2018 1932
rect 1998 1918 2002 1922
rect 2110 1918 2114 1922
rect 1982 1908 1986 1912
rect 2026 1903 2030 1907
rect 2033 1903 2037 1907
rect 2182 1938 2186 1942
rect 2158 1908 2162 1912
rect 2182 1908 2186 1912
rect 2142 1898 2146 1902
rect 2078 1888 2082 1892
rect 1974 1878 1978 1882
rect 1942 1828 1946 1832
rect 1910 1788 1914 1792
rect 1886 1768 1890 1772
rect 1902 1768 1906 1772
rect 1934 1788 1938 1792
rect 1966 1788 1970 1792
rect 1950 1758 1954 1762
rect 1710 1728 1714 1732
rect 1718 1728 1722 1732
rect 1726 1728 1730 1732
rect 1798 1728 1802 1732
rect 1830 1728 1834 1732
rect 1878 1728 1882 1732
rect 1702 1698 1706 1702
rect 1694 1688 1698 1692
rect 1750 1668 1754 1672
rect 1614 1608 1618 1612
rect 1630 1608 1634 1612
rect 1606 1598 1610 1602
rect 1534 1568 1538 1572
rect 1550 1568 1554 1572
rect 1574 1568 1578 1572
rect 1486 1538 1490 1542
rect 1470 1528 1474 1532
rect 1518 1538 1522 1542
rect 1494 1518 1498 1522
rect 1462 1468 1466 1472
rect 1478 1498 1482 1502
rect 1502 1498 1506 1502
rect 1470 1458 1474 1462
rect 1662 1638 1666 1642
rect 1638 1598 1642 1602
rect 1670 1568 1674 1572
rect 1638 1558 1642 1562
rect 1654 1548 1658 1552
rect 1542 1528 1546 1532
rect 1558 1528 1562 1532
rect 1606 1528 1610 1532
rect 1566 1518 1570 1522
rect 1630 1518 1634 1522
rect 1542 1478 1546 1482
rect 1486 1468 1490 1472
rect 1510 1468 1514 1472
rect 1558 1468 1562 1472
rect 1534 1458 1538 1462
rect 1606 1508 1610 1512
rect 1582 1498 1586 1502
rect 1622 1498 1626 1502
rect 1566 1458 1570 1462
rect 1486 1418 1490 1422
rect 1550 1418 1554 1422
rect 1454 1358 1458 1362
rect 1398 1338 1402 1342
rect 1414 1338 1418 1342
rect 1310 1328 1314 1332
rect 1286 1258 1290 1262
rect 1230 1248 1234 1252
rect 1310 1318 1314 1322
rect 1302 1278 1306 1282
rect 1422 1328 1426 1332
rect 1374 1298 1378 1302
rect 1310 1248 1314 1252
rect 1326 1238 1330 1242
rect 1294 1218 1298 1222
rect 1198 1198 1202 1202
rect 1326 1198 1330 1202
rect 1086 1168 1090 1172
rect 1174 1168 1178 1172
rect 1262 1168 1266 1172
rect 1062 1158 1066 1162
rect 1094 1158 1098 1162
rect 1118 1158 1122 1162
rect 1158 1158 1162 1162
rect 1230 1158 1234 1162
rect 1062 1148 1066 1152
rect 1078 1148 1082 1152
rect 1070 1138 1074 1142
rect 1102 1138 1106 1142
rect 1022 1078 1026 1082
rect 982 1058 986 1062
rect 998 1048 1002 1052
rect 974 1038 978 1042
rect 1118 1128 1122 1132
rect 1134 1148 1138 1152
rect 1206 1148 1210 1152
rect 1246 1148 1250 1152
rect 1302 1148 1306 1152
rect 1318 1148 1322 1152
rect 1142 1138 1146 1142
rect 1222 1138 1226 1142
rect 1238 1128 1242 1132
rect 1294 1128 1298 1132
rect 1038 1118 1042 1122
rect 1126 1118 1130 1122
rect 1230 1118 1234 1122
rect 1214 1108 1218 1112
rect 1118 1098 1122 1102
rect 1158 1098 1162 1102
rect 1046 1088 1050 1092
rect 1062 1078 1066 1082
rect 1070 1078 1074 1082
rect 1126 1088 1130 1092
rect 1142 1088 1146 1092
rect 1190 1078 1194 1082
rect 1174 1068 1178 1072
rect 1214 1068 1218 1072
rect 1038 1048 1042 1052
rect 1238 1108 1242 1112
rect 1174 1058 1178 1062
rect 1190 1058 1194 1062
rect 1030 1028 1034 1032
rect 1062 1028 1066 1032
rect 1142 1028 1146 1032
rect 974 998 978 1002
rect 1086 1018 1090 1022
rect 1126 978 1130 982
rect 1046 968 1050 972
rect 950 958 954 962
rect 974 958 978 962
rect 1022 958 1026 962
rect 926 948 930 952
rect 958 938 962 942
rect 990 938 994 942
rect 878 928 882 932
rect 878 918 882 922
rect 854 898 858 902
rect 950 898 954 902
rect 934 878 938 882
rect 966 888 970 892
rect 670 868 674 872
rect 694 868 698 872
rect 726 868 730 872
rect 742 868 746 872
rect 710 858 714 862
rect 822 859 826 863
rect 950 858 954 862
rect 662 848 666 852
rect 702 848 706 852
rect 734 848 738 852
rect 694 838 698 842
rect 726 828 730 832
rect 774 818 778 822
rect 646 808 650 812
rect 758 808 762 812
rect 630 768 634 772
rect 678 768 682 772
rect 870 808 874 812
rect 910 808 914 812
rect 702 758 706 762
rect 710 758 714 762
rect 638 748 642 752
rect 670 748 674 752
rect 702 738 706 742
rect 638 708 642 712
rect 630 688 634 692
rect 590 648 594 652
rect 614 648 618 652
rect 454 548 458 552
rect 662 698 666 702
rect 654 688 658 692
rect 670 688 674 692
rect 1002 903 1006 907
rect 1009 903 1013 907
rect 982 888 986 892
rect 1030 868 1034 872
rect 974 848 978 852
rect 1078 958 1082 962
rect 1054 948 1058 952
rect 1078 948 1082 952
rect 1214 1018 1218 1022
rect 1198 998 1202 1002
rect 1142 958 1146 962
rect 1150 958 1154 962
rect 1166 958 1170 962
rect 1182 958 1186 962
rect 1214 958 1218 962
rect 1054 898 1058 902
rect 1086 878 1090 882
rect 1038 838 1042 842
rect 1118 898 1122 902
rect 1158 948 1162 952
rect 1302 1098 1306 1102
rect 1358 1248 1362 1252
rect 1374 1248 1378 1252
rect 1366 1188 1370 1192
rect 1358 1158 1362 1162
rect 1350 1148 1354 1152
rect 1358 1118 1362 1122
rect 1342 1108 1346 1112
rect 1262 1088 1266 1092
rect 1294 1088 1298 1092
rect 1358 1088 1362 1092
rect 1310 1068 1314 1072
rect 1294 1058 1298 1062
rect 1318 1058 1322 1062
rect 1270 1048 1274 1052
rect 1302 1038 1306 1042
rect 1302 1028 1306 1032
rect 1278 1018 1282 1022
rect 1270 958 1274 962
rect 1262 948 1266 952
rect 1222 938 1226 942
rect 1230 938 1234 942
rect 1150 898 1154 902
rect 1142 888 1146 892
rect 1134 878 1138 882
rect 1142 868 1146 872
rect 1110 858 1114 862
rect 1102 818 1106 822
rect 1078 798 1082 802
rect 958 788 962 792
rect 750 748 754 752
rect 870 751 874 752
rect 870 748 874 751
rect 734 738 738 742
rect 750 738 754 742
rect 750 718 754 722
rect 710 678 714 682
rect 678 668 682 672
rect 702 658 706 662
rect 750 658 754 662
rect 654 648 658 652
rect 686 648 690 652
rect 734 648 738 652
rect 750 648 754 652
rect 654 628 658 632
rect 670 628 674 632
rect 654 598 658 602
rect 654 578 658 582
rect 662 568 666 572
rect 638 558 642 562
rect 406 518 410 522
rect 510 508 514 512
rect 486 488 490 492
rect 574 528 578 532
rect 542 508 546 512
rect 558 508 562 512
rect 590 508 594 512
rect 558 488 562 492
rect 390 478 394 482
rect 534 478 538 482
rect 630 478 634 482
rect 742 628 746 632
rect 742 608 746 612
rect 758 598 762 602
rect 694 558 698 562
rect 734 558 738 562
rect 742 548 746 552
rect 670 488 674 492
rect 366 468 370 472
rect 478 468 482 472
rect 566 468 570 472
rect 350 438 354 442
rect 350 428 354 432
rect 286 398 290 402
rect 326 398 330 402
rect 406 428 410 432
rect 374 418 378 422
rect 326 378 330 382
rect 310 368 314 372
rect 350 368 354 372
rect 254 348 258 352
rect 198 338 202 342
rect 238 338 242 342
rect 262 338 266 342
rect 270 338 274 342
rect 174 328 178 332
rect 118 268 122 272
rect 166 308 170 312
rect 214 308 218 312
rect 206 298 210 302
rect 486 408 490 412
rect 374 398 378 402
rect 406 388 410 392
rect 462 388 466 392
rect 422 368 426 372
rect 318 348 322 352
rect 342 348 346 352
rect 310 338 314 342
rect 406 338 410 342
rect 302 298 306 302
rect 310 298 314 302
rect 294 288 298 292
rect 158 278 162 282
rect 214 278 218 282
rect 286 278 290 282
rect 206 268 210 272
rect 294 268 298 272
rect 382 328 386 332
rect 406 318 410 322
rect 326 308 330 312
rect 382 298 386 302
rect 406 298 410 302
rect 318 278 322 282
rect 374 278 378 282
rect 310 268 314 272
rect 14 118 18 122
rect 22 118 26 122
rect 126 258 130 262
rect 158 258 162 262
rect 246 258 250 262
rect 270 258 274 262
rect 302 258 306 262
rect 190 248 194 252
rect 198 248 202 252
rect 310 248 314 252
rect 126 238 130 242
rect 150 218 154 222
rect 70 198 74 202
rect 94 188 98 192
rect 150 188 154 192
rect 86 148 90 152
rect 134 138 138 142
rect 54 118 58 122
rect 94 78 98 82
rect 118 68 122 72
rect 238 238 242 242
rect 246 238 250 242
rect 278 238 282 242
rect 214 228 218 232
rect 230 228 234 232
rect 222 198 226 202
rect 206 178 210 182
rect 238 178 242 182
rect 166 158 170 162
rect 182 68 186 72
rect 390 288 394 292
rect 350 258 354 262
rect 374 248 378 252
rect 342 238 346 242
rect 358 238 362 242
rect 334 228 338 232
rect 318 218 322 222
rect 262 178 266 182
rect 222 168 226 172
rect 222 158 226 162
rect 238 158 242 162
rect 230 148 234 152
rect 310 208 314 212
rect 294 168 298 172
rect 222 88 226 92
rect 230 88 234 92
rect 262 78 266 82
rect 278 68 282 72
rect 358 198 362 202
rect 366 188 370 192
rect 406 258 410 262
rect 478 358 482 362
rect 498 403 502 407
rect 505 403 509 407
rect 622 458 626 462
rect 558 378 562 382
rect 582 448 586 452
rect 606 448 610 452
rect 638 448 642 452
rect 646 448 650 452
rect 590 438 594 442
rect 606 418 610 422
rect 622 418 626 422
rect 590 388 594 392
rect 606 388 610 392
rect 590 378 594 382
rect 638 378 642 382
rect 622 368 626 372
rect 470 348 474 352
rect 558 348 562 352
rect 566 348 570 352
rect 574 348 578 352
rect 438 328 442 332
rect 470 328 474 332
rect 454 288 458 292
rect 430 258 434 262
rect 454 258 458 262
rect 422 208 426 212
rect 462 198 466 202
rect 390 178 394 182
rect 390 168 394 172
rect 350 158 354 162
rect 422 158 426 162
rect 326 148 330 152
rect 342 148 346 152
rect 366 148 370 152
rect 406 148 410 152
rect 358 88 362 92
rect 542 308 546 312
rect 486 298 490 302
rect 502 288 506 292
rect 478 278 482 282
rect 494 278 498 282
rect 526 278 530 282
rect 542 278 546 282
rect 478 258 482 262
rect 494 248 498 252
rect 498 203 502 207
rect 505 203 509 207
rect 510 168 514 172
rect 566 308 570 312
rect 550 258 554 262
rect 558 238 562 242
rect 542 218 546 222
rect 534 198 538 202
rect 558 178 562 182
rect 590 328 594 332
rect 614 328 618 332
rect 598 318 602 322
rect 582 288 586 292
rect 590 278 594 282
rect 598 258 602 262
rect 622 278 626 282
rect 646 338 650 342
rect 678 458 682 462
rect 710 488 714 492
rect 726 478 730 482
rect 726 468 730 472
rect 742 468 746 472
rect 790 698 794 702
rect 782 568 786 572
rect 782 558 786 562
rect 830 688 834 692
rect 1166 928 1170 932
rect 1190 908 1194 912
rect 1214 898 1218 902
rect 1166 878 1170 882
rect 1182 878 1186 882
rect 1254 928 1258 932
rect 1294 938 1298 942
rect 1286 918 1290 922
rect 1278 898 1282 902
rect 1254 888 1258 892
rect 1270 888 1274 892
rect 1286 878 1290 882
rect 1350 1068 1354 1072
rect 1374 1168 1378 1172
rect 1398 1308 1402 1312
rect 1414 1298 1418 1302
rect 1422 1298 1426 1302
rect 1406 1278 1410 1282
rect 1398 1268 1402 1272
rect 1398 1248 1402 1252
rect 1522 1403 1526 1407
rect 1529 1403 1533 1407
rect 1470 1368 1474 1372
rect 1494 1368 1498 1372
rect 1550 1368 1554 1372
rect 1462 1338 1466 1342
rect 1462 1328 1466 1332
rect 1446 1308 1450 1312
rect 1454 1298 1458 1302
rect 1462 1268 1466 1272
rect 1430 1188 1434 1192
rect 1446 1238 1450 1242
rect 1542 1358 1546 1362
rect 1502 1348 1506 1352
rect 1494 1338 1498 1342
rect 1542 1338 1546 1342
rect 1486 1288 1490 1292
rect 1470 1248 1474 1252
rect 1486 1248 1490 1252
rect 1462 1228 1466 1232
rect 1438 1178 1442 1182
rect 1478 1228 1482 1232
rect 1518 1318 1522 1322
rect 1534 1258 1538 1262
rect 1510 1248 1514 1252
rect 1526 1238 1530 1242
rect 1502 1208 1506 1212
rect 1494 1198 1498 1202
rect 1478 1168 1482 1172
rect 1398 1158 1402 1162
rect 1438 1158 1442 1162
rect 1454 1158 1458 1162
rect 1494 1158 1498 1162
rect 1406 1148 1410 1152
rect 1382 1138 1386 1142
rect 1414 1138 1418 1142
rect 1430 1138 1434 1142
rect 1522 1203 1526 1207
rect 1529 1203 1533 1207
rect 1542 1158 1546 1162
rect 1574 1438 1578 1442
rect 1622 1448 1626 1452
rect 2062 1878 2066 1882
rect 1982 1858 1986 1862
rect 1998 1858 2002 1862
rect 2014 1858 2018 1862
rect 2278 2128 2282 2132
rect 2366 2128 2370 2132
rect 2246 2078 2250 2082
rect 2326 2118 2330 2122
rect 2294 2088 2298 2092
rect 2350 2088 2354 2092
rect 2342 2078 2346 2082
rect 2294 2068 2298 2072
rect 2326 2068 2330 2072
rect 2278 2058 2282 2062
rect 2246 2028 2250 2032
rect 2278 2028 2282 2032
rect 2286 1998 2290 2002
rect 2294 1948 2298 1952
rect 2382 2118 2386 2122
rect 2446 2118 2450 2122
rect 2318 2058 2322 2062
rect 2310 1978 2314 1982
rect 2278 1938 2282 1942
rect 2326 2028 2330 2032
rect 2350 2028 2354 2032
rect 2342 1978 2346 1982
rect 2350 1978 2354 1982
rect 2318 1938 2322 1942
rect 2310 1888 2314 1892
rect 2182 1878 2186 1882
rect 2206 1878 2210 1882
rect 2302 1878 2306 1882
rect 2342 1878 2346 1882
rect 2062 1868 2066 1872
rect 2102 1868 2106 1872
rect 2078 1858 2082 1862
rect 2118 1858 2122 1862
rect 2070 1758 2074 1762
rect 2006 1748 2010 1752
rect 2054 1748 2058 1752
rect 1966 1738 1970 1742
rect 2230 1868 2234 1872
rect 2142 1858 2146 1862
rect 2214 1858 2218 1862
rect 2182 1848 2186 1852
rect 2166 1838 2170 1842
rect 2174 1838 2178 1842
rect 2230 1838 2234 1842
rect 2294 1858 2298 1862
rect 2478 2128 2482 2132
rect 2390 2088 2394 2092
rect 2462 2088 2466 2092
rect 2534 2108 2538 2112
rect 2494 2088 2498 2092
rect 2422 2068 2426 2072
rect 2470 2068 2474 2072
rect 2478 2068 2482 2072
rect 2526 2068 2530 2072
rect 2414 2058 2418 2062
rect 2438 2058 2442 2062
rect 2478 2058 2482 2062
rect 2518 2058 2522 2062
rect 2406 2048 2410 2052
rect 2494 2048 2498 2052
rect 2438 2028 2442 2032
rect 2478 1988 2482 1992
rect 2454 1958 2458 1962
rect 2470 1958 2474 1962
rect 2382 1948 2386 1952
rect 2422 1948 2426 1952
rect 2398 1928 2402 1932
rect 2422 1928 2426 1932
rect 2422 1918 2426 1922
rect 2398 1908 2402 1912
rect 2414 1878 2418 1882
rect 2462 1928 2466 1932
rect 2454 1908 2458 1912
rect 2470 1908 2474 1912
rect 2494 1948 2498 1952
rect 2494 1908 2498 1912
rect 2526 2048 2530 2052
rect 2582 2098 2586 2102
rect 2742 2098 2746 2102
rect 2678 2088 2682 2092
rect 2606 2078 2610 2082
rect 2702 2078 2706 2082
rect 2734 2078 2738 2082
rect 2758 2208 2762 2212
rect 2950 2658 2954 2662
rect 2990 2728 2994 2732
rect 2990 2708 2994 2712
rect 2982 2688 2986 2692
rect 2958 2648 2962 2652
rect 2934 2638 2938 2642
rect 2950 2628 2954 2632
rect 2958 2598 2962 2602
rect 2926 2568 2930 2572
rect 2926 2538 2930 2542
rect 3006 2778 3010 2782
rect 3006 2768 3010 2772
rect 3030 2768 3034 2772
rect 3014 2748 3018 2752
rect 3006 2648 3010 2652
rect 2982 2578 2986 2582
rect 2966 2548 2970 2552
rect 2974 2528 2978 2532
rect 2958 2518 2962 2522
rect 2934 2508 2938 2512
rect 2926 2498 2930 2502
rect 2926 2488 2930 2492
rect 2958 2508 2962 2512
rect 3070 2928 3074 2932
rect 3050 2903 3054 2907
rect 3057 2903 3061 2907
rect 3078 2898 3082 2902
rect 3086 2878 3090 2882
rect 3054 2858 3058 2862
rect 3094 2848 3098 2852
rect 3078 2768 3082 2772
rect 3062 2748 3066 2752
rect 3050 2703 3054 2707
rect 3057 2703 3061 2707
rect 3030 2678 3034 2682
rect 3158 2928 3162 2932
rect 3142 2858 3146 2862
rect 3190 2928 3194 2932
rect 3190 2908 3194 2912
rect 3198 2898 3202 2902
rect 3190 2868 3194 2872
rect 3158 2768 3162 2772
rect 3142 2758 3146 2762
rect 3134 2748 3138 2752
rect 3102 2718 3106 2722
rect 3094 2698 3098 2702
rect 3094 2688 3098 2692
rect 3094 2658 3098 2662
rect 3006 2568 3010 2572
rect 3022 2568 3026 2572
rect 2990 2538 2994 2542
rect 2974 2468 2978 2472
rect 2982 2468 2986 2472
rect 2974 2458 2978 2462
rect 2934 2408 2938 2412
rect 2918 2398 2922 2402
rect 2950 2398 2954 2402
rect 2918 2358 2922 2362
rect 2998 2378 3002 2382
rect 2974 2358 2978 2362
rect 2926 2348 2930 2352
rect 2958 2348 2962 2352
rect 2982 2348 2986 2352
rect 2918 2328 2922 2332
rect 3078 2558 3082 2562
rect 3222 2908 3226 2912
rect 3214 2898 3218 2902
rect 3206 2828 3210 2832
rect 3310 3048 3314 3052
rect 3294 2938 3298 2942
rect 3238 2928 3242 2932
rect 3350 3088 3354 3092
rect 3382 3068 3386 3072
rect 3334 2968 3338 2972
rect 3406 3278 3410 3282
rect 3422 3278 3426 3282
rect 3414 3258 3418 3262
rect 3570 3603 3574 3607
rect 3577 3603 3581 3607
rect 3718 3948 3722 3952
rect 3742 3938 3746 3942
rect 3710 3908 3714 3912
rect 3758 3968 3762 3972
rect 3830 4028 3834 4032
rect 3814 4018 3818 4022
rect 3806 3998 3810 4002
rect 3798 3978 3802 3982
rect 3806 3958 3810 3962
rect 3782 3938 3786 3942
rect 3774 3928 3778 3932
rect 3862 4018 3866 4022
rect 3838 3978 3842 3982
rect 3846 3958 3850 3962
rect 3854 3948 3858 3952
rect 3902 4038 3906 4042
rect 3990 4098 3994 4102
rect 3982 4088 3986 4092
rect 4082 4303 4086 4307
rect 4089 4303 4093 4307
rect 4134 4308 4138 4312
rect 4102 4298 4106 4302
rect 4134 4298 4138 4302
rect 4150 4298 4154 4302
rect 4094 4288 4098 4292
rect 4126 4288 4130 4292
rect 4102 4278 4106 4282
rect 4094 4258 4098 4262
rect 4110 4258 4114 4262
rect 4126 4258 4130 4262
rect 4070 4248 4074 4252
rect 4078 4228 4082 4232
rect 4038 4178 4042 4182
rect 4038 4158 4042 4162
rect 4062 4158 4066 4162
rect 4030 4118 4034 4122
rect 4054 4118 4058 4122
rect 3998 4068 4002 4072
rect 4006 4068 4010 4072
rect 4038 4108 4042 4112
rect 3974 4058 3978 4062
rect 3934 4038 3938 4042
rect 4014 4048 4018 4052
rect 4030 4048 4034 4052
rect 3958 4038 3962 4042
rect 3918 4028 3922 4032
rect 3950 4028 3954 4032
rect 3926 4018 3930 4022
rect 3966 4018 3970 4022
rect 3990 4018 3994 4022
rect 3958 4008 3962 4012
rect 3942 3968 3946 3972
rect 3878 3958 3882 3962
rect 3926 3958 3930 3962
rect 3878 3948 3882 3952
rect 3894 3948 3898 3952
rect 3902 3948 3906 3952
rect 3822 3938 3826 3942
rect 3838 3938 3842 3942
rect 3854 3938 3858 3942
rect 3774 3898 3778 3902
rect 3798 3898 3802 3902
rect 3678 3878 3682 3882
rect 3758 3878 3762 3882
rect 3702 3868 3706 3872
rect 3742 3866 3746 3870
rect 3694 3858 3698 3862
rect 3718 3858 3722 3862
rect 3678 3848 3682 3852
rect 3670 3778 3674 3782
rect 3926 3938 3930 3942
rect 3878 3928 3882 3932
rect 3894 3928 3898 3932
rect 3918 3928 3922 3932
rect 3822 3918 3826 3922
rect 3830 3918 3834 3922
rect 3910 3908 3914 3912
rect 3878 3888 3882 3892
rect 3950 3948 3954 3952
rect 3966 3978 3970 3982
rect 3982 3968 3986 3972
rect 4030 3998 4034 4002
rect 4006 3988 4010 3992
rect 4022 3968 4026 3972
rect 3982 3948 3986 3952
rect 3990 3948 3994 3952
rect 3958 3928 3962 3932
rect 3974 3928 3978 3932
rect 3974 3898 3978 3902
rect 3782 3878 3786 3882
rect 3846 3878 3850 3882
rect 3918 3878 3922 3882
rect 3934 3878 3938 3882
rect 3782 3868 3786 3872
rect 3926 3868 3930 3872
rect 3758 3848 3762 3852
rect 3630 3748 3634 3752
rect 3742 3748 3746 3752
rect 3734 3718 3738 3722
rect 3766 3828 3770 3832
rect 3822 3858 3826 3862
rect 3806 3828 3810 3832
rect 3806 3758 3810 3762
rect 4046 4068 4050 4072
rect 4082 4103 4086 4107
rect 4089 4103 4093 4107
rect 4118 4188 4122 4192
rect 4110 4158 4114 4162
rect 4102 4098 4106 4102
rect 4110 4078 4114 4082
rect 4078 4058 4082 4062
rect 4070 3998 4074 4002
rect 4062 3988 4066 3992
rect 4094 4048 4098 4052
rect 4150 4258 4154 4262
rect 4158 4258 4162 4262
rect 4166 4248 4170 4252
rect 4278 4368 4282 4372
rect 4238 4348 4242 4352
rect 4286 4348 4290 4352
rect 4198 4318 4202 4322
rect 4238 4298 4242 4302
rect 4246 4298 4250 4302
rect 4238 4288 4242 4292
rect 4278 4338 4282 4342
rect 4270 4318 4274 4322
rect 4262 4278 4266 4282
rect 4302 4338 4306 4342
rect 4326 4358 4330 4362
rect 4342 4358 4346 4362
rect 4430 4398 4434 4402
rect 4382 4388 4386 4392
rect 4502 4378 4506 4382
rect 4414 4368 4418 4372
rect 4358 4358 4362 4362
rect 4446 4358 4450 4362
rect 4390 4348 4394 4352
rect 4478 4348 4482 4352
rect 4486 4348 4490 4352
rect 4326 4338 4330 4342
rect 4358 4338 4362 4342
rect 4310 4288 4314 4292
rect 4358 4288 4362 4292
rect 4374 4288 4378 4292
rect 4294 4268 4298 4272
rect 4206 4258 4210 4262
rect 4254 4258 4258 4262
rect 4190 4238 4194 4242
rect 4142 4188 4146 4192
rect 4174 4178 4178 4182
rect 4134 4168 4138 4172
rect 4142 4158 4146 4162
rect 4158 4158 4162 4162
rect 4182 4168 4186 4172
rect 4238 4248 4242 4252
rect 4230 4178 4234 4182
rect 4286 4258 4290 4262
rect 4270 4248 4274 4252
rect 4262 4208 4266 4212
rect 4302 4248 4306 4252
rect 4302 4228 4306 4232
rect 4302 4208 4306 4212
rect 4246 4198 4250 4202
rect 4278 4198 4282 4202
rect 4294 4198 4298 4202
rect 4206 4158 4210 4162
rect 4198 4148 4202 4152
rect 4214 4148 4218 4152
rect 4126 4118 4130 4122
rect 4174 4118 4178 4122
rect 4134 4108 4138 4112
rect 4150 4098 4154 4102
rect 4126 4088 4130 4092
rect 4126 4078 4130 4082
rect 4182 4108 4186 4112
rect 4206 4108 4210 4112
rect 4222 4108 4226 4112
rect 4214 4098 4218 4102
rect 4166 4068 4170 4072
rect 4198 4068 4202 4072
rect 4134 4058 4138 4062
rect 4142 4058 4146 4062
rect 4118 4018 4122 4022
rect 4158 4018 4162 4022
rect 4150 4008 4154 4012
rect 4142 3958 4146 3962
rect 4054 3948 4058 3952
rect 4126 3948 4130 3952
rect 4046 3938 4050 3942
rect 4038 3918 4042 3922
rect 4006 3898 4010 3902
rect 3998 3878 4002 3882
rect 3886 3858 3890 3862
rect 3918 3858 3922 3862
rect 3942 3858 3946 3862
rect 3982 3858 3986 3862
rect 3838 3828 3842 3832
rect 3838 3758 3842 3762
rect 4102 3908 4106 3912
rect 4082 3903 4086 3907
rect 4089 3903 4093 3907
rect 4062 3888 4066 3892
rect 4102 3888 4106 3892
rect 4038 3878 4042 3882
rect 4078 3878 4082 3882
rect 4022 3868 4026 3872
rect 3862 3848 3866 3852
rect 3886 3848 3890 3852
rect 3862 3838 3866 3842
rect 4030 3838 4034 3842
rect 3982 3828 3986 3832
rect 3926 3808 3930 3812
rect 3966 3788 3970 3792
rect 4006 3788 4010 3792
rect 3854 3768 3858 3772
rect 3934 3768 3938 3772
rect 3926 3758 3930 3762
rect 3974 3778 3978 3782
rect 4054 3868 4058 3872
rect 4062 3858 4066 3862
rect 4070 3848 4074 3852
rect 4118 3848 4122 3852
rect 4166 3978 4170 3982
rect 4238 4098 4242 4102
rect 4238 4068 4242 4072
rect 4214 4058 4218 4062
rect 4254 4168 4258 4172
rect 4286 4168 4290 4172
rect 4262 4158 4266 4162
rect 4310 4158 4314 4162
rect 4254 4138 4258 4142
rect 4270 4138 4274 4142
rect 4262 4128 4266 4132
rect 4262 4068 4266 4072
rect 4294 4128 4298 4132
rect 4334 4258 4338 4262
rect 4350 4248 4354 4252
rect 4398 4338 4402 4342
rect 4414 4338 4418 4342
rect 4390 4328 4394 4332
rect 4406 4328 4410 4332
rect 4430 4328 4434 4332
rect 4390 4318 4394 4322
rect 4422 4298 4426 4302
rect 4406 4288 4410 4292
rect 4454 4338 4458 4342
rect 4478 4308 4482 4312
rect 4486 4308 4490 4312
rect 4446 4298 4450 4302
rect 4566 4368 4570 4372
rect 4510 4348 4514 4352
rect 4534 4348 4538 4352
rect 4582 4338 4586 4342
rect 4438 4278 4442 4282
rect 4462 4278 4466 4282
rect 4502 4278 4506 4282
rect 4494 4268 4498 4272
rect 4470 4258 4474 4262
rect 4382 4248 4386 4252
rect 4358 4238 4362 4242
rect 4326 4228 4330 4232
rect 4406 4228 4410 4232
rect 4398 4208 4402 4212
rect 4390 4198 4394 4202
rect 4334 4178 4338 4182
rect 4462 4248 4466 4252
rect 4478 4248 4482 4252
rect 4518 4288 4522 4292
rect 4550 4318 4554 4322
rect 4534 4308 4538 4312
rect 4526 4278 4530 4282
rect 4526 4268 4530 4272
rect 4566 4268 4570 4272
rect 4534 4258 4538 4262
rect 4510 4238 4514 4242
rect 4486 4228 4490 4232
rect 4454 4218 4458 4222
rect 4438 4208 4442 4212
rect 4430 4178 4434 4182
rect 4406 4168 4410 4172
rect 4366 4158 4370 4162
rect 4382 4158 4386 4162
rect 4398 4158 4402 4162
rect 4358 4148 4362 4152
rect 4446 4168 4450 4172
rect 4518 4208 4522 4212
rect 4502 4188 4506 4192
rect 4510 4158 4514 4162
rect 4542 4208 4546 4212
rect 4574 4228 4578 4232
rect 4438 4148 4442 4152
rect 4446 4148 4450 4152
rect 4470 4148 4474 4152
rect 4478 4148 4482 4152
rect 4526 4148 4530 4152
rect 4318 4138 4322 4142
rect 4326 4138 4330 4142
rect 4382 4138 4386 4142
rect 4422 4138 4426 4142
rect 4430 4138 4434 4142
rect 4334 4128 4338 4132
rect 4366 4128 4370 4132
rect 4302 4108 4306 4112
rect 4318 4098 4322 4102
rect 4286 4068 4290 4072
rect 4318 4068 4322 4072
rect 4254 4058 4258 4062
rect 4270 4058 4274 4062
rect 4294 4058 4298 4062
rect 4318 4058 4322 4062
rect 4222 4028 4226 4032
rect 4262 4048 4266 4052
rect 4286 4048 4290 4052
rect 4318 4048 4322 4052
rect 4374 4108 4378 4112
rect 4438 4108 4442 4112
rect 4366 4068 4370 4072
rect 4270 4038 4274 4042
rect 4246 3968 4250 3972
rect 4246 3958 4250 3962
rect 4350 3978 4354 3982
rect 4358 3968 4362 3972
rect 4454 4138 4458 4142
rect 4478 4118 4482 4122
rect 4486 4118 4490 4122
rect 4510 4098 4514 4102
rect 4542 4098 4546 4102
rect 4390 4088 4394 4092
rect 4422 4088 4426 4092
rect 4470 4088 4474 4092
rect 4534 4088 4538 4092
rect 4398 4078 4402 4082
rect 4430 4078 4434 4082
rect 4478 4078 4482 4082
rect 4510 4078 4514 4082
rect 4542 4078 4546 4082
rect 4502 4068 4506 4072
rect 4454 4058 4458 4062
rect 4510 4058 4514 4062
rect 4558 4148 4562 4152
rect 4590 4218 4594 4222
rect 4598 4158 4602 4162
rect 4558 4118 4562 4122
rect 4558 4108 4562 4112
rect 4590 4108 4594 4112
rect 4550 4068 4554 4072
rect 4566 4068 4570 4072
rect 4406 4048 4410 4052
rect 4422 4048 4426 4052
rect 4470 4048 4474 4052
rect 4494 4048 4498 4052
rect 4510 4048 4514 4052
rect 4526 4048 4530 4052
rect 4446 4038 4450 4042
rect 4390 3998 4394 4002
rect 4190 3948 4194 3952
rect 4230 3948 4234 3952
rect 4270 3948 4274 3952
rect 4366 3948 4370 3952
rect 4182 3938 4186 3942
rect 4222 3938 4226 3942
rect 4230 3938 4234 3942
rect 4246 3938 4250 3942
rect 4302 3938 4306 3942
rect 4190 3928 4194 3932
rect 4174 3908 4178 3912
rect 4142 3868 4146 3872
rect 4158 3858 4162 3862
rect 4174 3838 4178 3842
rect 4134 3828 4138 3832
rect 4054 3788 4058 3792
rect 4134 3768 4138 3772
rect 4102 3758 4106 3762
rect 4214 3908 4218 3912
rect 4222 3898 4226 3902
rect 4238 3928 4242 3932
rect 4294 3928 4298 3932
rect 4350 3928 4354 3932
rect 4238 3918 4242 3922
rect 4302 3918 4306 3922
rect 4206 3868 4210 3872
rect 4222 3868 4226 3872
rect 4190 3828 4194 3832
rect 4198 3808 4202 3812
rect 4270 3878 4274 3882
rect 4310 3878 4314 3882
rect 4318 3878 4322 3882
rect 4350 3898 4354 3902
rect 4262 3868 4266 3872
rect 4302 3868 4306 3872
rect 4262 3858 4266 3862
rect 4286 3858 4290 3862
rect 4214 3848 4218 3852
rect 4230 3848 4234 3852
rect 4246 3828 4250 3832
rect 4230 3808 4234 3812
rect 4198 3788 4202 3792
rect 4206 3788 4210 3792
rect 4254 3768 4258 3772
rect 4294 3768 4298 3772
rect 3830 3748 3834 3752
rect 3806 3738 3810 3742
rect 3822 3738 3826 3742
rect 3774 3728 3778 3732
rect 3798 3728 3802 3732
rect 3822 3728 3826 3732
rect 3838 3728 3842 3732
rect 3878 3728 3882 3732
rect 3782 3718 3786 3722
rect 3710 3708 3714 3712
rect 3758 3708 3762 3712
rect 3782 3708 3786 3712
rect 3814 3708 3818 3712
rect 3734 3678 3738 3682
rect 3630 3668 3634 3672
rect 3662 3668 3666 3672
rect 3726 3658 3730 3662
rect 3694 3608 3698 3612
rect 3462 3598 3466 3602
rect 3590 3598 3594 3602
rect 3510 3588 3514 3592
rect 3614 3578 3618 3582
rect 3542 3558 3546 3562
rect 3494 3538 3498 3542
rect 3510 3538 3514 3542
rect 3574 3538 3578 3542
rect 3462 3508 3466 3512
rect 3686 3538 3690 3542
rect 3654 3528 3658 3532
rect 3518 3498 3522 3502
rect 3518 3478 3522 3482
rect 3622 3478 3626 3482
rect 3470 3468 3474 3472
rect 3494 3468 3498 3472
rect 3510 3468 3514 3472
rect 3574 3468 3578 3472
rect 3654 3468 3658 3472
rect 3462 3458 3466 3462
rect 3478 3458 3482 3462
rect 3606 3458 3610 3462
rect 3526 3438 3530 3442
rect 3598 3438 3602 3442
rect 3606 3438 3610 3442
rect 3534 3408 3538 3412
rect 3570 3403 3574 3407
rect 3577 3403 3581 3407
rect 3462 3388 3466 3392
rect 3470 3378 3474 3382
rect 3502 3378 3506 3382
rect 3614 3378 3618 3382
rect 3638 3378 3642 3382
rect 3462 3358 3466 3362
rect 3478 3358 3482 3362
rect 3526 3348 3530 3352
rect 3550 3348 3554 3352
rect 3646 3348 3650 3352
rect 3486 3338 3490 3342
rect 3510 3338 3514 3342
rect 3534 3338 3538 3342
rect 3558 3338 3562 3342
rect 3582 3338 3586 3342
rect 3622 3338 3626 3342
rect 3646 3338 3650 3342
rect 3454 3328 3458 3332
rect 3510 3328 3514 3332
rect 3446 3228 3450 3232
rect 3454 3228 3458 3232
rect 3502 3248 3506 3252
rect 3518 3308 3522 3312
rect 3526 3278 3530 3282
rect 3558 3238 3562 3242
rect 3606 3248 3610 3252
rect 3518 3218 3522 3222
rect 3566 3218 3570 3222
rect 3570 3203 3574 3207
rect 3577 3203 3581 3207
rect 3574 3158 3578 3162
rect 3558 3148 3562 3152
rect 3430 3138 3434 3142
rect 3494 3138 3498 3142
rect 3502 3118 3506 3122
rect 3470 3108 3474 3112
rect 3462 3068 3466 3072
rect 3390 3028 3394 3032
rect 3510 3078 3514 3082
rect 3646 3298 3650 3302
rect 3670 3358 3674 3362
rect 3686 3348 3690 3352
rect 3694 3338 3698 3342
rect 3814 3668 3818 3672
rect 3742 3658 3746 3662
rect 3726 3588 3730 3592
rect 3726 3568 3730 3572
rect 3734 3568 3738 3572
rect 3742 3558 3746 3562
rect 3798 3568 3802 3572
rect 3750 3548 3754 3552
rect 3726 3488 3730 3492
rect 3806 3538 3810 3542
rect 3742 3478 3746 3482
rect 3742 3458 3746 3462
rect 3766 3458 3770 3462
rect 3782 3458 3786 3462
rect 3726 3448 3730 3452
rect 3750 3448 3754 3452
rect 3782 3448 3786 3452
rect 3734 3388 3738 3392
rect 3742 3358 3746 3362
rect 3726 3348 3730 3352
rect 3774 3338 3778 3342
rect 3670 3328 3674 3332
rect 3702 3328 3706 3332
rect 3750 3318 3754 3322
rect 3702 3288 3706 3292
rect 3662 3278 3666 3282
rect 3670 3278 3674 3282
rect 3702 3258 3706 3262
rect 3670 3238 3674 3242
rect 3662 3218 3666 3222
rect 3910 3748 3914 3752
rect 4022 3748 4026 3752
rect 4046 3748 4050 3752
rect 4078 3748 4082 3752
rect 3894 3738 3898 3742
rect 3886 3718 3890 3722
rect 3950 3738 3954 3742
rect 3982 3738 3986 3742
rect 4014 3738 4018 3742
rect 4086 3738 4090 3742
rect 3958 3728 3962 3732
rect 3958 3688 3962 3692
rect 3926 3668 3930 3672
rect 3910 3658 3914 3662
rect 3902 3588 3906 3592
rect 3878 3568 3882 3572
rect 3886 3558 3890 3562
rect 3998 3728 4002 3732
rect 4038 3728 4042 3732
rect 3998 3678 4002 3682
rect 4030 3668 4034 3672
rect 4110 3708 4114 3712
rect 4126 3708 4130 3712
rect 4082 3703 4086 3707
rect 4089 3703 4093 3707
rect 4022 3658 4026 3662
rect 4038 3658 4042 3662
rect 4198 3738 4202 3742
rect 4158 3708 4162 3712
rect 4118 3678 4122 3682
rect 4134 3678 4138 3682
rect 4166 3678 4170 3682
rect 4126 3668 4130 3672
rect 4142 3668 4146 3672
rect 4174 3668 4178 3672
rect 4222 3668 4226 3672
rect 4094 3658 4098 3662
rect 4118 3658 4122 3662
rect 4150 3658 4154 3662
rect 4182 3658 4186 3662
rect 4214 3658 4218 3662
rect 4022 3648 4026 3652
rect 4054 3648 4058 3652
rect 4070 3648 4074 3652
rect 4078 3648 4082 3652
rect 4150 3648 4154 3652
rect 4182 3648 4186 3652
rect 4030 3638 4034 3642
rect 3990 3628 3994 3632
rect 4022 3618 4026 3622
rect 4014 3578 4018 3582
rect 3982 3558 3986 3562
rect 3926 3547 3930 3551
rect 3998 3548 4002 3552
rect 3950 3538 3954 3542
rect 3862 3528 3866 3532
rect 3862 3478 3866 3482
rect 3862 3458 3866 3462
rect 3846 3368 3850 3372
rect 3886 3458 3890 3462
rect 3950 3459 3954 3463
rect 3886 3438 3890 3442
rect 4006 3468 4010 3472
rect 3990 3428 3994 3432
rect 3886 3378 3890 3382
rect 4038 3448 4042 3452
rect 3830 3348 3834 3352
rect 3886 3348 3890 3352
rect 4214 3628 4218 3632
rect 4110 3548 4114 3552
rect 4082 3503 4086 3507
rect 4089 3503 4093 3507
rect 4246 3738 4250 3742
rect 4262 3758 4266 3762
rect 4270 3748 4274 3752
rect 4310 3748 4314 3752
rect 4262 3738 4266 3742
rect 4302 3738 4306 3742
rect 4286 3728 4290 3732
rect 4254 3688 4258 3692
rect 4262 3678 4266 3682
rect 4310 3718 4314 3722
rect 4326 3868 4330 3872
rect 4334 3858 4338 3862
rect 4430 3988 4434 3992
rect 4494 3978 4498 3982
rect 4462 3968 4466 3972
rect 4446 3958 4450 3962
rect 4470 3958 4474 3962
rect 4406 3948 4410 3952
rect 4438 3948 4442 3952
rect 4470 3948 4474 3952
rect 4486 3948 4490 3952
rect 4390 3938 4394 3942
rect 4414 3938 4418 3942
rect 4382 3928 4386 3932
rect 4390 3928 4394 3932
rect 4398 3918 4402 3922
rect 4374 3878 4378 3882
rect 4350 3858 4354 3862
rect 4366 3858 4370 3862
rect 4382 3858 4386 3862
rect 4374 3848 4378 3852
rect 4342 3808 4346 3812
rect 4326 3758 4330 3762
rect 4334 3758 4338 3762
rect 4366 3758 4370 3762
rect 4406 3838 4410 3842
rect 4398 3758 4402 3762
rect 4326 3738 4330 3742
rect 4358 3738 4362 3742
rect 4390 3738 4394 3742
rect 4398 3728 4402 3732
rect 4398 3718 4402 3722
rect 4382 3688 4386 3692
rect 4454 3918 4458 3922
rect 4430 3888 4434 3892
rect 4446 3888 4450 3892
rect 4486 3888 4490 3892
rect 4470 3868 4474 3872
rect 4430 3858 4434 3862
rect 4446 3858 4450 3862
rect 4454 3848 4458 3852
rect 4502 3928 4506 3932
rect 4534 4038 4538 4042
rect 4542 4028 4546 4032
rect 4518 3978 4522 3982
rect 4542 3978 4546 3982
rect 4526 3968 4530 3972
rect 4534 3958 4538 3962
rect 4550 3948 4554 3952
rect 4574 4058 4578 4062
rect 4566 4048 4570 4052
rect 4598 4038 4602 4042
rect 4598 4028 4602 4032
rect 4582 3958 4586 3962
rect 4590 3958 4594 3962
rect 4566 3948 4570 3952
rect 4582 3948 4586 3952
rect 4558 3928 4562 3932
rect 4518 3908 4522 3912
rect 4534 3878 4538 3882
rect 4502 3868 4506 3872
rect 4550 3868 4554 3872
rect 4462 3838 4466 3842
rect 4438 3828 4442 3832
rect 4486 3808 4490 3812
rect 4462 3798 4466 3802
rect 4478 3798 4482 3802
rect 4438 3768 4442 3772
rect 4422 3748 4426 3752
rect 4430 3738 4434 3742
rect 4446 3738 4450 3742
rect 4454 3728 4458 3732
rect 4526 3848 4530 3852
rect 4518 3758 4522 3762
rect 4542 3798 4546 3802
rect 4582 3798 4586 3802
rect 4510 3748 4514 3752
rect 4534 3748 4538 3752
rect 4486 3738 4490 3742
rect 4502 3738 4506 3742
rect 4462 3718 4466 3722
rect 4478 3698 4482 3702
rect 4510 3668 4514 3672
rect 4542 3728 4546 3732
rect 4550 3728 4554 3732
rect 4534 3718 4538 3722
rect 4566 3718 4570 3722
rect 4566 3668 4570 3672
rect 4278 3658 4282 3662
rect 4406 3658 4410 3662
rect 4310 3648 4314 3652
rect 4326 3638 4330 3642
rect 4374 3638 4378 3642
rect 4542 3648 4546 3652
rect 4518 3638 4522 3642
rect 4502 3628 4506 3632
rect 4230 3618 4234 3622
rect 4366 3618 4370 3622
rect 4446 3618 4450 3622
rect 4574 3618 4578 3622
rect 4270 3598 4274 3602
rect 4238 3548 4242 3552
rect 4326 3578 4330 3582
rect 4342 3558 4346 3562
rect 4318 3548 4322 3552
rect 4206 3538 4210 3542
rect 4222 3538 4226 3542
rect 4182 3508 4186 3512
rect 4126 3488 4130 3492
rect 4110 3478 4114 3482
rect 4230 3508 4234 3512
rect 4254 3508 4258 3512
rect 4222 3468 4226 3472
rect 4102 3448 4106 3452
rect 4102 3388 4106 3392
rect 3918 3338 3922 3342
rect 3798 3248 3802 3252
rect 3718 3218 3722 3222
rect 3766 3218 3770 3222
rect 3686 3168 3690 3172
rect 3774 3188 3778 3192
rect 3662 3148 3666 3152
rect 3678 3148 3682 3152
rect 3734 3148 3738 3152
rect 3750 3148 3754 3152
rect 3638 3128 3642 3132
rect 3750 3128 3754 3132
rect 3638 3108 3642 3112
rect 3606 3098 3610 3102
rect 3486 3068 3490 3072
rect 3542 3068 3546 3072
rect 3502 3058 3506 3062
rect 3518 3058 3522 3062
rect 3534 3058 3538 3062
rect 3630 3058 3634 3062
rect 3510 3048 3514 3052
rect 3614 3048 3618 3052
rect 3454 3038 3458 3042
rect 3470 3008 3474 3012
rect 3462 2988 3466 2992
rect 3358 2948 3362 2952
rect 3414 2948 3418 2952
rect 3318 2938 3322 2942
rect 3342 2938 3346 2942
rect 3390 2938 3394 2942
rect 3270 2918 3274 2922
rect 3246 2908 3250 2912
rect 3238 2898 3242 2902
rect 3254 2888 3258 2892
rect 3278 2898 3282 2902
rect 3262 2868 3266 2872
rect 3230 2848 3234 2852
rect 3246 2818 3250 2822
rect 3246 2808 3250 2812
rect 3326 2928 3330 2932
rect 3310 2908 3314 2912
rect 3342 2898 3346 2902
rect 3454 2898 3458 2902
rect 3334 2888 3338 2892
rect 3318 2878 3322 2882
rect 3350 2868 3354 2872
rect 3334 2858 3338 2862
rect 3262 2848 3266 2852
rect 3294 2848 3298 2852
rect 3302 2848 3306 2852
rect 3334 2798 3338 2802
rect 3246 2768 3250 2772
rect 3254 2768 3258 2772
rect 3294 2768 3298 2772
rect 3222 2758 3226 2762
rect 3190 2748 3194 2752
rect 3222 2748 3226 2752
rect 3238 2748 3242 2752
rect 3278 2738 3282 2742
rect 3174 2708 3178 2712
rect 3198 2698 3202 2702
rect 3182 2678 3186 2682
rect 3278 2678 3282 2682
rect 3198 2668 3202 2672
rect 3150 2658 3154 2662
rect 3150 2628 3154 2632
rect 3150 2568 3154 2572
rect 3050 2503 3054 2507
rect 3057 2503 3061 2507
rect 3078 2498 3082 2502
rect 3110 2478 3114 2482
rect 3062 2468 3066 2472
rect 3014 2358 3018 2362
rect 3054 2358 3058 2362
rect 3006 2338 3010 2342
rect 3038 2338 3042 2342
rect 3070 2338 3074 2342
rect 3006 2328 3010 2332
rect 2950 2318 2954 2322
rect 2982 2318 2986 2322
rect 2990 2298 2994 2302
rect 3050 2303 3054 2307
rect 3057 2303 3061 2307
rect 2998 2278 3002 2282
rect 3030 2278 3034 2282
rect 3006 2268 3010 2272
rect 3062 2268 3066 2272
rect 2918 2258 2922 2262
rect 2934 2258 2938 2262
rect 2958 2258 2962 2262
rect 2974 2258 2978 2262
rect 3022 2248 3026 2252
rect 3046 2248 3050 2252
rect 2942 2238 2946 2242
rect 2966 2238 2970 2242
rect 2910 2218 2914 2222
rect 3038 2198 3042 2202
rect 2910 2188 2914 2192
rect 2918 2188 2922 2192
rect 3006 2178 3010 2182
rect 2782 2158 2786 2162
rect 2806 2158 2810 2162
rect 2838 2158 2842 2162
rect 2926 2158 2930 2162
rect 2798 2138 2802 2142
rect 2838 2148 2842 2152
rect 2910 2138 2914 2142
rect 2782 2128 2786 2132
rect 2798 2128 2802 2132
rect 2822 2128 2826 2132
rect 2838 2128 2842 2132
rect 2758 2118 2762 2122
rect 2766 2118 2770 2122
rect 2782 2118 2786 2122
rect 2758 2098 2762 2102
rect 2590 2068 2594 2072
rect 2598 2068 2602 2072
rect 2622 2068 2626 2072
rect 2686 2068 2690 2072
rect 2710 2068 2714 2072
rect 2718 2068 2722 2072
rect 2758 2068 2762 2072
rect 2574 2048 2578 2052
rect 2598 2018 2602 2022
rect 2630 2058 2634 2062
rect 2646 2058 2650 2062
rect 2678 2058 2682 2062
rect 2758 2058 2762 2062
rect 2862 2088 2866 2092
rect 3062 2178 3066 2182
rect 3006 2148 3010 2152
rect 3022 2148 3026 2152
rect 3038 2148 3042 2152
rect 3118 2458 3122 2462
rect 3206 2648 3210 2652
rect 3222 2618 3226 2622
rect 3206 2568 3210 2572
rect 3214 2568 3218 2572
rect 3198 2558 3202 2562
rect 3198 2518 3202 2522
rect 3182 2478 3186 2482
rect 3174 2448 3178 2452
rect 3182 2428 3186 2432
rect 3222 2488 3226 2492
rect 3270 2648 3274 2652
rect 3278 2628 3282 2632
rect 3286 2558 3290 2562
rect 3262 2538 3266 2542
rect 3262 2508 3266 2512
rect 3254 2498 3258 2502
rect 3238 2488 3242 2492
rect 3310 2728 3314 2732
rect 3390 2858 3394 2862
rect 3398 2828 3402 2832
rect 3390 2818 3394 2822
rect 3358 2808 3362 2812
rect 3366 2758 3370 2762
rect 3414 2758 3418 2762
rect 3398 2738 3402 2742
rect 3570 3003 3574 3007
rect 3577 3003 3581 3007
rect 3686 3078 3690 3082
rect 3702 3068 3706 3072
rect 3822 3158 3826 3162
rect 3726 3058 3730 3062
rect 3686 3018 3690 3022
rect 3662 2978 3666 2982
rect 3646 2968 3650 2972
rect 3710 3008 3714 3012
rect 3742 2978 3746 2982
rect 3510 2948 3514 2952
rect 3630 2948 3634 2952
rect 3670 2948 3674 2952
rect 3702 2948 3706 2952
rect 3718 2948 3722 2952
rect 3534 2938 3538 2942
rect 3566 2938 3570 2942
rect 3710 2938 3714 2942
rect 3510 2918 3514 2922
rect 3502 2898 3506 2902
rect 3438 2858 3442 2862
rect 3526 2898 3530 2902
rect 3518 2868 3522 2872
rect 3502 2848 3506 2852
rect 3470 2758 3474 2762
rect 3454 2748 3458 2752
rect 3422 2728 3426 2732
rect 3502 2728 3506 2732
rect 3518 2728 3522 2732
rect 3342 2688 3346 2692
rect 3318 2588 3322 2592
rect 3358 2708 3362 2712
rect 3430 2718 3434 2722
rect 3558 2918 3562 2922
rect 3678 2908 3682 2912
rect 3606 2868 3610 2872
rect 3646 2868 3650 2872
rect 3570 2803 3574 2807
rect 3577 2803 3581 2807
rect 3670 2858 3674 2862
rect 3670 2828 3674 2832
rect 3646 2768 3650 2772
rect 3662 2748 3666 2752
rect 3702 2858 3706 2862
rect 3726 2858 3730 2862
rect 3726 2838 3730 2842
rect 3686 2748 3690 2752
rect 3582 2738 3586 2742
rect 3598 2738 3602 2742
rect 3566 2728 3570 2732
rect 3406 2668 3410 2672
rect 3446 2668 3450 2672
rect 3470 2668 3474 2672
rect 3534 2668 3538 2672
rect 3366 2648 3370 2652
rect 3390 2658 3394 2662
rect 3382 2648 3386 2652
rect 3398 2648 3402 2652
rect 3422 2648 3426 2652
rect 3446 2648 3450 2652
rect 3462 2648 3466 2652
rect 3374 2638 3378 2642
rect 3350 2598 3354 2602
rect 3366 2598 3370 2602
rect 3350 2588 3354 2592
rect 3334 2568 3338 2572
rect 3302 2558 3306 2562
rect 3326 2558 3330 2562
rect 3318 2548 3322 2552
rect 3334 2538 3338 2542
rect 3318 2528 3322 2532
rect 3398 2638 3402 2642
rect 3534 2608 3538 2612
rect 3494 2578 3498 2582
rect 3462 2568 3466 2572
rect 3486 2568 3490 2572
rect 3470 2558 3474 2562
rect 3414 2548 3418 2552
rect 3534 2558 3538 2562
rect 3710 2698 3714 2702
rect 3662 2688 3666 2692
rect 3726 2688 3730 2692
rect 3694 2678 3698 2682
rect 3646 2668 3650 2672
rect 3686 2668 3690 2672
rect 3622 2638 3626 2642
rect 3782 2938 3786 2942
rect 3806 2898 3810 2902
rect 3774 2868 3778 2872
rect 3758 2838 3762 2842
rect 3806 2798 3810 2802
rect 3750 2778 3754 2782
rect 3774 2738 3778 2742
rect 3742 2708 3746 2712
rect 3742 2678 3746 2682
rect 3766 2678 3770 2682
rect 3734 2668 3738 2672
rect 3782 2728 3786 2732
rect 3798 2718 3802 2722
rect 3790 2688 3794 2692
rect 3798 2688 3802 2692
rect 3814 2738 3818 2742
rect 3862 3288 3866 3292
rect 3934 3328 3938 3332
rect 4030 3328 4034 3332
rect 3982 3298 3986 3302
rect 4014 3288 4018 3292
rect 3894 3268 3898 3272
rect 3990 3268 3994 3272
rect 4022 3258 4026 3262
rect 3894 3147 3898 3151
rect 3918 3138 3922 3142
rect 4082 3303 4086 3307
rect 4089 3303 4093 3307
rect 4190 3438 4194 3442
rect 4222 3428 4226 3432
rect 4126 3368 4130 3372
rect 4246 3498 4250 3502
rect 4294 3498 4298 3502
rect 4206 3338 4210 3342
rect 4126 3318 4130 3322
rect 4214 3278 4218 3282
rect 4070 3198 4074 3202
rect 4006 3178 4010 3182
rect 4070 3168 4074 3172
rect 3950 3158 3954 3162
rect 3966 3148 3970 3152
rect 4046 3148 4050 3152
rect 4078 3148 4082 3152
rect 3982 3118 3986 3122
rect 3998 3078 4002 3082
rect 4214 3258 4218 3262
rect 4222 3208 4226 3212
rect 4142 3188 4146 3192
rect 4190 3188 4194 3192
rect 4206 3188 4210 3192
rect 4198 3158 4202 3162
rect 4078 3118 4082 3122
rect 4082 3103 4086 3107
rect 4089 3103 4093 3107
rect 3878 3058 3882 3062
rect 3854 2968 3858 2972
rect 3854 2958 3858 2962
rect 3846 2868 3850 2872
rect 3934 2988 3938 2992
rect 3998 2968 4002 2972
rect 3862 2888 3866 2892
rect 4094 3058 4098 3062
rect 4062 3048 4066 3052
rect 4030 3038 4034 3042
rect 4118 3128 4122 3132
rect 4110 3078 4114 3082
rect 4150 3088 4154 3092
rect 4150 3068 4154 3072
rect 4118 3058 4122 3062
rect 4174 3108 4178 3112
rect 4166 3058 4170 3062
rect 4158 3048 4162 3052
rect 4030 2928 4034 2932
rect 4082 2903 4086 2907
rect 4089 2903 4093 2907
rect 4142 2888 4146 2892
rect 3918 2878 3922 2882
rect 4206 3018 4210 3022
rect 4166 2948 4170 2952
rect 4182 2948 4186 2952
rect 4198 2918 4202 2922
rect 3966 2868 3970 2872
rect 4110 2868 4114 2872
rect 3870 2858 3874 2862
rect 3910 2858 3914 2862
rect 3926 2848 3930 2852
rect 3854 2838 3858 2842
rect 3950 2838 3954 2842
rect 3838 2798 3842 2802
rect 3982 2808 3986 2812
rect 3942 2758 3946 2762
rect 3998 2758 4002 2762
rect 3878 2747 3882 2751
rect 3918 2748 3922 2752
rect 3838 2718 3842 2722
rect 3830 2698 3834 2702
rect 4158 2858 4162 2862
rect 4078 2808 4082 2812
rect 4102 2788 4106 2792
rect 4174 2788 4178 2792
rect 4030 2768 4034 2772
rect 4038 2747 4042 2751
rect 4078 2748 4082 2752
rect 4142 2748 4146 2752
rect 4126 2738 4130 2742
rect 3926 2718 3930 2722
rect 3934 2698 3938 2702
rect 3966 2698 3970 2702
rect 3790 2668 3794 2672
rect 3894 2668 3898 2672
rect 3902 2668 3906 2672
rect 3750 2658 3754 2662
rect 3710 2648 3714 2652
rect 3742 2648 3746 2652
rect 3774 2648 3778 2652
rect 3838 2648 3842 2652
rect 3670 2628 3674 2632
rect 3886 2618 3890 2622
rect 3630 2608 3634 2612
rect 3646 2608 3650 2612
rect 3570 2603 3574 2607
rect 3577 2603 3581 2607
rect 3598 2578 3602 2582
rect 3622 2578 3626 2582
rect 3574 2568 3578 2572
rect 3566 2558 3570 2562
rect 3550 2548 3554 2552
rect 3430 2538 3434 2542
rect 3518 2538 3522 2542
rect 3558 2538 3562 2542
rect 3430 2528 3434 2532
rect 3486 2528 3490 2532
rect 3294 2488 3298 2492
rect 3430 2488 3434 2492
rect 3486 2488 3490 2492
rect 3342 2478 3346 2482
rect 3310 2468 3314 2472
rect 3230 2458 3234 2462
rect 3206 2448 3210 2452
rect 3214 2438 3218 2442
rect 3230 2408 3234 2412
rect 3246 2398 3250 2402
rect 3190 2388 3194 2392
rect 3214 2388 3218 2392
rect 3174 2378 3178 2382
rect 3094 2348 3098 2352
rect 3134 2348 3138 2352
rect 3110 2338 3114 2342
rect 3158 2338 3162 2342
rect 3438 2478 3442 2482
rect 3462 2478 3466 2482
rect 3478 2478 3482 2482
rect 3510 2478 3514 2482
rect 3478 2468 3482 2472
rect 3542 2528 3546 2532
rect 3598 2498 3602 2502
rect 3558 2488 3562 2492
rect 3574 2478 3578 2482
rect 3526 2468 3530 2472
rect 3542 2468 3546 2472
rect 3582 2468 3586 2472
rect 3694 2598 3698 2602
rect 3638 2568 3642 2572
rect 3646 2558 3650 2562
rect 3630 2538 3634 2542
rect 3670 2538 3674 2542
rect 3830 2568 3834 2572
rect 3734 2558 3738 2562
rect 3750 2558 3754 2562
rect 3758 2558 3762 2562
rect 3798 2558 3802 2562
rect 3822 2558 3826 2562
rect 3926 2658 3930 2662
rect 3902 2598 3906 2602
rect 3918 2628 3922 2632
rect 3982 2688 3986 2692
rect 3942 2678 3946 2682
rect 3982 2668 3986 2672
rect 3958 2658 3962 2662
rect 4350 3548 4354 3552
rect 4334 3518 4338 3522
rect 4462 3588 4466 3592
rect 4534 3578 4538 3582
rect 4566 3578 4570 3582
rect 4422 3568 4426 3572
rect 4518 3558 4522 3562
rect 4590 3558 4594 3562
rect 4510 3538 4514 3542
rect 4494 3528 4498 3532
rect 4406 3508 4410 3512
rect 4366 3478 4370 3482
rect 4382 3478 4386 3482
rect 4278 3468 4282 3472
rect 4350 3468 4354 3472
rect 4358 3468 4362 3472
rect 4254 3458 4258 3462
rect 4294 3458 4298 3462
rect 4326 3458 4330 3462
rect 4246 3268 4250 3272
rect 4310 3448 4314 3452
rect 4318 3378 4322 3382
rect 4310 3358 4314 3362
rect 4358 3448 4362 3452
rect 4374 3448 4378 3452
rect 4390 3458 4394 3462
rect 4382 3438 4386 3442
rect 4390 3438 4394 3442
rect 4334 3368 4338 3372
rect 4278 3348 4282 3352
rect 4326 3348 4330 3352
rect 4358 3348 4362 3352
rect 4270 3328 4274 3332
rect 4262 3268 4266 3272
rect 4254 3258 4258 3262
rect 4246 3248 4250 3252
rect 4254 3238 4258 3242
rect 4294 3338 4298 3342
rect 4310 3338 4314 3342
rect 4318 3308 4322 3312
rect 4342 3288 4346 3292
rect 4278 3258 4282 3262
rect 4262 3168 4266 3172
rect 4286 3158 4290 3162
rect 4278 3148 4282 3152
rect 4270 3108 4274 3112
rect 4294 3138 4298 3142
rect 4294 3108 4298 3112
rect 4278 3098 4282 3102
rect 4270 3078 4274 3082
rect 4302 3098 4306 3102
rect 4278 3068 4282 3072
rect 4302 3058 4306 3062
rect 4286 3048 4290 3052
rect 4278 3028 4282 3032
rect 4326 3218 4330 3222
rect 4326 3151 4330 3152
rect 4326 3148 4330 3151
rect 4366 3308 4370 3312
rect 4366 3278 4370 3282
rect 4366 3268 4370 3272
rect 4430 3468 4434 3472
rect 4454 3468 4458 3472
rect 4502 3458 4506 3462
rect 4518 3468 4522 3472
rect 4542 3458 4546 3462
rect 4430 3448 4434 3452
rect 4550 3448 4554 3452
rect 4398 3338 4402 3342
rect 4390 3228 4394 3232
rect 4350 3138 4354 3142
rect 4350 3128 4354 3132
rect 4390 3098 4394 3102
rect 4390 3078 4394 3082
rect 4350 3048 4354 3052
rect 4318 3038 4322 3042
rect 4294 2948 4298 2952
rect 4254 2938 4258 2942
rect 4270 2938 4274 2942
rect 4286 2938 4290 2942
rect 4254 2918 4258 2922
rect 4238 2908 4242 2912
rect 4318 2958 4322 2962
rect 4374 3048 4378 3052
rect 4414 3258 4418 3262
rect 4430 3238 4434 3242
rect 4406 3188 4410 3192
rect 4430 3178 4434 3182
rect 4414 3148 4418 3152
rect 4502 3438 4506 3442
rect 4526 3428 4530 3432
rect 4486 3378 4490 3382
rect 4454 3358 4458 3362
rect 4510 3358 4514 3362
rect 4542 3358 4546 3362
rect 4518 3348 4522 3352
rect 4478 3328 4482 3332
rect 4534 3328 4538 3332
rect 4566 3388 4570 3392
rect 4558 3348 4562 3352
rect 4478 3308 4482 3312
rect 4494 3308 4498 3312
rect 4510 3308 4514 3312
rect 4494 3298 4498 3302
rect 4526 3278 4530 3282
rect 4526 3268 4530 3272
rect 4558 3298 4562 3302
rect 4566 3288 4570 3292
rect 4542 3248 4546 3252
rect 4534 3168 4538 3172
rect 4566 3248 4570 3252
rect 4550 3158 4554 3162
rect 4566 3158 4570 3162
rect 4590 3158 4594 3162
rect 4438 3148 4442 3152
rect 4502 3148 4506 3152
rect 4406 3138 4410 3142
rect 4422 3138 4426 3142
rect 4462 3138 4466 3142
rect 4486 3138 4490 3142
rect 4510 3138 4514 3142
rect 4558 3138 4562 3142
rect 4446 3108 4450 3112
rect 4438 3088 4442 3092
rect 4486 3098 4490 3102
rect 4454 3068 4458 3072
rect 4478 3068 4482 3072
rect 4510 3068 4514 3072
rect 4542 3068 4546 3072
rect 4486 3058 4490 3062
rect 4534 3058 4538 3062
rect 4462 3038 4466 3042
rect 4470 3038 4474 3042
rect 4446 3028 4450 3032
rect 4406 2958 4410 2962
rect 4422 2958 4426 2962
rect 4326 2948 4330 2952
rect 4350 2948 4354 2952
rect 4406 2948 4410 2952
rect 4334 2938 4338 2942
rect 4310 2908 4314 2912
rect 4318 2868 4322 2872
rect 4398 2928 4402 2932
rect 4382 2918 4386 2922
rect 4358 2898 4362 2902
rect 4342 2878 4346 2882
rect 4358 2868 4362 2872
rect 4326 2858 4330 2862
rect 4382 2908 4386 2912
rect 4398 2878 4402 2882
rect 4566 3078 4570 3082
rect 4518 3048 4522 3052
rect 4526 3038 4530 3042
rect 4582 3058 4586 3062
rect 4558 3028 4562 3032
rect 4574 3028 4578 3032
rect 4558 2978 4562 2982
rect 4510 2968 4514 2972
rect 4574 2968 4578 2972
rect 4550 2948 4554 2952
rect 4462 2938 4466 2942
rect 4454 2918 4458 2922
rect 4518 2938 4522 2942
rect 4542 2938 4546 2942
rect 4566 2938 4570 2942
rect 4558 2898 4562 2902
rect 4486 2888 4490 2892
rect 4470 2878 4474 2882
rect 4582 2878 4586 2882
rect 4422 2868 4426 2872
rect 4398 2858 4402 2862
rect 4374 2848 4378 2852
rect 4414 2848 4418 2852
rect 4270 2828 4274 2832
rect 4238 2798 4242 2802
rect 4238 2758 4242 2762
rect 4262 2758 4266 2762
rect 4310 2758 4314 2762
rect 4206 2738 4210 2742
rect 4238 2738 4242 2742
rect 4038 2728 4042 2732
rect 4158 2728 4162 2732
rect 4082 2703 4086 2707
rect 4089 2703 4093 2707
rect 4126 2698 4130 2702
rect 4142 2698 4146 2702
rect 4230 2698 4234 2702
rect 4038 2688 4042 2692
rect 3998 2678 4002 2682
rect 4022 2678 4026 2682
rect 4118 2678 4122 2682
rect 4014 2668 4018 2672
rect 4046 2668 4050 2672
rect 4086 2668 4090 2672
rect 4086 2658 4090 2662
rect 3942 2648 3946 2652
rect 3966 2648 3970 2652
rect 4054 2648 4058 2652
rect 4062 2648 4066 2652
rect 3910 2568 3914 2572
rect 3926 2568 3930 2572
rect 4062 2638 4066 2642
rect 3958 2618 3962 2622
rect 4038 2578 4042 2582
rect 3942 2558 3946 2562
rect 3974 2558 3978 2562
rect 4006 2558 4010 2562
rect 3846 2538 3850 2542
rect 3894 2538 3898 2542
rect 3910 2538 3914 2542
rect 3926 2538 3930 2542
rect 3958 2538 3962 2542
rect 3974 2538 3978 2542
rect 3646 2518 3650 2522
rect 3686 2488 3690 2492
rect 3702 2518 3706 2522
rect 3718 2518 3722 2522
rect 3702 2498 3706 2502
rect 3638 2478 3642 2482
rect 3638 2468 3642 2472
rect 3686 2468 3690 2472
rect 3750 2508 3754 2512
rect 3822 2528 3826 2532
rect 3902 2518 3906 2522
rect 3966 2518 3970 2522
rect 3782 2498 3786 2502
rect 3814 2488 3818 2492
rect 3782 2478 3786 2482
rect 3838 2478 3842 2482
rect 3966 2488 3970 2492
rect 3894 2478 3898 2482
rect 3934 2478 3938 2482
rect 3750 2468 3754 2472
rect 3790 2468 3794 2472
rect 3814 2468 3818 2472
rect 3830 2468 3834 2472
rect 3334 2458 3338 2462
rect 3358 2458 3362 2462
rect 3518 2458 3522 2462
rect 3606 2458 3610 2462
rect 3662 2458 3666 2462
rect 3694 2458 3698 2462
rect 3286 2448 3290 2452
rect 3302 2448 3306 2452
rect 3326 2448 3330 2452
rect 3350 2448 3354 2452
rect 3302 2438 3306 2442
rect 3326 2438 3330 2442
rect 3358 2398 3362 2402
rect 3302 2388 3306 2392
rect 3350 2388 3354 2392
rect 3262 2368 3266 2372
rect 3438 2448 3442 2452
rect 3646 2448 3650 2452
rect 3654 2448 3658 2452
rect 3670 2448 3674 2452
rect 3710 2448 3714 2452
rect 3766 2458 3770 2462
rect 3806 2458 3810 2462
rect 3942 2458 3946 2462
rect 3750 2448 3754 2452
rect 3774 2448 3778 2452
rect 3846 2448 3850 2452
rect 3414 2438 3418 2442
rect 3526 2438 3530 2442
rect 3494 2428 3498 2432
rect 3398 2408 3402 2412
rect 3470 2388 3474 2392
rect 3366 2368 3370 2372
rect 3374 2368 3378 2372
rect 3206 2358 3210 2362
rect 3230 2358 3234 2362
rect 3310 2358 3314 2362
rect 3350 2358 3354 2362
rect 3262 2348 3266 2352
rect 3510 2378 3514 2382
rect 3558 2428 3562 2432
rect 3550 2378 3554 2382
rect 3570 2403 3574 2407
rect 3577 2403 3581 2407
rect 3798 2438 3802 2442
rect 3854 2438 3858 2442
rect 3838 2428 3842 2432
rect 3822 2398 3826 2402
rect 3742 2388 3746 2392
rect 3638 2378 3642 2382
rect 3670 2378 3674 2382
rect 3598 2358 3602 2362
rect 3630 2358 3634 2362
rect 3686 2358 3690 2362
rect 3710 2358 3714 2362
rect 3750 2358 3754 2362
rect 3806 2358 3810 2362
rect 3350 2348 3354 2352
rect 3406 2348 3410 2352
rect 3454 2348 3458 2352
rect 3486 2348 3490 2352
rect 3518 2348 3522 2352
rect 3550 2348 3554 2352
rect 3238 2338 3242 2342
rect 3270 2338 3274 2342
rect 3302 2338 3306 2342
rect 3366 2338 3370 2342
rect 3398 2338 3402 2342
rect 3438 2338 3442 2342
rect 3094 2328 3098 2332
rect 3118 2328 3122 2332
rect 3206 2328 3210 2332
rect 3270 2328 3274 2332
rect 3318 2328 3322 2332
rect 3374 2328 3378 2332
rect 3094 2268 3098 2272
rect 3102 2258 3106 2262
rect 3118 2258 3122 2262
rect 3150 2308 3154 2312
rect 3254 2318 3258 2322
rect 3174 2298 3178 2302
rect 3246 2298 3250 2302
rect 3302 2308 3306 2312
rect 3150 2278 3154 2282
rect 3206 2278 3210 2282
rect 3222 2278 3226 2282
rect 3238 2278 3242 2282
rect 3270 2278 3274 2282
rect 3142 2268 3146 2272
rect 3174 2268 3178 2272
rect 3190 2268 3194 2272
rect 3286 2268 3290 2272
rect 3182 2258 3186 2262
rect 3110 2248 3114 2252
rect 3134 2248 3138 2252
rect 3158 2248 3162 2252
rect 3174 2248 3178 2252
rect 3262 2248 3266 2252
rect 3230 2238 3234 2242
rect 3182 2218 3186 2222
rect 3230 2198 3234 2202
rect 3134 2188 3138 2192
rect 3118 2178 3122 2182
rect 3142 2178 3146 2182
rect 3078 2168 3082 2172
rect 2998 2138 3002 2142
rect 3030 2138 3034 2142
rect 2942 2128 2946 2132
rect 2878 2108 2882 2112
rect 2894 2108 2898 2112
rect 2870 2078 2874 2082
rect 2934 2098 2938 2102
rect 2958 2098 2962 2102
rect 2982 2118 2986 2122
rect 3038 2118 3042 2122
rect 2950 2088 2954 2092
rect 2942 2078 2946 2082
rect 2854 2068 2858 2072
rect 2878 2068 2882 2072
rect 2950 2068 2954 2072
rect 2774 2048 2778 2052
rect 2710 2028 2714 2032
rect 2750 2028 2754 2032
rect 2766 2028 2770 2032
rect 2662 2018 2666 2022
rect 2606 2008 2610 2012
rect 2646 2008 2650 2012
rect 2546 2003 2550 2007
rect 2553 2003 2557 2007
rect 2534 1988 2538 1992
rect 2630 1988 2634 1992
rect 2518 1958 2522 1962
rect 2534 1948 2538 1952
rect 2534 1928 2538 1932
rect 2478 1878 2482 1882
rect 2486 1878 2490 1882
rect 2366 1868 2370 1872
rect 2422 1858 2426 1862
rect 2446 1858 2450 1862
rect 2254 1848 2258 1852
rect 2262 1848 2266 1852
rect 2302 1848 2306 1852
rect 2526 1858 2530 1862
rect 2246 1828 2250 1832
rect 2254 1828 2258 1832
rect 2094 1808 2098 1812
rect 2134 1808 2138 1812
rect 2150 1808 2154 1812
rect 2238 1808 2242 1812
rect 2126 1768 2130 1772
rect 2134 1768 2138 1772
rect 2030 1738 2034 1742
rect 2118 1728 2122 1732
rect 2198 1798 2202 1802
rect 2158 1788 2162 1792
rect 2174 1768 2178 1772
rect 2286 1838 2290 1842
rect 2182 1758 2186 1762
rect 2214 1758 2218 1762
rect 2230 1758 2234 1762
rect 2246 1758 2250 1762
rect 2318 1758 2322 1762
rect 2174 1748 2178 1752
rect 2230 1748 2234 1752
rect 2262 1748 2266 1752
rect 2270 1748 2274 1752
rect 2246 1738 2250 1742
rect 2254 1738 2258 1742
rect 2318 1738 2322 1742
rect 2422 1848 2426 1852
rect 2430 1848 2434 1852
rect 2486 1848 2490 1852
rect 2510 1848 2514 1852
rect 2382 1768 2386 1772
rect 2406 1788 2410 1792
rect 2342 1758 2346 1762
rect 2486 1838 2490 1842
rect 2446 1768 2450 1772
rect 2470 1758 2474 1762
rect 2502 1828 2506 1832
rect 2358 1738 2362 1742
rect 2142 1728 2146 1732
rect 2190 1728 2194 1732
rect 2246 1728 2250 1732
rect 2294 1728 2298 1732
rect 2326 1728 2330 1732
rect 2366 1728 2370 1732
rect 1870 1718 1874 1722
rect 1894 1718 1898 1722
rect 1982 1718 1986 1722
rect 2078 1718 2082 1722
rect 2334 1718 2338 1722
rect 2342 1718 2346 1722
rect 1814 1688 1818 1692
rect 2286 1708 2290 1712
rect 2026 1703 2030 1707
rect 2033 1703 2037 1707
rect 1982 1698 1986 1702
rect 2278 1698 2282 1702
rect 1894 1688 1898 1692
rect 1790 1678 1794 1682
rect 1726 1648 1730 1652
rect 1694 1638 1698 1642
rect 1718 1638 1722 1642
rect 1734 1638 1738 1642
rect 1846 1678 1850 1682
rect 2046 1688 2050 1692
rect 2142 1688 2146 1692
rect 2150 1688 2154 1692
rect 2166 1688 2170 1692
rect 2262 1688 2266 1692
rect 1902 1678 1906 1682
rect 1966 1678 1970 1682
rect 1982 1678 1986 1682
rect 2110 1678 2114 1682
rect 1798 1668 1802 1672
rect 1830 1668 1834 1672
rect 1878 1668 1882 1672
rect 1934 1668 1938 1672
rect 1950 1668 1954 1672
rect 1990 1668 1994 1672
rect 2094 1668 2098 1672
rect 1910 1658 1914 1662
rect 1766 1648 1770 1652
rect 1774 1648 1778 1652
rect 1854 1648 1858 1652
rect 1758 1638 1762 1642
rect 1830 1638 1834 1642
rect 1886 1638 1890 1642
rect 1742 1608 1746 1612
rect 1702 1588 1706 1592
rect 1718 1588 1722 1592
rect 1654 1528 1658 1532
rect 1678 1518 1682 1522
rect 1694 1518 1698 1522
rect 1726 1578 1730 1582
rect 1718 1538 1722 1542
rect 1710 1508 1714 1512
rect 1646 1488 1650 1492
rect 1702 1488 1706 1492
rect 1654 1478 1658 1482
rect 1662 1468 1666 1472
rect 1702 1468 1706 1472
rect 1750 1548 1754 1552
rect 1766 1548 1770 1552
rect 1742 1488 1746 1492
rect 1750 1478 1754 1482
rect 1710 1458 1714 1462
rect 1726 1458 1730 1462
rect 1678 1448 1682 1452
rect 1646 1438 1650 1442
rect 1638 1428 1642 1432
rect 1598 1418 1602 1422
rect 1646 1418 1650 1422
rect 1590 1378 1594 1382
rect 1678 1378 1682 1382
rect 1598 1368 1602 1372
rect 1590 1358 1594 1362
rect 1670 1348 1674 1352
rect 1630 1338 1634 1342
rect 1558 1328 1562 1332
rect 1590 1328 1594 1332
rect 1606 1328 1610 1332
rect 1662 1328 1666 1332
rect 1582 1298 1586 1302
rect 1654 1288 1658 1292
rect 1558 1278 1562 1282
rect 1574 1278 1578 1282
rect 1614 1278 1618 1282
rect 1630 1278 1634 1282
rect 1638 1268 1642 1272
rect 1614 1258 1618 1262
rect 1670 1258 1674 1262
rect 1590 1248 1594 1252
rect 1606 1248 1610 1252
rect 1614 1248 1618 1252
rect 1630 1248 1634 1252
rect 1654 1248 1658 1252
rect 1590 1238 1594 1242
rect 1598 1188 1602 1192
rect 1630 1238 1634 1242
rect 1614 1228 1618 1232
rect 1606 1178 1610 1182
rect 1606 1168 1610 1172
rect 1550 1148 1554 1152
rect 1526 1138 1530 1142
rect 1446 1128 1450 1132
rect 1486 1118 1490 1122
rect 1422 1098 1426 1102
rect 1430 1088 1434 1092
rect 1382 1078 1386 1082
rect 1406 1078 1410 1082
rect 1326 1048 1330 1052
rect 1342 1038 1346 1042
rect 1382 1058 1386 1062
rect 1422 1058 1426 1062
rect 1390 1028 1394 1032
rect 1414 1028 1418 1032
rect 1478 1098 1482 1102
rect 1494 1088 1498 1092
rect 1446 1068 1450 1072
rect 1470 1068 1474 1072
rect 1550 1108 1554 1112
rect 1622 1158 1626 1162
rect 1542 1098 1546 1102
rect 1614 1098 1618 1102
rect 1438 1058 1442 1062
rect 1478 1058 1482 1062
rect 1462 1038 1466 1042
rect 1374 978 1378 982
rect 1446 978 1450 982
rect 1366 958 1370 962
rect 1438 958 1442 962
rect 1430 948 1434 952
rect 1558 1078 1562 1082
rect 1502 1058 1506 1062
rect 1494 1048 1498 1052
rect 1486 978 1490 982
rect 1470 958 1474 962
rect 1478 958 1482 962
rect 1522 1003 1526 1007
rect 1529 1003 1533 1007
rect 1510 988 1514 992
rect 1582 1058 1586 1062
rect 1558 1008 1562 1012
rect 1566 968 1570 972
rect 1542 958 1546 962
rect 1478 948 1482 952
rect 1494 948 1498 952
rect 1350 938 1354 942
rect 1414 928 1418 932
rect 1398 918 1402 922
rect 1462 918 1466 922
rect 1398 898 1402 902
rect 1334 888 1338 892
rect 1382 888 1386 892
rect 1318 878 1322 882
rect 1190 868 1194 872
rect 1206 868 1210 872
rect 1246 868 1250 872
rect 1294 868 1298 872
rect 1326 868 1330 872
rect 1166 858 1170 862
rect 1230 858 1234 862
rect 1190 848 1194 852
rect 1222 848 1226 852
rect 1158 768 1162 772
rect 1094 748 1098 752
rect 1206 758 1210 762
rect 1070 738 1074 742
rect 1158 738 1162 742
rect 1174 738 1178 742
rect 1278 858 1282 862
rect 1270 848 1274 852
rect 1318 848 1322 852
rect 1326 818 1330 822
rect 1270 768 1274 772
rect 1254 748 1258 752
rect 1246 738 1250 742
rect 1350 878 1354 882
rect 1430 878 1434 882
rect 1438 868 1442 872
rect 1494 918 1498 922
rect 1550 948 1554 952
rect 1470 908 1474 912
rect 1510 908 1514 912
rect 1518 908 1522 912
rect 1566 898 1570 902
rect 1574 898 1578 902
rect 1470 888 1474 892
rect 1598 1048 1602 1052
rect 1590 1028 1594 1032
rect 1590 948 1594 952
rect 1598 888 1602 892
rect 1470 868 1474 872
rect 1350 848 1354 852
rect 1398 848 1402 852
rect 1462 858 1466 862
rect 1422 838 1426 842
rect 1462 838 1466 842
rect 1342 818 1346 822
rect 1342 768 1346 772
rect 1366 768 1370 772
rect 1350 758 1354 762
rect 1374 758 1378 762
rect 1374 748 1378 752
rect 1422 748 1426 752
rect 1470 768 1474 772
rect 1342 738 1346 742
rect 1430 738 1434 742
rect 1022 718 1026 722
rect 1002 703 1006 707
rect 1009 703 1013 707
rect 990 688 994 692
rect 1014 688 1018 692
rect 966 678 970 682
rect 894 668 898 672
rect 806 658 810 662
rect 902 648 906 652
rect 894 598 898 602
rect 902 598 906 602
rect 846 568 850 572
rect 798 558 802 562
rect 838 558 842 562
rect 774 538 778 542
rect 774 488 778 492
rect 702 458 706 462
rect 686 448 690 452
rect 670 438 674 442
rect 678 438 682 442
rect 702 438 706 442
rect 694 428 698 432
rect 702 428 706 432
rect 710 428 714 432
rect 686 358 690 362
rect 798 538 802 542
rect 814 498 818 502
rect 790 458 794 462
rect 798 458 802 462
rect 766 448 770 452
rect 734 378 738 382
rect 742 378 746 382
rect 790 378 794 382
rect 750 348 754 352
rect 662 318 666 322
rect 742 338 746 342
rect 758 338 762 342
rect 790 328 794 332
rect 726 318 730 322
rect 702 308 706 312
rect 646 298 650 302
rect 678 298 682 302
rect 702 298 706 302
rect 630 268 634 272
rect 630 248 634 252
rect 614 198 618 202
rect 574 168 578 172
rect 582 168 586 172
rect 486 138 490 142
rect 526 138 530 142
rect 558 148 562 152
rect 606 148 610 152
rect 574 138 578 142
rect 598 138 602 142
rect 550 128 554 132
rect 646 258 650 262
rect 750 288 754 292
rect 702 258 706 262
rect 726 248 730 252
rect 662 208 666 212
rect 806 358 810 362
rect 878 558 882 562
rect 862 518 866 522
rect 902 548 906 552
rect 878 478 882 482
rect 982 618 986 622
rect 950 598 954 602
rect 902 538 906 542
rect 942 538 946 542
rect 934 478 938 482
rect 894 468 898 472
rect 886 458 890 462
rect 878 448 882 452
rect 894 448 898 452
rect 862 398 866 402
rect 998 568 1002 572
rect 998 558 1002 562
rect 1086 728 1090 732
rect 1118 718 1122 722
rect 1030 708 1034 712
rect 1126 708 1130 712
rect 1046 688 1050 692
rect 1070 688 1074 692
rect 1054 678 1058 682
rect 1158 708 1162 712
rect 1174 708 1178 712
rect 1142 698 1146 702
rect 1198 728 1202 732
rect 1222 728 1226 732
rect 1246 728 1250 732
rect 1214 718 1218 722
rect 1286 718 1290 722
rect 1206 708 1210 712
rect 1182 688 1186 692
rect 1190 678 1194 682
rect 1222 708 1226 712
rect 1238 698 1242 702
rect 1238 678 1242 682
rect 1062 668 1066 672
rect 1126 668 1130 672
rect 1198 668 1202 672
rect 1342 728 1346 732
rect 1398 708 1402 712
rect 1302 698 1306 702
rect 1326 698 1330 702
rect 1398 698 1402 702
rect 1286 688 1290 692
rect 1310 688 1314 692
rect 1278 678 1282 682
rect 1318 668 1322 672
rect 1118 658 1122 662
rect 1174 658 1178 662
rect 1366 678 1370 682
rect 1382 678 1386 682
rect 1438 698 1442 702
rect 1334 668 1338 672
rect 1342 668 1346 672
rect 1358 668 1362 672
rect 1422 668 1426 672
rect 1590 878 1594 882
rect 1662 1218 1666 1222
rect 1646 1178 1650 1182
rect 1678 1208 1682 1212
rect 1702 1438 1706 1442
rect 1718 1388 1722 1392
rect 1742 1378 1746 1382
rect 1766 1468 1770 1472
rect 1798 1618 1802 1622
rect 1886 1598 1890 1602
rect 1910 1598 1914 1602
rect 1862 1578 1866 1582
rect 1870 1578 1874 1582
rect 1886 1578 1890 1582
rect 1814 1568 1818 1572
rect 1830 1568 1834 1572
rect 1862 1558 1866 1562
rect 1790 1548 1794 1552
rect 1814 1548 1818 1552
rect 1782 1508 1786 1512
rect 1790 1498 1794 1502
rect 1854 1548 1858 1552
rect 1838 1538 1842 1542
rect 1870 1538 1874 1542
rect 1990 1648 1994 1652
rect 1990 1638 1994 1642
rect 2174 1678 2178 1682
rect 2182 1678 2186 1682
rect 2222 1678 2226 1682
rect 2246 1678 2250 1682
rect 2070 1658 2074 1662
rect 2110 1658 2114 1662
rect 2142 1658 2146 1662
rect 2206 1658 2210 1662
rect 2126 1648 2130 1652
rect 2238 1648 2242 1652
rect 2078 1638 2082 1642
rect 2094 1638 2098 1642
rect 2006 1618 2010 1622
rect 2054 1618 2058 1622
rect 1950 1578 1954 1582
rect 2006 1578 2010 1582
rect 1966 1568 1970 1572
rect 1950 1558 1954 1562
rect 2078 1568 2082 1572
rect 2022 1558 2026 1562
rect 1926 1548 1930 1552
rect 1966 1548 1970 1552
rect 1974 1548 1978 1552
rect 1894 1538 1898 1542
rect 1910 1538 1914 1542
rect 1918 1488 1922 1492
rect 1926 1488 1930 1492
rect 1902 1468 1906 1472
rect 1918 1468 1922 1472
rect 1814 1458 1818 1462
rect 1878 1458 1882 1462
rect 1830 1448 1834 1452
rect 1862 1448 1866 1452
rect 1958 1538 1962 1542
rect 2030 1538 2034 1542
rect 1982 1508 1986 1512
rect 1990 1488 1994 1492
rect 1934 1478 1938 1482
rect 1974 1478 1978 1482
rect 2026 1503 2030 1507
rect 2033 1503 2037 1507
rect 2150 1598 2154 1602
rect 2134 1568 2138 1572
rect 2238 1588 2242 1592
rect 2246 1588 2250 1592
rect 2246 1558 2250 1562
rect 2126 1548 2130 1552
rect 2142 1548 2146 1552
rect 2158 1548 2162 1552
rect 2198 1548 2202 1552
rect 2214 1548 2218 1552
rect 2238 1548 2242 1552
rect 2078 1538 2082 1542
rect 2118 1538 2122 1542
rect 2198 1538 2202 1542
rect 2230 1538 2234 1542
rect 2262 1538 2266 1542
rect 2102 1528 2106 1532
rect 2166 1518 2170 1522
rect 2054 1488 2058 1492
rect 2014 1478 2018 1482
rect 2086 1478 2090 1482
rect 2102 1478 2106 1482
rect 2142 1478 2146 1482
rect 1950 1468 1954 1472
rect 2070 1468 2074 1472
rect 2086 1466 2090 1470
rect 1958 1458 1962 1462
rect 2086 1458 2090 1462
rect 2102 1458 2106 1462
rect 1982 1448 1986 1452
rect 2030 1448 2034 1452
rect 1798 1438 1802 1442
rect 1870 1438 1874 1442
rect 1886 1438 1890 1442
rect 1766 1398 1770 1402
rect 1758 1358 1762 1362
rect 1798 1388 1802 1392
rect 1870 1408 1874 1412
rect 1878 1388 1882 1392
rect 1902 1388 1906 1392
rect 1814 1378 1818 1382
rect 1862 1368 1866 1372
rect 1894 1368 1898 1372
rect 1774 1358 1778 1362
rect 1790 1358 1794 1362
rect 1814 1358 1818 1362
rect 1702 1348 1706 1352
rect 1742 1348 1746 1352
rect 1758 1348 1762 1352
rect 1790 1348 1794 1352
rect 1814 1348 1818 1352
rect 1846 1348 1850 1352
rect 1886 1348 1890 1352
rect 1774 1328 1778 1332
rect 1830 1328 1834 1332
rect 1846 1328 1850 1332
rect 1726 1308 1730 1312
rect 1694 1298 1698 1302
rect 1702 1258 1706 1262
rect 1750 1308 1754 1312
rect 1886 1328 1890 1332
rect 1902 1318 1906 1322
rect 1830 1288 1834 1292
rect 1862 1288 1866 1292
rect 1870 1288 1874 1292
rect 1902 1288 1906 1292
rect 1822 1278 1826 1282
rect 1886 1278 1890 1282
rect 1718 1258 1722 1262
rect 1726 1258 1730 1262
rect 1742 1258 1746 1262
rect 1750 1258 1754 1262
rect 1798 1258 1802 1262
rect 1710 1238 1714 1242
rect 1750 1248 1754 1252
rect 1734 1228 1738 1232
rect 1742 1208 1746 1212
rect 1718 1198 1722 1202
rect 1686 1188 1690 1192
rect 1718 1188 1722 1192
rect 1670 1178 1674 1182
rect 1734 1158 1738 1162
rect 1694 1148 1698 1152
rect 1662 1138 1666 1142
rect 1686 1138 1690 1142
rect 1646 1128 1650 1132
rect 1678 1128 1682 1132
rect 1638 1068 1642 1072
rect 1630 1058 1634 1062
rect 1622 1048 1626 1052
rect 1678 1108 1682 1112
rect 1686 1108 1690 1112
rect 1654 1088 1658 1092
rect 1654 1078 1658 1082
rect 1694 1098 1698 1102
rect 1646 1038 1650 1042
rect 1686 1028 1690 1032
rect 1670 978 1674 982
rect 1726 1058 1730 1062
rect 1710 1048 1714 1052
rect 1710 998 1714 1002
rect 1702 968 1706 972
rect 1670 958 1674 962
rect 1726 958 1730 962
rect 1614 948 1618 952
rect 1694 948 1698 952
rect 1662 938 1666 942
rect 1710 938 1714 942
rect 1718 938 1722 942
rect 1670 928 1674 932
rect 1630 908 1634 912
rect 1638 898 1642 902
rect 1622 868 1626 872
rect 1638 868 1642 872
rect 1558 858 1562 862
rect 1574 858 1578 862
rect 1534 838 1538 842
rect 1510 818 1514 822
rect 1522 803 1526 807
rect 1529 803 1533 807
rect 1486 768 1490 772
rect 1518 768 1522 772
rect 1502 728 1506 732
rect 1478 698 1482 702
rect 1494 678 1498 682
rect 1382 658 1386 662
rect 1158 648 1162 652
rect 1102 618 1106 622
rect 1134 618 1138 622
rect 1150 608 1154 612
rect 1070 578 1074 582
rect 966 538 970 542
rect 1102 538 1106 542
rect 1142 528 1146 532
rect 1166 548 1170 552
rect 1002 503 1006 507
rect 1009 503 1013 507
rect 958 468 962 472
rect 1030 468 1034 472
rect 910 438 914 442
rect 982 438 986 442
rect 902 368 906 372
rect 902 358 906 362
rect 934 368 938 372
rect 854 338 858 342
rect 838 298 842 302
rect 814 268 818 272
rect 782 258 786 262
rect 798 258 802 262
rect 846 288 850 292
rect 870 318 874 322
rect 870 288 874 292
rect 854 278 858 282
rect 798 248 802 252
rect 830 248 834 252
rect 846 248 850 252
rect 814 238 818 242
rect 774 228 778 232
rect 718 198 722 202
rect 678 188 682 192
rect 702 188 706 192
rect 910 268 914 272
rect 934 268 938 272
rect 886 258 890 262
rect 918 258 922 262
rect 1006 378 1010 382
rect 1014 318 1018 322
rect 1002 303 1006 307
rect 1009 303 1013 307
rect 958 298 962 302
rect 894 248 898 252
rect 934 248 938 252
rect 878 218 882 222
rect 622 158 626 162
rect 630 158 634 162
rect 758 178 762 182
rect 646 148 650 152
rect 614 138 618 142
rect 638 138 642 142
rect 702 138 706 142
rect 718 138 722 142
rect 622 128 626 132
rect 710 128 714 132
rect 598 118 602 122
rect 446 88 450 92
rect 406 78 410 82
rect 198 58 202 62
rect 350 58 354 62
rect 398 59 402 63
rect 486 58 490 62
rect 6 48 10 52
rect 498 3 502 7
rect 505 3 509 7
rect 574 78 578 82
rect 734 98 738 102
rect 654 78 658 82
rect 582 58 586 62
rect 630 58 634 62
rect 678 59 682 63
rect 862 168 866 172
rect 902 158 906 162
rect 854 148 858 152
rect 950 248 954 252
rect 1094 458 1098 462
rect 1406 648 1410 652
rect 1390 638 1394 642
rect 1270 628 1274 632
rect 1262 568 1266 572
rect 1222 538 1226 542
rect 1246 528 1250 532
rect 1206 488 1210 492
rect 1326 618 1330 622
rect 1470 588 1474 592
rect 1486 588 1490 592
rect 1390 578 1394 582
rect 1398 578 1402 582
rect 1382 568 1386 572
rect 1326 528 1330 532
rect 1366 528 1370 532
rect 1382 508 1386 512
rect 1278 498 1282 502
rect 1342 498 1346 502
rect 1390 498 1394 502
rect 1326 478 1330 482
rect 1382 478 1386 482
rect 1438 568 1442 572
rect 1470 568 1474 572
rect 1550 728 1554 732
rect 1566 758 1570 762
rect 1782 1168 1786 1172
rect 1974 1438 1978 1442
rect 2030 1438 2034 1442
rect 1958 1418 1962 1422
rect 1918 1368 1922 1372
rect 1942 1348 1946 1352
rect 1934 1328 1938 1332
rect 1918 1318 1922 1322
rect 1926 1318 1930 1322
rect 1910 1278 1914 1282
rect 1838 1268 1842 1272
rect 1870 1268 1874 1272
rect 1894 1268 1898 1272
rect 1902 1268 1906 1272
rect 1926 1268 1930 1272
rect 1862 1258 1866 1262
rect 1806 1248 1810 1252
rect 1838 1248 1842 1252
rect 1894 1228 1898 1232
rect 1854 1218 1858 1222
rect 1886 1218 1890 1222
rect 1822 1178 1826 1182
rect 1798 1158 1802 1162
rect 1766 1138 1770 1142
rect 1766 1088 1770 1092
rect 1790 1148 1794 1152
rect 1790 1108 1794 1112
rect 1782 1088 1786 1092
rect 1790 1088 1794 1092
rect 1774 1078 1778 1082
rect 1774 1068 1778 1072
rect 1758 1048 1762 1052
rect 1766 1018 1770 1022
rect 1750 978 1754 982
rect 1806 1148 1810 1152
rect 1782 978 1786 982
rect 1798 958 1802 962
rect 1766 948 1770 952
rect 1766 938 1770 942
rect 1742 928 1746 932
rect 1702 918 1706 922
rect 1734 918 1738 922
rect 1782 928 1786 932
rect 1686 888 1690 892
rect 1686 878 1690 882
rect 1702 868 1706 872
rect 1726 868 1730 872
rect 1758 868 1762 872
rect 1630 858 1634 862
rect 1734 858 1738 862
rect 1598 788 1602 792
rect 1622 848 1626 852
rect 1694 848 1698 852
rect 1734 848 1738 852
rect 1718 838 1722 842
rect 1726 838 1730 842
rect 1694 778 1698 782
rect 1574 728 1578 732
rect 1522 603 1526 607
rect 1529 603 1533 607
rect 1566 668 1570 672
rect 1574 658 1578 662
rect 1510 568 1514 572
rect 1558 568 1562 572
rect 1414 548 1418 552
rect 1494 548 1498 552
rect 1518 548 1522 552
rect 1606 758 1610 762
rect 1654 748 1658 752
rect 1622 738 1626 742
rect 1646 738 1650 742
rect 1662 738 1666 742
rect 1678 738 1682 742
rect 1670 728 1674 732
rect 1622 718 1626 722
rect 1630 688 1634 692
rect 1646 688 1650 692
rect 1614 678 1618 682
rect 1694 708 1698 712
rect 1678 688 1682 692
rect 1686 678 1690 682
rect 1638 668 1642 672
rect 1654 668 1658 672
rect 1630 658 1634 662
rect 1646 658 1650 662
rect 1606 628 1610 632
rect 1718 758 1722 762
rect 1726 748 1730 752
rect 1750 848 1754 852
rect 1782 848 1786 852
rect 1790 848 1794 852
rect 1798 838 1802 842
rect 1838 1168 1842 1172
rect 1846 1148 1850 1152
rect 1830 1128 1834 1132
rect 1846 1088 1850 1092
rect 1846 1078 1850 1082
rect 1886 1188 1890 1192
rect 1870 1168 1874 1172
rect 1878 1148 1882 1152
rect 1894 1178 1898 1182
rect 1894 1138 1898 1142
rect 1870 1108 1874 1112
rect 1990 1368 1994 1372
rect 2014 1368 2018 1372
rect 1950 1328 1954 1332
rect 1942 1308 1946 1312
rect 1958 1298 1962 1302
rect 1950 1278 1954 1282
rect 1910 1258 1914 1262
rect 1934 1258 1938 1262
rect 1918 1248 1922 1252
rect 1926 1228 1930 1232
rect 1974 1328 1978 1332
rect 2006 1328 2010 1332
rect 1990 1318 1994 1322
rect 2006 1318 2010 1322
rect 1966 1288 1970 1292
rect 1974 1278 1978 1282
rect 1974 1270 1978 1272
rect 1974 1268 1978 1270
rect 1990 1258 1994 1262
rect 1950 1218 1954 1222
rect 1926 1198 1930 1202
rect 1942 1188 1946 1192
rect 1926 1178 1930 1182
rect 1934 1158 1938 1162
rect 1918 1128 1922 1132
rect 1918 1118 1922 1122
rect 1886 1078 1890 1082
rect 1934 1078 1938 1082
rect 1846 1058 1850 1062
rect 1830 1048 1834 1052
rect 1854 1048 1858 1052
rect 1830 1008 1834 1012
rect 1814 968 1818 972
rect 1838 998 1842 1002
rect 1902 1068 1906 1072
rect 1926 1058 1930 1062
rect 1878 1028 1882 1032
rect 1886 1028 1890 1032
rect 1886 998 1890 1002
rect 1982 1238 1986 1242
rect 1974 1208 1978 1212
rect 1958 1158 1962 1162
rect 1950 1148 1954 1152
rect 1966 1148 1970 1152
rect 1958 1128 1962 1132
rect 2006 1218 2010 1222
rect 1998 1188 2002 1192
rect 1982 1108 1986 1112
rect 1998 1128 2002 1132
rect 1990 1098 1994 1102
rect 1998 1078 2002 1082
rect 1990 1068 1994 1072
rect 1958 1058 1962 1062
rect 1998 1008 2002 1012
rect 1854 988 1858 992
rect 1870 988 1874 992
rect 1902 988 1906 992
rect 1846 968 1850 972
rect 1886 968 1890 972
rect 1942 968 1946 972
rect 2046 1318 2050 1322
rect 2026 1303 2030 1307
rect 2033 1303 2037 1307
rect 2174 1508 2178 1512
rect 2190 1508 2194 1512
rect 2246 1508 2250 1512
rect 2206 1488 2210 1492
rect 2238 1488 2242 1492
rect 2174 1478 2178 1482
rect 2150 1468 2154 1472
rect 2206 1468 2210 1472
rect 2222 1468 2226 1472
rect 2142 1458 2146 1462
rect 2158 1458 2162 1462
rect 2190 1458 2194 1462
rect 2214 1458 2218 1462
rect 2222 1448 2226 1452
rect 2198 1438 2202 1442
rect 2206 1438 2210 1442
rect 2230 1438 2234 1442
rect 2126 1428 2130 1432
rect 2166 1408 2170 1412
rect 2102 1398 2106 1402
rect 2070 1368 2074 1372
rect 2110 1378 2114 1382
rect 2182 1388 2186 1392
rect 2214 1378 2218 1382
rect 2198 1368 2202 1372
rect 2142 1358 2146 1362
rect 2182 1358 2186 1362
rect 2134 1348 2138 1352
rect 2150 1348 2154 1352
rect 2302 1688 2306 1692
rect 2358 1698 2362 1702
rect 2382 1698 2386 1702
rect 2350 1678 2354 1682
rect 2310 1668 2314 1672
rect 2350 1658 2354 1662
rect 2382 1668 2386 1672
rect 2470 1738 2474 1742
rect 2486 1738 2490 1742
rect 2606 1938 2610 1942
rect 2622 1940 2626 1944
rect 2558 1928 2562 1932
rect 2598 1908 2602 1912
rect 2566 1888 2570 1892
rect 2598 1858 2602 1862
rect 2558 1848 2562 1852
rect 2598 1848 2602 1852
rect 2622 1908 2626 1912
rect 2670 1958 2674 1962
rect 2670 1948 2674 1952
rect 2686 1948 2690 1952
rect 2686 1928 2690 1932
rect 2654 1918 2658 1922
rect 2638 1908 2642 1912
rect 2630 1888 2634 1892
rect 2630 1868 2634 1872
rect 2662 1868 2666 1872
rect 2726 2008 2730 2012
rect 2710 1948 2714 1952
rect 2750 1988 2754 1992
rect 2934 2058 2938 2062
rect 2862 2048 2866 2052
rect 2894 2048 2898 2052
rect 2918 2048 2922 2052
rect 2926 2048 2930 2052
rect 2950 2048 2954 2052
rect 3050 2103 3054 2107
rect 3057 2103 3061 2107
rect 3078 2138 3082 2142
rect 3134 2148 3138 2152
rect 3110 2128 3114 2132
rect 3118 2128 3122 2132
rect 3102 2118 3106 2122
rect 3118 2118 3122 2122
rect 3094 2098 3098 2102
rect 3134 2108 3138 2112
rect 3046 2088 3050 2092
rect 3102 2088 3106 2092
rect 3134 2088 3138 2092
rect 2982 2068 2986 2072
rect 3006 2068 3010 2072
rect 3014 2058 3018 2062
rect 3078 2058 3082 2062
rect 3094 2058 3098 2062
rect 3110 2058 3114 2062
rect 2814 2028 2818 2032
rect 2870 2028 2874 2032
rect 2974 2028 2978 2032
rect 2886 2018 2890 2022
rect 3022 2018 3026 2022
rect 3086 2018 3090 2022
rect 2878 2008 2882 2012
rect 2862 1978 2866 1982
rect 2838 1958 2842 1962
rect 2894 1998 2898 2002
rect 2766 1948 2770 1952
rect 2878 1948 2882 1952
rect 2886 1948 2890 1952
rect 2726 1940 2730 1944
rect 2854 1938 2858 1942
rect 2734 1928 2738 1932
rect 2750 1928 2754 1932
rect 2798 1928 2802 1932
rect 2838 1928 2842 1932
rect 2702 1918 2706 1922
rect 2886 1918 2890 1922
rect 2694 1878 2698 1882
rect 2694 1858 2698 1862
rect 2614 1838 2618 1842
rect 2646 1838 2650 1842
rect 2670 1838 2674 1842
rect 2566 1818 2570 1822
rect 2546 1803 2550 1807
rect 2553 1803 2557 1807
rect 2534 1798 2538 1802
rect 2494 1728 2498 1732
rect 2518 1728 2522 1732
rect 2534 1728 2538 1732
rect 2446 1718 2450 1722
rect 2430 1688 2434 1692
rect 2398 1668 2402 1672
rect 2422 1668 2426 1672
rect 2390 1658 2394 1662
rect 2390 1638 2394 1642
rect 2286 1598 2290 1602
rect 2294 1578 2298 1582
rect 2278 1558 2282 1562
rect 2286 1558 2290 1562
rect 2318 1558 2322 1562
rect 2278 1538 2282 1542
rect 2294 1538 2298 1542
rect 2310 1528 2314 1532
rect 2278 1518 2282 1522
rect 2270 1478 2274 1482
rect 2254 1468 2258 1472
rect 2286 1508 2290 1512
rect 2302 1508 2306 1512
rect 2286 1478 2290 1482
rect 2262 1458 2266 1462
rect 2390 1588 2394 1592
rect 2366 1578 2370 1582
rect 2398 1558 2402 1562
rect 2342 1548 2346 1552
rect 2382 1548 2386 1552
rect 2414 1548 2418 1552
rect 2350 1538 2354 1542
rect 2398 1538 2402 1542
rect 2358 1528 2362 1532
rect 2334 1518 2338 1522
rect 2326 1508 2330 1512
rect 2350 1498 2354 1502
rect 2318 1468 2322 1472
rect 2342 1468 2346 1472
rect 2326 1458 2330 1462
rect 2358 1458 2362 1462
rect 2310 1448 2314 1452
rect 2350 1448 2354 1452
rect 2342 1438 2346 1442
rect 2390 1508 2394 1512
rect 2414 1488 2418 1492
rect 2430 1618 2434 1622
rect 2454 1678 2458 1682
rect 2470 1678 2474 1682
rect 2438 1588 2442 1592
rect 2430 1518 2434 1522
rect 2438 1488 2442 1492
rect 2454 1668 2458 1672
rect 2518 1688 2522 1692
rect 2574 1808 2578 1812
rect 2646 1798 2650 1802
rect 2614 1768 2618 1772
rect 2646 1768 2650 1772
rect 2670 1768 2674 1772
rect 2590 1758 2594 1762
rect 2734 1908 2738 1912
rect 2710 1888 2714 1892
rect 2798 1888 2802 1892
rect 2870 1888 2874 1892
rect 2742 1878 2746 1882
rect 2766 1878 2770 1882
rect 2878 1878 2882 1882
rect 3150 2168 3154 2172
rect 3246 2168 3250 2172
rect 3182 2138 3186 2142
rect 3158 2128 3162 2132
rect 3174 2128 3178 2132
rect 3158 2098 3162 2102
rect 3222 2148 3226 2152
rect 3294 2238 3298 2242
rect 3262 2188 3266 2192
rect 3270 2168 3274 2172
rect 3214 2138 3218 2142
rect 3206 2098 3210 2102
rect 3214 2098 3218 2102
rect 3238 2098 3242 2102
rect 3214 2088 3218 2092
rect 3278 2138 3282 2142
rect 3254 2128 3258 2132
rect 3270 2128 3274 2132
rect 3310 2278 3314 2282
rect 3430 2328 3434 2332
rect 3454 2328 3458 2332
rect 3382 2298 3386 2302
rect 3406 2298 3410 2302
rect 3502 2328 3506 2332
rect 3430 2278 3434 2282
rect 3334 2268 3338 2272
rect 3366 2268 3370 2272
rect 3326 2258 3330 2262
rect 3302 2218 3306 2222
rect 3302 2178 3306 2182
rect 3342 2248 3346 2252
rect 3358 2238 3362 2242
rect 3318 2138 3322 2142
rect 3334 2128 3338 2132
rect 3318 2118 3322 2122
rect 3278 2088 3282 2092
rect 3182 2068 3186 2072
rect 3190 2058 3194 2062
rect 3222 2058 3226 2062
rect 3150 2048 3154 2052
rect 3174 2048 3178 2052
rect 3230 2048 3234 2052
rect 3254 2058 3258 2062
rect 3286 2058 3290 2062
rect 3182 2028 3186 2032
rect 3246 2028 3250 2032
rect 3262 2028 3266 2032
rect 3142 1998 3146 2002
rect 3014 1988 3018 1992
rect 3174 1988 3178 1992
rect 2966 1978 2970 1982
rect 2910 1958 2914 1962
rect 2902 1948 2906 1952
rect 2942 1938 2946 1942
rect 2934 1928 2938 1932
rect 2942 1878 2946 1882
rect 2774 1858 2778 1862
rect 2790 1858 2794 1862
rect 2718 1848 2722 1852
rect 2710 1808 2714 1812
rect 2694 1798 2698 1802
rect 2662 1758 2666 1762
rect 2686 1758 2690 1762
rect 2606 1748 2610 1752
rect 2614 1738 2618 1742
rect 2590 1728 2594 1732
rect 2630 1728 2634 1732
rect 2790 1838 2794 1842
rect 2750 1828 2754 1832
rect 2678 1748 2682 1752
rect 2718 1748 2722 1752
rect 2734 1748 2738 1752
rect 2654 1728 2658 1732
rect 2726 1738 2730 1742
rect 2766 1798 2770 1802
rect 2766 1748 2770 1752
rect 2702 1728 2706 1732
rect 2686 1708 2690 1712
rect 2582 1698 2586 1702
rect 2638 1698 2642 1702
rect 2622 1688 2626 1692
rect 2678 1688 2682 1692
rect 2566 1678 2570 1682
rect 2654 1678 2658 1682
rect 2694 1678 2698 1682
rect 2518 1668 2522 1672
rect 2590 1668 2594 1672
rect 2622 1668 2626 1672
rect 2630 1668 2634 1672
rect 2470 1658 2474 1662
rect 2502 1658 2506 1662
rect 2534 1658 2538 1662
rect 2614 1658 2618 1662
rect 2750 1718 2754 1722
rect 2718 1708 2722 1712
rect 2710 1668 2714 1672
rect 2558 1648 2562 1652
rect 2694 1648 2698 1652
rect 2590 1618 2594 1622
rect 2646 1618 2650 1622
rect 2622 1608 2626 1612
rect 2546 1603 2550 1607
rect 2553 1603 2557 1607
rect 2462 1598 2466 1602
rect 2494 1588 2498 1592
rect 2542 1578 2546 1582
rect 2526 1568 2530 1572
rect 2534 1558 2538 1562
rect 2454 1548 2458 1552
rect 2478 1548 2482 1552
rect 2486 1538 2490 1542
rect 2502 1538 2506 1542
rect 2518 1538 2522 1542
rect 2470 1528 2474 1532
rect 2446 1468 2450 1472
rect 2462 1468 2466 1472
rect 2502 1458 2506 1462
rect 2526 1458 2530 1462
rect 2406 1438 2410 1442
rect 2422 1438 2426 1442
rect 2246 1418 2250 1422
rect 2382 1418 2386 1422
rect 2278 1408 2282 1412
rect 2366 1408 2370 1412
rect 2294 1378 2298 1382
rect 2350 1378 2354 1382
rect 2278 1358 2282 1362
rect 2262 1348 2266 1352
rect 2142 1338 2146 1342
rect 2198 1338 2202 1342
rect 2062 1328 2066 1332
rect 2070 1328 2074 1332
rect 2030 1268 2034 1272
rect 2054 1268 2058 1272
rect 2022 1248 2026 1252
rect 2014 1188 2018 1192
rect 2038 1168 2042 1172
rect 2150 1318 2154 1322
rect 2102 1288 2106 1292
rect 2126 1288 2130 1292
rect 2142 1288 2146 1292
rect 2110 1278 2114 1282
rect 2118 1278 2122 1282
rect 2110 1268 2114 1272
rect 2102 1258 2106 1262
rect 2118 1258 2122 1262
rect 2070 1248 2074 1252
rect 2094 1238 2098 1242
rect 2134 1208 2138 1212
rect 2046 1148 2050 1152
rect 2062 1148 2066 1152
rect 2086 1138 2090 1142
rect 2102 1138 2106 1142
rect 2118 1138 2122 1142
rect 2022 1128 2026 1132
rect 2054 1128 2058 1132
rect 2110 1128 2114 1132
rect 2026 1103 2030 1107
rect 2033 1103 2037 1107
rect 2166 1278 2170 1282
rect 2190 1278 2194 1282
rect 2214 1278 2218 1282
rect 2150 1268 2154 1272
rect 2262 1328 2266 1332
rect 2262 1318 2266 1322
rect 2246 1298 2250 1302
rect 2262 1298 2266 1302
rect 2254 1278 2258 1282
rect 2214 1268 2218 1272
rect 2230 1268 2234 1272
rect 2190 1258 2194 1262
rect 2198 1258 2202 1262
rect 2238 1266 2242 1270
rect 2230 1258 2234 1262
rect 2302 1358 2306 1362
rect 2342 1358 2346 1362
rect 2318 1328 2322 1332
rect 2366 1338 2370 1342
rect 2358 1328 2362 1332
rect 2326 1318 2330 1322
rect 2286 1258 2290 1262
rect 2270 1248 2274 1252
rect 2278 1248 2282 1252
rect 2198 1238 2202 1242
rect 2222 1228 2226 1232
rect 2190 1198 2194 1202
rect 2182 1188 2186 1192
rect 2214 1188 2218 1192
rect 2166 1158 2170 1162
rect 2158 1148 2162 1152
rect 2166 1148 2170 1152
rect 2238 1208 2242 1212
rect 2342 1288 2346 1292
rect 2446 1408 2450 1412
rect 2462 1448 2466 1452
rect 2478 1448 2482 1452
rect 2454 1398 2458 1402
rect 2486 1398 2490 1402
rect 2430 1388 2434 1392
rect 2486 1388 2490 1392
rect 2390 1358 2394 1362
rect 2422 1358 2426 1362
rect 2430 1358 2434 1362
rect 2462 1358 2466 1362
rect 2398 1348 2402 1352
rect 2414 1348 2418 1352
rect 2462 1348 2466 1352
rect 2390 1338 2394 1342
rect 2406 1338 2410 1342
rect 2366 1308 2370 1312
rect 2470 1338 2474 1342
rect 2446 1328 2450 1332
rect 2438 1308 2442 1312
rect 2494 1368 2498 1372
rect 2494 1348 2498 1352
rect 2446 1288 2450 1292
rect 2582 1558 2586 1562
rect 2566 1548 2570 1552
rect 2574 1538 2578 1542
rect 2558 1468 2562 1472
rect 2518 1378 2522 1382
rect 2526 1358 2530 1362
rect 2510 1328 2514 1332
rect 2526 1328 2530 1332
rect 2510 1308 2514 1312
rect 2358 1268 2362 1272
rect 2318 1248 2322 1252
rect 2342 1248 2346 1252
rect 2302 1208 2306 1212
rect 2310 1208 2314 1212
rect 2278 1188 2282 1192
rect 2262 1158 2266 1162
rect 2270 1148 2274 1152
rect 2158 1118 2162 1122
rect 2214 1138 2218 1142
rect 2190 1108 2194 1112
rect 2134 1088 2138 1092
rect 2142 1088 2146 1092
rect 2054 1078 2058 1082
rect 2014 1068 2018 1072
rect 2094 1068 2098 1072
rect 2086 1058 2090 1062
rect 2102 1058 2106 1062
rect 1886 958 1890 962
rect 1982 958 1986 962
rect 1822 948 1826 952
rect 1846 948 1850 952
rect 1918 948 1922 952
rect 1830 938 1834 942
rect 1822 928 1826 932
rect 1838 908 1842 912
rect 1814 878 1818 882
rect 1886 928 1890 932
rect 1910 928 1914 932
rect 1942 928 1946 932
rect 1870 918 1874 922
rect 1870 898 1874 902
rect 1926 878 1930 882
rect 1854 868 1858 872
rect 1886 868 1890 872
rect 1814 848 1818 852
rect 1886 838 1890 842
rect 1966 928 1970 932
rect 1982 928 1986 932
rect 1982 918 1986 922
rect 1966 908 1970 912
rect 1958 898 1962 902
rect 1934 858 1938 862
rect 1942 858 1946 862
rect 1950 848 1954 852
rect 1910 838 1914 842
rect 1902 828 1906 832
rect 1806 778 1810 782
rect 1774 758 1778 762
rect 1790 758 1794 762
rect 1814 758 1818 762
rect 1886 798 1890 802
rect 1894 798 1898 802
rect 1830 768 1834 772
rect 1742 748 1746 752
rect 1750 748 1754 752
rect 1766 748 1770 752
rect 1822 748 1826 752
rect 1766 738 1770 742
rect 1726 728 1730 732
rect 1750 728 1754 732
rect 1734 718 1738 722
rect 1734 708 1738 712
rect 1726 698 1730 702
rect 1718 688 1722 692
rect 1742 678 1746 682
rect 1790 738 1794 742
rect 1830 738 1834 742
rect 1766 688 1770 692
rect 1854 728 1858 732
rect 1798 698 1802 702
rect 1822 698 1826 702
rect 1758 678 1762 682
rect 1782 678 1786 682
rect 1750 668 1754 672
rect 1806 688 1810 692
rect 1974 808 1978 812
rect 1966 758 1970 762
rect 1902 748 1906 752
rect 1926 748 1930 752
rect 1934 748 1938 752
rect 1974 748 1978 752
rect 1878 738 1882 742
rect 1902 708 1906 712
rect 1846 668 1850 672
rect 1854 668 1858 672
rect 1886 668 1890 672
rect 1774 658 1778 662
rect 1910 658 1914 662
rect 1718 648 1722 652
rect 1822 648 1826 652
rect 1870 648 1874 652
rect 1766 638 1770 642
rect 1758 618 1762 622
rect 1790 618 1794 622
rect 1702 578 1706 582
rect 1654 568 1658 572
rect 1702 568 1706 572
rect 1598 558 1602 562
rect 1654 558 1658 562
rect 1734 558 1738 562
rect 1582 548 1586 552
rect 1646 548 1650 552
rect 1414 528 1418 532
rect 1430 498 1434 502
rect 1414 478 1418 482
rect 1334 458 1338 462
rect 1206 448 1210 452
rect 1070 438 1074 442
rect 1110 438 1114 442
rect 1166 438 1170 442
rect 1294 438 1298 442
rect 1102 388 1106 392
rect 1134 338 1138 342
rect 1078 318 1082 322
rect 1166 428 1170 432
rect 1206 348 1210 352
rect 1318 418 1322 422
rect 1350 418 1354 422
rect 1302 408 1306 412
rect 1310 348 1314 352
rect 1230 338 1234 342
rect 1270 318 1274 322
rect 1062 288 1066 292
rect 1166 288 1170 292
rect 1262 288 1266 292
rect 1038 278 1042 282
rect 1102 278 1106 282
rect 966 268 970 272
rect 1062 268 1066 272
rect 974 258 978 262
rect 1014 258 1018 262
rect 1030 258 1034 262
rect 1046 258 1050 262
rect 966 248 970 252
rect 1038 248 1042 252
rect 982 218 986 222
rect 958 178 962 182
rect 942 168 946 172
rect 934 158 938 162
rect 950 158 954 162
rect 790 118 794 122
rect 774 108 778 112
rect 846 108 850 112
rect 838 98 842 102
rect 782 88 786 92
rect 774 78 778 82
rect 806 78 810 82
rect 878 138 882 142
rect 878 128 882 132
rect 894 108 898 112
rect 870 78 874 82
rect 742 58 746 62
rect 790 58 794 62
rect 822 58 826 62
rect 870 59 874 63
rect 974 108 978 112
rect 934 88 938 92
rect 958 88 962 92
rect 934 78 938 82
rect 958 68 962 72
rect 1054 218 1058 222
rect 1134 268 1138 272
rect 1166 268 1170 272
rect 1294 268 1298 272
rect 1310 268 1314 272
rect 1078 258 1082 262
rect 1086 258 1090 262
rect 1110 258 1114 262
rect 1230 258 1234 262
rect 1278 258 1282 262
rect 1030 178 1034 182
rect 1038 178 1042 182
rect 1070 178 1074 182
rect 998 158 1002 162
rect 1078 168 1082 172
rect 1102 248 1106 252
rect 1118 238 1122 242
rect 1230 228 1234 232
rect 1166 208 1170 212
rect 1102 168 1106 172
rect 1086 148 1090 152
rect 1102 138 1106 142
rect 1110 128 1114 132
rect 1158 128 1162 132
rect 1014 118 1018 122
rect 1002 103 1006 107
rect 1009 103 1013 107
rect 1134 118 1138 122
rect 1110 78 1114 82
rect 894 58 898 62
rect 1238 188 1242 192
rect 1174 178 1178 182
rect 1182 158 1186 162
rect 1214 158 1218 162
rect 1174 138 1178 142
rect 1366 398 1370 402
rect 1398 398 1402 402
rect 1414 358 1418 362
rect 1478 528 1482 532
rect 1486 528 1490 532
rect 1574 528 1578 532
rect 1470 508 1474 512
rect 1502 518 1506 522
rect 1486 478 1490 482
rect 1438 458 1442 462
rect 1454 458 1458 462
rect 1438 448 1442 452
rect 1510 468 1514 472
rect 1518 468 1522 472
rect 1462 428 1466 432
rect 1454 398 1458 402
rect 1446 378 1450 382
rect 1550 508 1554 512
rect 1614 538 1618 542
rect 1646 528 1650 532
rect 1614 508 1618 512
rect 1654 498 1658 502
rect 1630 488 1634 492
rect 1886 648 1890 652
rect 1878 628 1882 632
rect 1862 618 1866 622
rect 1830 598 1834 602
rect 1902 598 1906 602
rect 1790 568 1794 572
rect 1822 568 1826 572
rect 1894 568 1898 572
rect 1814 558 1818 562
rect 1910 568 1914 572
rect 1694 548 1698 552
rect 1702 548 1706 552
rect 1718 548 1722 552
rect 1774 548 1778 552
rect 1782 548 1786 552
rect 1878 548 1882 552
rect 1686 538 1690 542
rect 1670 498 1674 502
rect 1614 478 1618 482
rect 1646 478 1650 482
rect 1662 478 1666 482
rect 1638 468 1642 472
rect 1694 478 1698 482
rect 1662 468 1666 472
rect 1670 458 1674 462
rect 1686 458 1690 462
rect 1606 448 1610 452
rect 1646 448 1650 452
rect 1598 428 1602 432
rect 1542 418 1546 422
rect 1522 403 1526 407
rect 1529 403 1533 407
rect 1502 388 1506 392
rect 1526 388 1530 392
rect 1494 378 1498 382
rect 1438 338 1442 342
rect 1470 338 1474 342
rect 1326 278 1330 282
rect 1358 278 1362 282
rect 1342 258 1346 262
rect 1318 198 1322 202
rect 1206 138 1210 142
rect 1270 128 1274 132
rect 1198 108 1202 112
rect 1326 168 1330 172
rect 1374 318 1378 322
rect 1198 68 1202 72
rect 1294 58 1298 62
rect 1046 48 1050 52
rect 790 8 794 12
rect 1030 8 1034 12
rect 1390 308 1394 312
rect 1422 308 1426 312
rect 1502 328 1506 332
rect 1526 318 1530 322
rect 1670 378 1674 382
rect 1694 378 1698 382
rect 1606 368 1610 372
rect 1726 538 1730 542
rect 1734 478 1738 482
rect 1718 468 1722 472
rect 1718 458 1722 462
rect 1734 458 1738 462
rect 1710 368 1714 372
rect 1766 468 1770 472
rect 1950 688 1954 692
rect 1942 678 1946 682
rect 1934 658 1938 662
rect 2062 1048 2066 1052
rect 2038 1008 2042 1012
rect 2030 938 2034 942
rect 2026 903 2030 907
rect 2033 903 2037 907
rect 2006 888 2010 892
rect 2054 998 2058 1002
rect 2094 1038 2098 1042
rect 2102 1038 2106 1042
rect 2054 978 2058 982
rect 2158 1078 2162 1082
rect 2182 1078 2186 1082
rect 2158 1068 2162 1072
rect 2182 1068 2186 1072
rect 2126 1058 2130 1062
rect 2150 1048 2154 1052
rect 2182 1048 2186 1052
rect 2182 1038 2186 1042
rect 2174 1008 2178 1012
rect 2166 998 2170 1002
rect 2094 958 2098 962
rect 2062 928 2066 932
rect 1998 878 2002 882
rect 2046 878 2050 882
rect 1998 868 2002 872
rect 1990 828 1994 832
rect 1990 748 1994 752
rect 1982 708 1986 712
rect 2022 868 2026 872
rect 2054 866 2058 870
rect 2022 848 2026 852
rect 2046 848 2050 852
rect 2006 838 2010 842
rect 2014 768 2018 772
rect 2030 728 2034 732
rect 2102 948 2106 952
rect 2078 928 2082 932
rect 2070 838 2074 842
rect 2070 818 2074 822
rect 2126 938 2130 942
rect 2110 928 2114 932
rect 2158 948 2162 952
rect 2174 948 2178 952
rect 2206 1128 2210 1132
rect 2246 1128 2250 1132
rect 2230 1118 2234 1122
rect 2214 1078 2218 1082
rect 2206 1068 2210 1072
rect 2246 1068 2250 1072
rect 2206 1058 2210 1062
rect 2222 1058 2226 1062
rect 2206 1048 2210 1052
rect 2222 1048 2226 1052
rect 2198 1028 2202 1032
rect 2254 1058 2258 1062
rect 2310 1198 2314 1202
rect 2334 1198 2338 1202
rect 2318 1188 2322 1192
rect 2318 1178 2322 1182
rect 2326 1178 2330 1182
rect 2334 1178 2338 1182
rect 2286 1138 2290 1142
rect 2342 1158 2346 1162
rect 2350 1158 2354 1162
rect 2310 1128 2314 1132
rect 2382 1278 2386 1282
rect 2494 1278 2498 1282
rect 2374 1258 2378 1262
rect 2390 1258 2394 1262
rect 2374 1248 2378 1252
rect 2486 1268 2490 1272
rect 2518 1268 2522 1272
rect 2462 1258 2466 1262
rect 2422 1248 2426 1252
rect 2390 1228 2394 1232
rect 2446 1228 2450 1232
rect 2438 1198 2442 1202
rect 2366 1168 2370 1172
rect 2454 1218 2458 1222
rect 2462 1188 2466 1192
rect 2494 1188 2498 1192
rect 2486 1168 2490 1172
rect 2454 1158 2458 1162
rect 2390 1148 2394 1152
rect 2358 1108 2362 1112
rect 2302 1098 2306 1102
rect 2334 1098 2338 1102
rect 2350 1098 2354 1102
rect 2366 1098 2370 1102
rect 2438 1148 2442 1152
rect 2406 1138 2410 1142
rect 2414 1138 2418 1142
rect 2486 1148 2490 1152
rect 2546 1403 2550 1407
rect 2553 1403 2557 1407
rect 2574 1388 2578 1392
rect 2542 1378 2546 1382
rect 2654 1598 2658 1602
rect 2646 1558 2650 1562
rect 2670 1558 2674 1562
rect 2598 1548 2602 1552
rect 2606 1548 2610 1552
rect 2630 1548 2634 1552
rect 2662 1548 2666 1552
rect 2590 1538 2594 1542
rect 2590 1508 2594 1512
rect 2638 1538 2642 1542
rect 2670 1508 2674 1512
rect 2606 1478 2610 1482
rect 2654 1478 2658 1482
rect 2670 1478 2674 1482
rect 2606 1468 2610 1472
rect 2598 1388 2602 1392
rect 2638 1438 2642 1442
rect 2670 1448 2674 1452
rect 2686 1448 2690 1452
rect 2670 1438 2674 1442
rect 2710 1518 2714 1522
rect 2702 1458 2706 1462
rect 2630 1428 2634 1432
rect 2654 1428 2658 1432
rect 2702 1428 2706 1432
rect 2694 1418 2698 1422
rect 2646 1408 2650 1412
rect 2670 1398 2674 1402
rect 2606 1378 2610 1382
rect 2566 1328 2570 1332
rect 2590 1368 2594 1372
rect 2614 1368 2618 1372
rect 2638 1358 2642 1362
rect 2550 1268 2554 1272
rect 2534 1258 2538 1262
rect 2526 1238 2530 1242
rect 2558 1238 2562 1242
rect 2574 1238 2578 1242
rect 2518 1218 2522 1222
rect 2598 1338 2602 1342
rect 2614 1338 2618 1342
rect 2742 1708 2746 1712
rect 2758 1708 2762 1712
rect 2814 1858 2818 1862
rect 2830 1858 2834 1862
rect 2862 1858 2866 1862
rect 2886 1858 2890 1862
rect 2902 1858 2906 1862
rect 2910 1858 2914 1862
rect 2934 1858 2938 1862
rect 2950 1858 2954 1862
rect 2806 1848 2810 1852
rect 2846 1818 2850 1822
rect 2830 1808 2834 1812
rect 2814 1778 2818 1782
rect 2822 1758 2826 1762
rect 2814 1738 2818 1742
rect 3166 1968 3170 1972
rect 3030 1958 3034 1962
rect 3046 1958 3050 1962
rect 2974 1938 2978 1942
rect 2998 1928 3002 1932
rect 2974 1878 2978 1882
rect 3150 1948 3154 1952
rect 3038 1928 3042 1932
rect 3038 1918 3042 1922
rect 3050 1903 3054 1907
rect 3057 1903 3061 1907
rect 3038 1898 3042 1902
rect 3142 1938 3146 1942
rect 3222 1968 3226 1972
rect 3254 1958 3258 1962
rect 3206 1948 3210 1952
rect 3214 1948 3218 1952
rect 3230 1948 3234 1952
rect 3254 1938 3258 1942
rect 3110 1928 3114 1932
rect 3166 1928 3170 1932
rect 3118 1908 3122 1912
rect 3022 1888 3026 1892
rect 3078 1888 3082 1892
rect 3086 1888 3090 1892
rect 3038 1878 3042 1882
rect 3166 1878 3170 1882
rect 2998 1858 3002 1862
rect 3070 1848 3074 1852
rect 2918 1838 2922 1842
rect 2942 1838 2946 1842
rect 2902 1828 2906 1832
rect 2910 1808 2914 1812
rect 2854 1798 2858 1802
rect 2878 1798 2882 1802
rect 2862 1748 2866 1752
rect 2942 1828 2946 1832
rect 3166 1848 3170 1852
rect 3198 1878 3202 1882
rect 3190 1868 3194 1872
rect 3206 1858 3210 1862
rect 3182 1828 3186 1832
rect 3158 1798 3162 1802
rect 3102 1788 3106 1792
rect 3142 1788 3146 1792
rect 3190 1788 3194 1792
rect 3006 1768 3010 1772
rect 3134 1768 3138 1772
rect 2934 1758 2938 1762
rect 3158 1758 3162 1762
rect 2974 1748 2978 1752
rect 2998 1748 3002 1752
rect 3126 1748 3130 1752
rect 2910 1738 2914 1742
rect 2934 1738 2938 1742
rect 2862 1728 2866 1732
rect 2798 1718 2802 1722
rect 2854 1718 2858 1722
rect 2902 1718 2906 1722
rect 2790 1688 2794 1692
rect 2806 1698 2810 1702
rect 2782 1678 2786 1682
rect 2838 1688 2842 1692
rect 2838 1678 2842 1682
rect 2766 1658 2770 1662
rect 2790 1658 2794 1662
rect 2806 1648 2810 1652
rect 2814 1648 2818 1652
rect 2726 1618 2730 1622
rect 2734 1568 2738 1572
rect 2734 1548 2738 1552
rect 2838 1628 2842 1632
rect 2870 1708 2874 1712
rect 2894 1698 2898 1702
rect 2854 1678 2858 1682
rect 2918 1678 2922 1682
rect 2926 1668 2930 1672
rect 2934 1668 2938 1672
rect 2942 1668 2946 1672
rect 2950 1658 2954 1662
rect 2998 1718 3002 1722
rect 3022 1718 3026 1722
rect 3014 1708 3018 1712
rect 3030 1708 3034 1712
rect 2966 1698 2970 1702
rect 2974 1698 2978 1702
rect 3006 1698 3010 1702
rect 2982 1678 2986 1682
rect 2974 1658 2978 1662
rect 2886 1648 2890 1652
rect 2958 1648 2962 1652
rect 2870 1628 2874 1632
rect 3006 1648 3010 1652
rect 3014 1648 3018 1652
rect 3094 1738 3098 1742
rect 3062 1728 3066 1732
rect 3050 1703 3054 1707
rect 3057 1703 3061 1707
rect 3118 1728 3122 1732
rect 3126 1728 3130 1732
rect 3094 1678 3098 1682
rect 3022 1628 3026 1632
rect 3038 1628 3042 1632
rect 2990 1618 2994 1622
rect 3030 1618 3034 1622
rect 2774 1578 2778 1582
rect 2830 1578 2834 1582
rect 2846 1578 2850 1582
rect 2822 1568 2826 1572
rect 2750 1558 2754 1562
rect 2806 1548 2810 1552
rect 2750 1518 2754 1522
rect 2750 1478 2754 1482
rect 2638 1348 2642 1352
rect 2662 1348 2666 1352
rect 2646 1328 2650 1332
rect 2670 1328 2674 1332
rect 2678 1318 2682 1322
rect 2646 1308 2650 1312
rect 2622 1288 2626 1292
rect 2638 1288 2642 1292
rect 2614 1278 2618 1282
rect 2622 1268 2626 1272
rect 2614 1248 2618 1252
rect 2614 1238 2618 1242
rect 2670 1288 2674 1292
rect 2662 1258 2666 1262
rect 2638 1228 2642 1232
rect 2546 1203 2550 1207
rect 2553 1203 2557 1207
rect 2494 1138 2498 1142
rect 2510 1138 2514 1142
rect 2470 1128 2474 1132
rect 2502 1128 2506 1132
rect 2398 1118 2402 1122
rect 2454 1118 2458 1122
rect 2414 1108 2418 1112
rect 2438 1108 2442 1112
rect 2374 1078 2378 1082
rect 2406 1078 2410 1082
rect 2350 1068 2354 1072
rect 2246 1048 2250 1052
rect 2270 1048 2274 1052
rect 2262 1028 2266 1032
rect 2278 1028 2282 1032
rect 2230 998 2234 1002
rect 2238 998 2242 1002
rect 2214 988 2218 992
rect 2198 958 2202 962
rect 2206 958 2210 962
rect 2150 938 2154 942
rect 2174 938 2178 942
rect 2182 938 2186 942
rect 2190 938 2194 942
rect 2110 918 2114 922
rect 2134 918 2138 922
rect 2118 908 2122 912
rect 2246 968 2250 972
rect 2158 928 2162 932
rect 2230 948 2234 952
rect 2246 948 2250 952
rect 2230 928 2234 932
rect 2222 918 2226 922
rect 2206 898 2210 902
rect 2174 888 2178 892
rect 2110 878 2114 882
rect 2134 878 2138 882
rect 2198 868 2202 872
rect 2158 858 2162 862
rect 2110 848 2114 852
rect 2126 848 2130 852
rect 2102 838 2106 842
rect 2134 828 2138 832
rect 2118 798 2122 802
rect 2230 908 2234 912
rect 2222 878 2226 882
rect 2190 858 2194 862
rect 2326 1058 2330 1062
rect 2342 1058 2346 1062
rect 2390 1068 2394 1072
rect 2406 1068 2410 1072
rect 2286 1008 2290 1012
rect 2278 978 2282 982
rect 2318 1048 2322 1052
rect 2310 1008 2314 1012
rect 2294 968 2298 972
rect 2278 958 2282 962
rect 2286 958 2290 962
rect 2278 938 2282 942
rect 2254 918 2258 922
rect 2230 858 2234 862
rect 2238 858 2242 862
rect 2262 878 2266 882
rect 2318 968 2322 972
rect 2302 928 2306 932
rect 2486 1098 2490 1102
rect 2502 1078 2506 1082
rect 2558 1138 2562 1142
rect 2582 1158 2586 1162
rect 2622 1158 2626 1162
rect 2646 1148 2650 1152
rect 2606 1138 2610 1142
rect 2622 1138 2626 1142
rect 2654 1138 2658 1142
rect 2550 1118 2554 1122
rect 2566 1128 2570 1132
rect 2534 1078 2538 1082
rect 2510 1068 2514 1072
rect 2486 1058 2490 1062
rect 2382 1048 2386 1052
rect 2422 1048 2426 1052
rect 2518 1048 2522 1052
rect 2558 1048 2562 1052
rect 2478 1028 2482 1032
rect 2510 1028 2514 1032
rect 2350 998 2354 1002
rect 2398 988 2402 992
rect 2358 968 2362 972
rect 2334 938 2338 942
rect 2326 918 2330 922
rect 2294 908 2298 912
rect 2278 898 2282 902
rect 2294 878 2298 882
rect 2254 868 2258 872
rect 2270 868 2274 872
rect 2182 848 2186 852
rect 2214 848 2218 852
rect 2238 848 2242 852
rect 2198 838 2202 842
rect 2230 838 2234 842
rect 2174 808 2178 812
rect 2070 778 2074 782
rect 2158 778 2162 782
rect 2110 748 2114 752
rect 2102 738 2106 742
rect 2054 718 2058 722
rect 2026 703 2030 707
rect 2033 703 2037 707
rect 2014 688 2018 692
rect 2046 688 2050 692
rect 2014 678 2018 682
rect 2006 658 2010 662
rect 1950 648 1954 652
rect 1950 628 1954 632
rect 1926 618 1930 622
rect 2014 628 2018 632
rect 1958 598 1962 602
rect 1974 598 1978 602
rect 1990 548 1994 552
rect 1846 538 1850 542
rect 1862 538 1866 542
rect 1830 528 1834 532
rect 1854 528 1858 532
rect 1910 528 1914 532
rect 1934 528 1938 532
rect 1782 488 1786 492
rect 1854 508 1858 512
rect 1942 518 1946 522
rect 1918 508 1922 512
rect 1894 478 1898 482
rect 1790 468 1794 472
rect 1830 468 1834 472
rect 1886 468 1890 472
rect 1750 438 1754 442
rect 1806 458 1810 462
rect 1846 458 1850 462
rect 1862 458 1866 462
rect 1798 418 1802 422
rect 1822 398 1826 402
rect 1870 428 1874 432
rect 1758 388 1762 392
rect 1726 368 1730 372
rect 1766 368 1770 372
rect 1806 368 1810 372
rect 1742 358 1746 362
rect 1790 358 1794 362
rect 1870 358 1874 362
rect 1566 348 1570 352
rect 1590 348 1594 352
rect 1646 348 1650 352
rect 1702 348 1706 352
rect 1558 338 1562 342
rect 1582 328 1586 332
rect 1638 328 1642 332
rect 1662 328 1666 332
rect 1726 348 1730 352
rect 1814 348 1818 352
rect 1854 348 1858 352
rect 1734 338 1738 342
rect 1806 338 1810 342
rect 1574 318 1578 322
rect 1662 318 1666 322
rect 1694 318 1698 322
rect 1542 308 1546 312
rect 1550 298 1554 302
rect 1598 298 1602 302
rect 1654 298 1658 302
rect 1478 288 1482 292
rect 1510 288 1514 292
rect 1582 278 1586 282
rect 1390 268 1394 272
rect 1494 268 1498 272
rect 1430 218 1434 222
rect 1522 203 1526 207
rect 1529 203 1533 207
rect 1454 188 1458 192
rect 1526 188 1530 192
rect 1614 258 1618 262
rect 1694 288 1698 292
rect 1670 278 1674 282
rect 1718 278 1722 282
rect 1734 308 1738 312
rect 1758 308 1762 312
rect 1750 298 1754 302
rect 1742 288 1746 292
rect 1766 288 1770 292
rect 1782 278 1786 282
rect 1742 268 1746 272
rect 1726 258 1730 262
rect 1758 258 1762 262
rect 1782 258 1786 262
rect 1646 188 1650 192
rect 1558 138 1562 142
rect 1630 138 1634 142
rect 1398 118 1402 122
rect 1406 118 1410 122
rect 1462 108 1466 112
rect 1566 108 1570 112
rect 1590 108 1594 112
rect 1790 158 1794 162
rect 1662 148 1666 152
rect 1678 148 1682 152
rect 1694 138 1698 142
rect 1710 138 1714 142
rect 1774 128 1778 132
rect 1718 88 1722 92
rect 1614 68 1618 72
rect 1974 528 1978 532
rect 1990 528 1994 532
rect 1934 468 1938 472
rect 1894 448 1898 452
rect 1886 348 1890 352
rect 1822 338 1826 342
rect 1846 338 1850 342
rect 1878 338 1882 342
rect 1846 328 1850 332
rect 1878 328 1882 332
rect 1822 288 1826 292
rect 1870 308 1874 312
rect 1838 268 1842 272
rect 1846 268 1850 272
rect 1830 258 1834 262
rect 1814 148 1818 152
rect 1798 118 1802 122
rect 1814 68 1818 72
rect 1854 218 1858 222
rect 1934 368 1938 372
rect 1910 358 1914 362
rect 2142 748 2146 752
rect 2134 738 2138 742
rect 2150 738 2154 742
rect 2118 708 2122 712
rect 2134 708 2138 712
rect 2118 698 2122 702
rect 2086 678 2090 682
rect 2094 668 2098 672
rect 2070 658 2074 662
rect 2110 658 2114 662
rect 2062 648 2066 652
rect 2094 628 2098 632
rect 2062 618 2066 622
rect 2022 558 2026 562
rect 2006 518 2010 522
rect 1998 488 2002 492
rect 2190 768 2194 772
rect 2222 758 2226 762
rect 2174 748 2178 752
rect 2278 838 2282 842
rect 2286 838 2290 842
rect 2246 808 2250 812
rect 2262 768 2266 772
rect 2254 758 2258 762
rect 2278 748 2282 752
rect 2302 868 2306 872
rect 2310 868 2314 872
rect 2374 958 2378 962
rect 2374 948 2378 952
rect 2350 898 2354 902
rect 2390 938 2394 942
rect 2374 888 2378 892
rect 2454 1008 2458 1012
rect 2422 958 2426 962
rect 2454 958 2458 962
rect 2406 948 2410 952
rect 2422 948 2426 952
rect 2406 938 2410 942
rect 2406 918 2410 922
rect 2358 868 2362 872
rect 2374 868 2378 872
rect 2390 868 2394 872
rect 2310 838 2314 842
rect 2342 838 2346 842
rect 2318 798 2322 802
rect 2310 768 2314 772
rect 2358 848 2362 852
rect 2366 848 2370 852
rect 2374 838 2378 842
rect 2350 788 2354 792
rect 2310 748 2314 752
rect 2326 748 2330 752
rect 2182 738 2186 742
rect 2214 738 2218 742
rect 2238 738 2242 742
rect 2254 738 2258 742
rect 2166 728 2170 732
rect 2158 718 2162 722
rect 2142 658 2146 662
rect 2190 728 2194 732
rect 2214 728 2218 732
rect 2238 728 2242 732
rect 2174 718 2178 722
rect 2286 728 2290 732
rect 2302 688 2306 692
rect 2174 668 2178 672
rect 2190 668 2194 672
rect 2214 668 2218 672
rect 2270 668 2274 672
rect 2294 668 2298 672
rect 2198 658 2202 662
rect 2174 648 2178 652
rect 2158 638 2162 642
rect 2150 618 2154 622
rect 2126 608 2130 612
rect 2126 598 2130 602
rect 2086 578 2090 582
rect 2134 578 2138 582
rect 2070 558 2074 562
rect 2054 538 2058 542
rect 2046 518 2050 522
rect 2026 503 2030 507
rect 2033 503 2037 507
rect 2070 528 2074 532
rect 2078 508 2082 512
rect 2030 488 2034 492
rect 2070 488 2074 492
rect 2022 478 2026 482
rect 1966 458 1970 462
rect 1974 458 1978 462
rect 1950 448 1954 452
rect 2006 448 2010 452
rect 2006 428 2010 432
rect 1982 378 1986 382
rect 1974 358 1978 362
rect 1926 348 1930 352
rect 1926 338 1930 342
rect 1942 338 1946 342
rect 1958 338 1962 342
rect 1918 328 1922 332
rect 1910 318 1914 322
rect 1950 308 1954 312
rect 1998 368 2002 372
rect 2014 408 2018 412
rect 2062 478 2066 482
rect 2046 448 2050 452
rect 1998 348 2002 352
rect 2006 348 2010 352
rect 2078 398 2082 402
rect 2070 368 2074 372
rect 2054 358 2058 362
rect 2118 558 2122 562
rect 2102 538 2106 542
rect 2094 498 2098 502
rect 2110 478 2114 482
rect 2102 468 2106 472
rect 2118 468 2122 472
rect 2118 458 2122 462
rect 2118 418 2122 422
rect 2094 408 2098 412
rect 2190 568 2194 572
rect 2230 648 2234 652
rect 2238 618 2242 622
rect 2174 528 2178 532
rect 2158 488 2162 492
rect 2166 488 2170 492
rect 2158 458 2162 462
rect 2190 498 2194 502
rect 2182 488 2186 492
rect 2174 478 2178 482
rect 2230 538 2234 542
rect 2222 528 2226 532
rect 2214 508 2218 512
rect 2222 488 2226 492
rect 2238 488 2242 492
rect 2230 468 2234 472
rect 2174 448 2178 452
rect 2198 448 2202 452
rect 2214 448 2218 452
rect 2190 428 2194 432
rect 2190 378 2194 382
rect 2174 368 2178 372
rect 2134 358 2138 362
rect 2158 358 2162 362
rect 2014 338 2018 342
rect 2078 338 2082 342
rect 2046 308 2050 312
rect 2026 303 2030 307
rect 2033 303 2037 307
rect 2054 298 2058 302
rect 2086 298 2090 302
rect 2006 288 2010 292
rect 1910 278 1914 282
rect 1918 268 1922 272
rect 1942 268 1946 272
rect 1958 268 1962 272
rect 2022 268 2026 272
rect 2070 268 2074 272
rect 1894 258 1898 262
rect 1886 208 1890 212
rect 1926 208 1930 212
rect 1918 188 1922 192
rect 1910 168 1914 172
rect 1846 158 1850 162
rect 1854 158 1858 162
rect 1878 148 1882 152
rect 1894 128 1898 132
rect 1878 118 1882 122
rect 1830 68 1834 72
rect 1822 58 1826 62
rect 1846 58 1850 62
rect 1798 48 1802 52
rect 2102 308 2106 312
rect 2126 318 2130 322
rect 2134 318 2138 322
rect 2214 358 2218 362
rect 2278 658 2282 662
rect 2294 648 2298 652
rect 2294 628 2298 632
rect 2254 608 2258 612
rect 2262 568 2266 572
rect 2270 558 2274 562
rect 2286 558 2290 562
rect 2326 738 2330 742
rect 2350 738 2354 742
rect 2382 798 2386 802
rect 2382 788 2386 792
rect 2430 938 2434 942
rect 2454 928 2458 932
rect 2550 1038 2554 1042
rect 2566 1028 2570 1032
rect 2546 1003 2550 1007
rect 2553 1003 2557 1007
rect 2510 968 2514 972
rect 2518 958 2522 962
rect 2606 1128 2610 1132
rect 2646 1128 2650 1132
rect 2638 1118 2642 1122
rect 2662 1108 2666 1112
rect 2614 1098 2618 1102
rect 2686 1288 2690 1292
rect 2678 1278 2682 1282
rect 2686 1238 2690 1242
rect 2726 1438 2730 1442
rect 2750 1438 2754 1442
rect 2734 1378 2738 1382
rect 2766 1508 2770 1512
rect 2774 1508 2778 1512
rect 2766 1498 2770 1502
rect 2782 1438 2786 1442
rect 2774 1428 2778 1432
rect 2774 1418 2778 1422
rect 3022 1608 3026 1612
rect 3046 1608 3050 1612
rect 2902 1598 2906 1602
rect 3046 1598 3050 1602
rect 2838 1568 2842 1572
rect 2854 1568 2858 1572
rect 2926 1568 2930 1572
rect 2870 1558 2874 1562
rect 2862 1548 2866 1552
rect 2894 1548 2898 1552
rect 2918 1538 2922 1542
rect 2878 1528 2882 1532
rect 2822 1518 2826 1522
rect 2910 1518 2914 1522
rect 2878 1488 2882 1492
rect 2806 1478 2810 1482
rect 2838 1478 2842 1482
rect 2862 1478 2866 1482
rect 2902 1468 2906 1472
rect 2806 1458 2810 1462
rect 2862 1458 2866 1462
rect 2878 1458 2882 1462
rect 2806 1448 2810 1452
rect 2838 1448 2842 1452
rect 2830 1428 2834 1432
rect 2814 1418 2818 1422
rect 2790 1408 2794 1412
rect 2790 1378 2794 1382
rect 2742 1358 2746 1362
rect 2766 1358 2770 1362
rect 2750 1348 2754 1352
rect 2782 1348 2786 1352
rect 2710 1338 2714 1342
rect 2718 1338 2722 1342
rect 2702 1308 2706 1312
rect 2726 1318 2730 1322
rect 2718 1278 2722 1282
rect 2726 1268 2730 1272
rect 2774 1328 2778 1332
rect 2806 1408 2810 1412
rect 2822 1378 2826 1382
rect 2846 1428 2850 1432
rect 2862 1368 2866 1372
rect 2822 1328 2826 1332
rect 2846 1328 2850 1332
rect 2854 1328 2858 1332
rect 2814 1318 2818 1322
rect 2798 1308 2802 1312
rect 2766 1288 2770 1292
rect 2798 1288 2802 1292
rect 2742 1268 2746 1272
rect 2710 1258 2714 1262
rect 2734 1258 2738 1262
rect 2702 1248 2706 1252
rect 2750 1248 2754 1252
rect 2774 1268 2778 1272
rect 2782 1268 2786 1272
rect 2782 1248 2786 1252
rect 2814 1248 2818 1252
rect 2702 1218 2706 1222
rect 2766 1218 2770 1222
rect 2806 1218 2810 1222
rect 2694 1208 2698 1212
rect 2678 1168 2682 1172
rect 2726 1198 2730 1202
rect 2790 1198 2794 1202
rect 2782 1168 2786 1172
rect 2750 1158 2754 1162
rect 2694 1138 2698 1142
rect 2702 1108 2706 1112
rect 2670 1088 2674 1092
rect 2774 1148 2778 1152
rect 2838 1308 2842 1312
rect 2862 1308 2866 1312
rect 2950 1558 2954 1562
rect 3030 1558 3034 1562
rect 2966 1548 2970 1552
rect 3006 1548 3010 1552
rect 2942 1528 2946 1532
rect 2974 1538 2978 1542
rect 2998 1528 3002 1532
rect 2982 1488 2986 1492
rect 2990 1488 2994 1492
rect 2942 1478 2946 1482
rect 2966 1478 2970 1482
rect 2910 1458 2914 1462
rect 2894 1448 2898 1452
rect 2894 1388 2898 1392
rect 2950 1438 2954 1442
rect 2926 1378 2930 1382
rect 2950 1348 2954 1352
rect 2910 1328 2914 1332
rect 2886 1308 2890 1312
rect 2870 1298 2874 1302
rect 2870 1288 2874 1292
rect 2846 1258 2850 1262
rect 2854 1258 2858 1262
rect 2830 1238 2834 1242
rect 2846 1238 2850 1242
rect 2862 1238 2866 1242
rect 2830 1188 2834 1192
rect 2814 1168 2818 1172
rect 2822 1168 2826 1172
rect 2838 1168 2842 1172
rect 2742 1118 2746 1122
rect 2798 1108 2802 1112
rect 2782 1098 2786 1102
rect 2862 1168 2866 1172
rect 2934 1328 2938 1332
rect 2918 1298 2922 1302
rect 2990 1468 2994 1472
rect 3030 1528 3034 1532
rect 3062 1538 3066 1542
rect 3050 1503 3054 1507
rect 3057 1503 3061 1507
rect 3038 1488 3042 1492
rect 3054 1488 3058 1492
rect 3078 1668 3082 1672
rect 3102 1658 3106 1662
rect 3102 1648 3106 1652
rect 3110 1648 3114 1652
rect 3094 1628 3098 1632
rect 3086 1578 3090 1582
rect 3078 1528 3082 1532
rect 3102 1558 3106 1562
rect 3086 1518 3090 1522
rect 3070 1478 3074 1482
rect 3046 1468 3050 1472
rect 3062 1468 3066 1472
rect 3006 1448 3010 1452
rect 2974 1438 2978 1442
rect 2990 1428 2994 1432
rect 2974 1348 2978 1352
rect 3006 1348 3010 1352
rect 2950 1328 2954 1332
rect 2942 1288 2946 1292
rect 2950 1288 2954 1292
rect 2974 1298 2978 1302
rect 3006 1298 3010 1302
rect 3222 1838 3226 1842
rect 3238 1848 3242 1852
rect 3254 1828 3258 1832
rect 3230 1818 3234 1822
rect 3254 1768 3258 1772
rect 3198 1748 3202 1752
rect 3158 1738 3162 1742
rect 3190 1738 3194 1742
rect 3230 1738 3234 1742
rect 3182 1728 3186 1732
rect 3206 1728 3210 1732
rect 3142 1698 3146 1702
rect 3182 1698 3186 1702
rect 3134 1678 3138 1682
rect 3150 1658 3154 1662
rect 3166 1658 3170 1662
rect 3142 1648 3146 1652
rect 3118 1548 3122 1552
rect 3134 1548 3138 1552
rect 3150 1578 3154 1582
rect 3150 1568 3154 1572
rect 3158 1558 3162 1562
rect 3190 1678 3194 1682
rect 3198 1668 3202 1672
rect 3174 1568 3178 1572
rect 3190 1568 3194 1572
rect 3174 1548 3178 1552
rect 3110 1538 3114 1542
rect 3142 1538 3146 1542
rect 3166 1528 3170 1532
rect 3222 1708 3226 1712
rect 3230 1698 3234 1702
rect 3334 2058 3338 2062
rect 3350 2178 3354 2182
rect 3358 2148 3362 2152
rect 3382 2228 3386 2232
rect 3422 2258 3426 2262
rect 3446 2258 3450 2262
rect 3398 2248 3402 2252
rect 3430 2248 3434 2252
rect 3422 2238 3426 2242
rect 3446 2238 3450 2242
rect 3390 2208 3394 2212
rect 3478 2258 3482 2262
rect 3462 2198 3466 2202
rect 3534 2308 3538 2312
rect 3510 2288 3514 2292
rect 3494 2278 3498 2282
rect 3534 2268 3538 2272
rect 3454 2178 3458 2182
rect 3486 2178 3490 2182
rect 3382 2168 3386 2172
rect 3502 2168 3506 2172
rect 3438 2158 3442 2162
rect 3486 2158 3490 2162
rect 3382 2148 3386 2152
rect 3398 2148 3402 2152
rect 3454 2148 3458 2152
rect 3406 2138 3410 2142
rect 3422 2138 3426 2142
rect 3366 2118 3370 2122
rect 3430 2118 3434 2122
rect 3374 2108 3378 2112
rect 3398 2098 3402 2102
rect 3438 2088 3442 2092
rect 3494 2148 3498 2152
rect 3534 2248 3538 2252
rect 3518 2178 3522 2182
rect 3518 2158 3522 2162
rect 3510 2128 3514 2132
rect 3502 2118 3506 2122
rect 3494 2108 3498 2112
rect 3494 2088 3498 2092
rect 3366 2078 3370 2082
rect 3374 2068 3378 2072
rect 3518 2118 3522 2122
rect 3590 2328 3594 2332
rect 3550 2288 3554 2292
rect 3590 2288 3594 2292
rect 3582 2278 3586 2282
rect 3622 2348 3626 2352
rect 3646 2348 3650 2352
rect 3702 2348 3706 2352
rect 3606 2338 3610 2342
rect 3654 2338 3658 2342
rect 3726 2338 3730 2342
rect 3766 2338 3770 2342
rect 3622 2318 3626 2322
rect 3638 2298 3642 2302
rect 3646 2278 3650 2282
rect 3598 2268 3602 2272
rect 3686 2328 3690 2332
rect 3742 2328 3746 2332
rect 3694 2318 3698 2322
rect 3686 2308 3690 2312
rect 3702 2298 3706 2302
rect 3678 2278 3682 2282
rect 3726 2278 3730 2282
rect 3814 2348 3818 2352
rect 3830 2348 3834 2352
rect 3782 2338 3786 2342
rect 3790 2328 3794 2332
rect 3782 2318 3786 2322
rect 3774 2308 3778 2312
rect 3758 2278 3762 2282
rect 3750 2268 3754 2272
rect 3550 2258 3554 2262
rect 3662 2258 3666 2262
rect 3686 2258 3690 2262
rect 3742 2258 3746 2262
rect 3798 2298 3802 2302
rect 3990 2508 3994 2512
rect 3974 2478 3978 2482
rect 3982 2468 3986 2472
rect 3926 2448 3930 2452
rect 3958 2448 3962 2452
rect 4046 2568 4050 2572
rect 4078 2558 4082 2562
rect 4126 2658 4130 2662
rect 4206 2678 4210 2682
rect 4382 2748 4386 2752
rect 4390 2748 4394 2752
rect 4278 2738 4282 2742
rect 4302 2738 4306 2742
rect 4342 2738 4346 2742
rect 4286 2728 4290 2732
rect 4302 2728 4306 2732
rect 4318 2718 4322 2722
rect 4270 2678 4274 2682
rect 4286 2678 4290 2682
rect 4310 2678 4314 2682
rect 4246 2668 4250 2672
rect 4254 2668 4258 2672
rect 4270 2668 4274 2672
rect 4358 2708 4362 2712
rect 4358 2678 4362 2682
rect 4334 2668 4338 2672
rect 4206 2658 4210 2662
rect 4214 2658 4218 2662
rect 4326 2658 4330 2662
rect 4102 2568 4106 2572
rect 4134 2568 4138 2572
rect 4134 2558 4138 2562
rect 4166 2648 4170 2652
rect 4214 2648 4218 2652
rect 4158 2638 4162 2642
rect 4150 2598 4154 2602
rect 4062 2538 4066 2542
rect 4142 2538 4146 2542
rect 4086 2528 4090 2532
rect 4062 2518 4066 2522
rect 4030 2478 4034 2482
rect 4046 2468 4050 2472
rect 4082 2503 4086 2507
rect 4089 2503 4093 2507
rect 4134 2498 4138 2502
rect 4086 2488 4090 2492
rect 4110 2488 4114 2492
rect 4078 2468 4082 2472
rect 4118 2468 4122 2472
rect 4134 2468 4138 2472
rect 4158 2568 4162 2572
rect 4182 2638 4186 2642
rect 4174 2628 4178 2632
rect 4302 2648 4306 2652
rect 4318 2648 4322 2652
rect 4286 2578 4290 2582
rect 4302 2568 4306 2572
rect 4326 2568 4330 2572
rect 4230 2558 4234 2562
rect 4254 2558 4258 2562
rect 4278 2558 4282 2562
rect 4214 2548 4218 2552
rect 4238 2548 4242 2552
rect 4190 2538 4194 2542
rect 4182 2528 4186 2532
rect 4198 2528 4202 2532
rect 4190 2518 4194 2522
rect 4174 2498 4178 2502
rect 4166 2478 4170 2482
rect 4174 2468 4178 2472
rect 4070 2458 4074 2462
rect 4158 2458 4162 2462
rect 3974 2438 3978 2442
rect 3990 2438 3994 2442
rect 4006 2438 4010 2442
rect 3910 2398 3914 2402
rect 4006 2408 4010 2412
rect 4046 2408 4050 2412
rect 4046 2398 4050 2402
rect 3918 2388 3922 2392
rect 3878 2378 3882 2382
rect 3926 2378 3930 2382
rect 4030 2378 4034 2382
rect 3846 2358 3850 2362
rect 3870 2358 3874 2362
rect 3918 2358 3922 2362
rect 3966 2358 3970 2362
rect 3854 2348 3858 2352
rect 3822 2288 3826 2292
rect 3838 2298 3842 2302
rect 3806 2278 3810 2282
rect 3790 2268 3794 2272
rect 3814 2268 3818 2272
rect 3862 2338 3866 2342
rect 3862 2328 3866 2332
rect 3870 2308 3874 2312
rect 3942 2348 3946 2352
rect 3974 2348 3978 2352
rect 3998 2348 4002 2352
rect 4022 2348 4026 2352
rect 4062 2378 4066 2382
rect 4118 2368 4122 2372
rect 4150 2358 4154 2362
rect 3966 2338 3970 2342
rect 4006 2338 4010 2342
rect 4014 2338 4018 2342
rect 3918 2328 3922 2332
rect 3910 2298 3914 2302
rect 4150 2348 4154 2352
rect 4198 2478 4202 2482
rect 4254 2538 4258 2542
rect 4270 2538 4274 2542
rect 4374 2668 4378 2672
rect 4350 2658 4354 2662
rect 4406 2678 4410 2682
rect 4542 2868 4546 2872
rect 4558 2868 4562 2872
rect 4470 2848 4474 2852
rect 4462 2778 4466 2782
rect 4454 2758 4458 2762
rect 4582 2858 4586 2862
rect 4558 2838 4562 2842
rect 4350 2648 4354 2652
rect 4374 2648 4378 2652
rect 4398 2648 4402 2652
rect 4454 2648 4458 2652
rect 4342 2568 4346 2572
rect 4438 2568 4442 2572
rect 4310 2558 4314 2562
rect 4334 2558 4338 2562
rect 4342 2558 4346 2562
rect 4406 2558 4410 2562
rect 4318 2538 4322 2542
rect 4334 2528 4338 2532
rect 4470 2558 4474 2562
rect 4518 2558 4522 2562
rect 4534 2558 4538 2562
rect 4470 2548 4474 2552
rect 4486 2548 4490 2552
rect 4350 2538 4354 2542
rect 4438 2538 4442 2542
rect 4518 2538 4522 2542
rect 4382 2528 4386 2532
rect 4398 2528 4402 2532
rect 4414 2528 4418 2532
rect 4438 2528 4442 2532
rect 4446 2528 4450 2532
rect 4254 2508 4258 2512
rect 4278 2498 4282 2502
rect 4326 2498 4330 2502
rect 4286 2478 4290 2482
rect 4254 2468 4258 2472
rect 4342 2478 4346 2482
rect 4366 2478 4370 2482
rect 4358 2468 4362 2472
rect 4190 2458 4194 2462
rect 4214 2458 4218 2462
rect 4230 2458 4234 2462
rect 4246 2458 4250 2462
rect 4334 2458 4338 2462
rect 4342 2448 4346 2452
rect 4286 2438 4290 2442
rect 4390 2498 4394 2502
rect 4430 2478 4434 2482
rect 4462 2508 4466 2512
rect 4494 2508 4498 2512
rect 4518 2508 4522 2512
rect 4446 2478 4450 2482
rect 4486 2478 4490 2482
rect 4382 2468 4386 2472
rect 4430 2468 4434 2472
rect 4406 2458 4410 2462
rect 4414 2458 4418 2462
rect 4446 2458 4450 2462
rect 4542 2548 4546 2552
rect 4558 2518 4562 2522
rect 4558 2478 4562 2482
rect 4598 2858 4602 2862
rect 4598 2848 4602 2852
rect 4598 2768 4602 2772
rect 4582 2488 4586 2492
rect 4590 2488 4594 2492
rect 4366 2448 4370 2452
rect 4454 2448 4458 2452
rect 4486 2448 4490 2452
rect 4526 2448 4530 2452
rect 4374 2438 4378 2442
rect 4358 2418 4362 2422
rect 4318 2408 4322 2412
rect 4206 2388 4210 2392
rect 4438 2408 4442 2412
rect 4430 2378 4434 2382
rect 4214 2368 4218 2372
rect 4238 2368 4242 2372
rect 4278 2368 4282 2372
rect 4342 2368 4346 2372
rect 4190 2358 4194 2362
rect 4174 2338 4178 2342
rect 4126 2328 4130 2332
rect 4158 2328 4162 2332
rect 4166 2328 4170 2332
rect 4086 2318 4090 2322
rect 4082 2303 4086 2307
rect 4089 2303 4093 2307
rect 4190 2318 4194 2322
rect 3870 2278 3874 2282
rect 3894 2278 3898 2282
rect 3910 2278 3914 2282
rect 3966 2278 3970 2282
rect 3982 2278 3986 2282
rect 3998 2278 4002 2282
rect 4166 2278 4170 2282
rect 3910 2268 3914 2272
rect 3942 2268 3946 2272
rect 3974 2268 3978 2272
rect 4006 2268 4010 2272
rect 4094 2268 4098 2272
rect 3798 2258 3802 2262
rect 3822 2258 3826 2262
rect 3846 2258 3850 2262
rect 3558 2248 3562 2252
rect 3606 2248 3610 2252
rect 3622 2248 3626 2252
rect 3654 2248 3658 2252
rect 3894 2248 3898 2252
rect 3942 2248 3946 2252
rect 3750 2238 3754 2242
rect 3950 2238 3954 2242
rect 3638 2218 3642 2222
rect 3570 2203 3574 2207
rect 3577 2203 3581 2207
rect 3590 2178 3594 2182
rect 3542 2148 3546 2152
rect 3558 2148 3562 2152
rect 3598 2168 3602 2172
rect 3622 2158 3626 2162
rect 3606 2148 3610 2152
rect 3822 2228 3826 2232
rect 3870 2208 3874 2212
rect 3662 2168 3666 2172
rect 3766 2168 3770 2172
rect 3790 2168 3794 2172
rect 3990 2218 3994 2222
rect 3982 2188 3986 2192
rect 3974 2168 3978 2172
rect 3702 2158 3706 2162
rect 3710 2158 3714 2162
rect 3782 2158 3786 2162
rect 3814 2158 3818 2162
rect 3830 2158 3834 2162
rect 3726 2148 3730 2152
rect 3758 2148 3762 2152
rect 3798 2148 3802 2152
rect 3822 2148 3826 2152
rect 3862 2148 3866 2152
rect 3894 2148 3898 2152
rect 3926 2148 3930 2152
rect 3646 2138 3650 2142
rect 3670 2138 3674 2142
rect 3750 2138 3754 2142
rect 3814 2138 3818 2142
rect 3854 2138 3858 2142
rect 3934 2138 3938 2142
rect 4014 2248 4018 2252
rect 4134 2268 4138 2272
rect 4046 2258 4050 2262
rect 4118 2258 4122 2262
rect 4174 2258 4178 2262
rect 4046 2248 4050 2252
rect 4070 2248 4074 2252
rect 4062 2238 4066 2242
rect 4022 2228 4026 2232
rect 4030 2228 4034 2232
rect 4030 2218 4034 2222
rect 4014 2198 4018 2202
rect 4094 2248 4098 2252
rect 4118 2248 4122 2252
rect 4174 2248 4178 2252
rect 4078 2208 4082 2212
rect 4126 2238 4130 2242
rect 4150 2238 4154 2242
rect 4126 2218 4130 2222
rect 4158 2218 4162 2222
rect 4094 2198 4098 2202
rect 4054 2178 4058 2182
rect 3998 2148 4002 2152
rect 3550 2128 3554 2132
rect 3558 2128 3562 2132
rect 3678 2128 3682 2132
rect 3734 2128 3738 2132
rect 3782 2128 3786 2132
rect 3846 2128 3850 2132
rect 3542 2078 3546 2082
rect 3518 2068 3522 2072
rect 3382 2058 3386 2062
rect 3390 2058 3394 2062
rect 3406 2058 3410 2062
rect 3470 2058 3474 2062
rect 3366 2048 3370 2052
rect 3302 2018 3306 2022
rect 3326 2018 3330 2022
rect 3350 2018 3354 2022
rect 3374 1958 3378 1962
rect 3286 1948 3290 1952
rect 3294 1948 3298 1952
rect 3270 1878 3274 1882
rect 3270 1818 3274 1822
rect 3270 1758 3274 1762
rect 3318 1948 3322 1952
rect 3302 1938 3306 1942
rect 3342 1938 3346 1942
rect 3302 1918 3306 1922
rect 3310 1918 3314 1922
rect 3334 1918 3338 1922
rect 3374 1928 3378 1932
rect 3350 1898 3354 1902
rect 3438 2048 3442 2052
rect 3398 2008 3402 2012
rect 3646 2118 3650 2122
rect 3654 2118 3658 2122
rect 3622 2088 3626 2092
rect 3638 2078 3642 2082
rect 3702 2118 3706 2122
rect 3766 2118 3770 2122
rect 3694 2108 3698 2112
rect 3710 2088 3714 2092
rect 3678 2078 3682 2082
rect 3686 2078 3690 2082
rect 3814 2098 3818 2102
rect 3782 2088 3786 2092
rect 3814 2088 3818 2092
rect 3822 2078 3826 2082
rect 3846 2078 3850 2082
rect 3614 2068 3618 2072
rect 3630 2068 3634 2072
rect 3702 2068 3706 2072
rect 3718 2068 3722 2072
rect 3742 2068 3746 2072
rect 3902 2128 3906 2132
rect 3910 2128 3914 2132
rect 3966 2128 3970 2132
rect 3862 2098 3866 2102
rect 3878 2108 3882 2112
rect 3974 2098 3978 2102
rect 3870 2078 3874 2082
rect 3894 2078 3898 2082
rect 3958 2078 3962 2082
rect 3590 2058 3594 2062
rect 3654 2058 3658 2062
rect 3686 2058 3690 2062
rect 3726 2058 3730 2062
rect 3766 2058 3770 2062
rect 3494 2038 3498 2042
rect 3454 1978 3458 1982
rect 3574 2048 3578 2052
rect 3622 2048 3626 2052
rect 3630 2048 3634 2052
rect 3614 2018 3618 2022
rect 3570 2003 3574 2007
rect 3577 2003 3581 2007
rect 3614 1978 3618 1982
rect 3518 1968 3522 1972
rect 3542 1968 3546 1972
rect 3550 1968 3554 1972
rect 3558 1968 3562 1972
rect 3486 1958 3490 1962
rect 3430 1948 3434 1952
rect 3414 1938 3418 1942
rect 3390 1868 3394 1872
rect 3382 1858 3386 1862
rect 3398 1858 3402 1862
rect 3438 1938 3442 1942
rect 3470 1938 3474 1942
rect 3438 1928 3442 1932
rect 3430 1868 3434 1872
rect 3414 1858 3418 1862
rect 3286 1838 3290 1842
rect 3310 1818 3314 1822
rect 3326 1808 3330 1812
rect 3302 1788 3306 1792
rect 3350 1838 3354 1842
rect 3342 1768 3346 1772
rect 3358 1828 3362 1832
rect 3382 1798 3386 1802
rect 3542 1948 3546 1952
rect 3494 1938 3498 1942
rect 3534 1938 3538 1942
rect 3534 1928 3538 1932
rect 3462 1858 3466 1862
rect 3494 1858 3498 1862
rect 3510 1858 3514 1862
rect 3598 1948 3602 1952
rect 3550 1878 3554 1882
rect 3766 2048 3770 2052
rect 3774 2048 3778 2052
rect 3798 2048 3802 2052
rect 3774 2038 3778 2042
rect 3782 2038 3786 2042
rect 3790 2038 3794 2042
rect 3782 2028 3786 2032
rect 3774 1998 3778 2002
rect 3678 1988 3682 1992
rect 3686 1988 3690 1992
rect 3670 1978 3674 1982
rect 3654 1958 3658 1962
rect 3638 1948 3642 1952
rect 3710 1968 3714 1972
rect 3718 1968 3722 1972
rect 3718 1948 3722 1952
rect 3750 1948 3754 1952
rect 3662 1938 3666 1942
rect 3742 1938 3746 1942
rect 3758 1938 3762 1942
rect 3718 1928 3722 1932
rect 3630 1878 3634 1882
rect 3574 1868 3578 1872
rect 3582 1868 3586 1872
rect 3646 1908 3650 1912
rect 3686 1908 3690 1912
rect 3718 1908 3722 1912
rect 3758 1918 3762 1922
rect 3678 1878 3682 1882
rect 3710 1878 3714 1882
rect 3734 1878 3738 1882
rect 3750 1878 3754 1882
rect 3654 1858 3658 1862
rect 3670 1858 3674 1862
rect 3566 1848 3570 1852
rect 3414 1838 3418 1842
rect 3518 1838 3522 1842
rect 3470 1828 3474 1832
rect 3638 1848 3642 1852
rect 3598 1828 3602 1832
rect 3574 1818 3578 1822
rect 3398 1798 3402 1802
rect 3366 1788 3370 1792
rect 3358 1768 3362 1772
rect 3286 1758 3290 1762
rect 3310 1758 3314 1762
rect 3350 1758 3354 1762
rect 3278 1748 3282 1752
rect 3318 1748 3322 1752
rect 3262 1738 3266 1742
rect 3302 1738 3306 1742
rect 3334 1748 3338 1752
rect 3334 1728 3338 1732
rect 3278 1678 3282 1682
rect 3414 1758 3418 1762
rect 3446 1808 3450 1812
rect 3494 1808 3498 1812
rect 3486 1798 3490 1802
rect 3526 1798 3530 1802
rect 3446 1758 3450 1762
rect 3462 1758 3466 1762
rect 3430 1748 3434 1752
rect 3510 1758 3514 1762
rect 3502 1748 3506 1752
rect 3390 1738 3394 1742
rect 3406 1738 3410 1742
rect 3422 1738 3426 1742
rect 3470 1738 3474 1742
rect 3494 1738 3498 1742
rect 3518 1738 3522 1742
rect 3366 1728 3370 1732
rect 3382 1708 3386 1712
rect 3454 1708 3458 1712
rect 3358 1698 3362 1702
rect 3398 1698 3402 1702
rect 3422 1698 3426 1702
rect 3438 1698 3442 1702
rect 3246 1668 3250 1672
rect 3406 1678 3410 1682
rect 3398 1668 3402 1672
rect 3342 1658 3346 1662
rect 3398 1658 3402 1662
rect 3238 1628 3242 1632
rect 3214 1618 3218 1622
rect 3238 1598 3242 1602
rect 3318 1648 3322 1652
rect 3310 1638 3314 1642
rect 3326 1638 3330 1642
rect 3294 1628 3298 1632
rect 3302 1628 3306 1632
rect 3310 1618 3314 1622
rect 3270 1588 3274 1592
rect 3214 1548 3218 1552
rect 3310 1578 3314 1582
rect 3278 1558 3282 1562
rect 3302 1558 3306 1562
rect 3286 1548 3290 1552
rect 3318 1568 3322 1572
rect 3414 1638 3418 1642
rect 3358 1558 3362 1562
rect 3318 1548 3322 1552
rect 3342 1548 3346 1552
rect 3222 1538 3226 1542
rect 3246 1538 3250 1542
rect 3262 1538 3266 1542
rect 3294 1538 3298 1542
rect 3214 1518 3218 1522
rect 3142 1488 3146 1492
rect 3174 1488 3178 1492
rect 3206 1488 3210 1492
rect 3118 1478 3122 1482
rect 3094 1468 3098 1472
rect 3126 1468 3130 1472
rect 3198 1468 3202 1472
rect 3110 1458 3114 1462
rect 3094 1448 3098 1452
rect 3078 1438 3082 1442
rect 3110 1388 3114 1392
rect 3062 1378 3066 1382
rect 3142 1428 3146 1432
rect 3126 1418 3130 1422
rect 3118 1378 3122 1382
rect 3150 1398 3154 1402
rect 3190 1458 3194 1462
rect 3206 1458 3210 1462
rect 3198 1438 3202 1442
rect 3198 1388 3202 1392
rect 3166 1378 3170 1382
rect 3126 1358 3130 1362
rect 3134 1358 3138 1362
rect 3174 1358 3178 1362
rect 3038 1348 3042 1352
rect 3062 1348 3066 1352
rect 3118 1348 3122 1352
rect 3150 1348 3154 1352
rect 3182 1348 3186 1352
rect 3046 1338 3050 1342
rect 3078 1338 3082 1342
rect 3038 1308 3042 1312
rect 3050 1303 3054 1307
rect 3057 1303 3061 1307
rect 3006 1288 3010 1292
rect 2902 1268 2906 1272
rect 2958 1268 2962 1272
rect 3014 1268 3018 1272
rect 3030 1268 3034 1272
rect 2894 1258 2898 1262
rect 2910 1258 2914 1262
rect 2926 1258 2930 1262
rect 2990 1258 2994 1262
rect 3038 1258 3042 1262
rect 2894 1248 2898 1252
rect 2942 1238 2946 1242
rect 2950 1238 2954 1242
rect 2918 1228 2922 1232
rect 3062 1248 3066 1252
rect 2894 1218 2898 1222
rect 2958 1218 2962 1222
rect 2998 1238 3002 1242
rect 3030 1228 3034 1232
rect 3006 1218 3010 1222
rect 2990 1208 2994 1212
rect 2982 1198 2986 1202
rect 2910 1188 2914 1192
rect 2966 1188 2970 1192
rect 2886 1168 2890 1172
rect 2926 1158 2930 1162
rect 2958 1158 2962 1162
rect 2918 1148 2922 1152
rect 2878 1138 2882 1142
rect 2910 1138 2914 1142
rect 2902 1118 2906 1122
rect 2742 1088 2746 1092
rect 2830 1088 2834 1092
rect 2846 1088 2850 1092
rect 2886 1088 2890 1092
rect 2910 1088 2914 1092
rect 2926 1088 2930 1092
rect 2678 1078 2682 1082
rect 2710 1078 2714 1082
rect 2774 1078 2778 1082
rect 2814 1078 2818 1082
rect 2614 1068 2618 1072
rect 2582 1058 2586 1062
rect 2590 1058 2594 1062
rect 2582 968 2586 972
rect 2510 948 2514 952
rect 2550 948 2554 952
rect 2574 948 2578 952
rect 2614 1038 2618 1042
rect 2662 1068 2666 1072
rect 2686 1068 2690 1072
rect 2654 1058 2658 1062
rect 2694 1058 2698 1062
rect 2702 1058 2706 1062
rect 2646 1018 2650 1022
rect 2670 1018 2674 1022
rect 2638 1008 2642 1012
rect 2630 998 2634 1002
rect 2630 958 2634 962
rect 2654 998 2658 1002
rect 2606 948 2610 952
rect 2494 928 2498 932
rect 2438 918 2442 922
rect 2446 918 2450 922
rect 2462 918 2466 922
rect 2502 918 2506 922
rect 2470 908 2474 912
rect 2422 858 2426 862
rect 2414 838 2418 842
rect 2414 788 2418 792
rect 2430 768 2434 772
rect 2390 738 2394 742
rect 2382 708 2386 712
rect 2726 1068 2730 1072
rect 2798 1068 2802 1072
rect 2822 1068 2826 1072
rect 2718 1018 2722 1022
rect 2766 1038 2770 1042
rect 2782 1058 2786 1062
rect 2806 1058 2810 1062
rect 2814 1058 2818 1062
rect 2790 1038 2794 1042
rect 2774 1018 2778 1022
rect 2750 1008 2754 1012
rect 2710 998 2714 1002
rect 2774 998 2778 1002
rect 2678 978 2682 982
rect 2710 978 2714 982
rect 2670 958 2674 962
rect 2798 948 2802 952
rect 2678 938 2682 942
rect 2582 928 2586 932
rect 2646 928 2650 932
rect 2534 918 2538 922
rect 2542 888 2546 892
rect 2598 888 2602 892
rect 2550 878 2554 882
rect 2478 868 2482 872
rect 2510 868 2514 872
rect 2574 868 2578 872
rect 2638 868 2642 872
rect 2454 848 2458 852
rect 2494 848 2498 852
rect 2446 838 2450 842
rect 2462 838 2466 842
rect 2478 838 2482 842
rect 2534 858 2538 862
rect 2606 858 2610 862
rect 2638 858 2642 862
rect 2526 838 2530 842
rect 2518 828 2522 832
rect 2518 798 2522 802
rect 2502 778 2506 782
rect 2478 768 2482 772
rect 2422 728 2426 732
rect 2438 728 2442 732
rect 2366 688 2370 692
rect 2398 688 2402 692
rect 2422 688 2426 692
rect 2342 668 2346 672
rect 2358 668 2362 672
rect 2486 758 2490 762
rect 2622 848 2626 852
rect 2606 838 2610 842
rect 2614 838 2618 842
rect 2546 803 2550 807
rect 2553 803 2557 807
rect 2582 798 2586 802
rect 2574 778 2578 782
rect 2598 768 2602 772
rect 2558 758 2562 762
rect 2622 798 2626 802
rect 2614 788 2618 792
rect 2470 748 2474 752
rect 2550 748 2554 752
rect 2454 728 2458 732
rect 2494 728 2498 732
rect 2510 728 2514 732
rect 2454 678 2458 682
rect 2326 658 2330 662
rect 2430 658 2434 662
rect 2382 648 2386 652
rect 2454 608 2458 612
rect 2438 598 2442 602
rect 2350 578 2354 582
rect 2318 558 2322 562
rect 2342 558 2346 562
rect 2270 538 2274 542
rect 2278 518 2282 522
rect 2286 518 2290 522
rect 2254 508 2258 512
rect 2270 508 2274 512
rect 2254 458 2258 462
rect 2246 358 2250 362
rect 2182 328 2186 332
rect 2174 318 2178 322
rect 2158 308 2162 312
rect 2110 288 2114 292
rect 2142 288 2146 292
rect 2150 288 2154 292
rect 2134 268 2138 272
rect 2166 268 2170 272
rect 2190 268 2194 272
rect 1998 258 2002 262
rect 2038 258 2042 262
rect 2086 258 2090 262
rect 2094 258 2098 262
rect 2110 258 2114 262
rect 2158 258 2162 262
rect 1942 248 1946 252
rect 1958 248 1962 252
rect 1990 248 1994 252
rect 2174 248 2178 252
rect 2198 248 2202 252
rect 1982 238 1986 242
rect 2110 238 2114 242
rect 1934 198 1938 202
rect 1974 198 1978 202
rect 1942 158 1946 162
rect 1886 88 1890 92
rect 1918 78 1922 82
rect 1870 68 1874 72
rect 2046 178 2050 182
rect 2102 178 2106 182
rect 2094 158 2098 162
rect 1998 148 2002 152
rect 2062 148 2066 152
rect 1982 138 1986 142
rect 2078 138 2082 142
rect 1974 128 1978 132
rect 1950 108 1954 112
rect 1998 118 2002 122
rect 1982 78 1986 82
rect 1998 78 2002 82
rect 1910 58 1914 62
rect 2078 128 2082 132
rect 2078 108 2082 112
rect 2026 103 2030 107
rect 2033 103 2037 107
rect 2046 98 2050 102
rect 2062 88 2066 92
rect 2126 228 2130 232
rect 2214 328 2218 332
rect 2230 328 2234 332
rect 2222 298 2226 302
rect 2390 568 2394 572
rect 2430 568 2434 572
rect 2494 708 2498 712
rect 2494 688 2498 692
rect 2518 688 2522 692
rect 2510 678 2514 682
rect 2494 658 2498 662
rect 2518 658 2522 662
rect 2486 648 2490 652
rect 2470 588 2474 592
rect 2462 578 2466 582
rect 2462 568 2466 572
rect 2342 538 2346 542
rect 2374 538 2378 542
rect 2382 538 2386 542
rect 2326 508 2330 512
rect 2310 488 2314 492
rect 2278 468 2282 472
rect 2382 518 2386 522
rect 2366 488 2370 492
rect 2358 478 2362 482
rect 2382 478 2386 482
rect 2342 468 2346 472
rect 2350 468 2354 472
rect 2294 458 2298 462
rect 2262 448 2266 452
rect 2318 448 2322 452
rect 2286 378 2290 382
rect 2262 358 2266 362
rect 2254 328 2258 332
rect 2254 308 2258 312
rect 2262 298 2266 302
rect 2230 268 2234 272
rect 2262 268 2266 272
rect 2342 408 2346 412
rect 2326 398 2330 402
rect 2358 458 2362 462
rect 2382 438 2386 442
rect 2438 538 2442 542
rect 2406 528 2410 532
rect 2414 508 2418 512
rect 2406 488 2410 492
rect 2414 488 2418 492
rect 2446 518 2450 522
rect 2406 468 2410 472
rect 2414 468 2418 472
rect 2438 458 2442 462
rect 2302 368 2306 372
rect 2422 428 2426 432
rect 2470 508 2474 512
rect 2494 638 2498 642
rect 2502 558 2506 562
rect 2494 528 2498 532
rect 2478 498 2482 502
rect 2502 498 2506 502
rect 2510 498 2514 502
rect 2550 668 2554 672
rect 2590 748 2594 752
rect 2574 708 2578 712
rect 2646 768 2650 772
rect 2662 898 2666 902
rect 2662 838 2666 842
rect 2702 928 2706 932
rect 2822 968 2826 972
rect 3006 1188 3010 1192
rect 3014 1188 3018 1192
rect 3030 1188 3034 1192
rect 3110 1298 3114 1302
rect 3126 1298 3130 1302
rect 3246 1488 3250 1492
rect 3262 1498 3266 1502
rect 3238 1468 3242 1472
rect 3254 1468 3258 1472
rect 3246 1458 3250 1462
rect 3222 1438 3226 1442
rect 3326 1538 3330 1542
rect 3350 1538 3354 1542
rect 3334 1508 3338 1512
rect 3302 1468 3306 1472
rect 3318 1468 3322 1472
rect 3342 1458 3346 1462
rect 3270 1448 3274 1452
rect 3278 1448 3282 1452
rect 3286 1438 3290 1442
rect 3350 1448 3354 1452
rect 3326 1408 3330 1412
rect 3342 1408 3346 1412
rect 3262 1378 3266 1382
rect 3262 1348 3266 1352
rect 3166 1328 3170 1332
rect 3166 1318 3170 1322
rect 3206 1318 3210 1322
rect 3134 1288 3138 1292
rect 3158 1288 3162 1292
rect 3174 1288 3178 1292
rect 3190 1308 3194 1312
rect 3174 1268 3178 1272
rect 3118 1258 3122 1262
rect 3150 1258 3154 1262
rect 3094 1248 3098 1252
rect 3102 1248 3106 1252
rect 3142 1248 3146 1252
rect 3158 1248 3162 1252
rect 3174 1258 3178 1262
rect 3094 1218 3098 1222
rect 3030 1158 3034 1162
rect 3038 1158 3042 1162
rect 3150 1198 3154 1202
rect 3118 1158 3122 1162
rect 3126 1158 3130 1162
rect 3046 1148 3050 1152
rect 3174 1218 3178 1222
rect 3286 1338 3290 1342
rect 3294 1338 3298 1342
rect 3310 1328 3314 1332
rect 3230 1318 3234 1322
rect 3238 1288 3242 1292
rect 3238 1268 3242 1272
rect 3230 1238 3234 1242
rect 3222 1228 3226 1232
rect 3174 1188 3178 1192
rect 3214 1188 3218 1192
rect 2990 1138 2994 1142
rect 3014 1138 3018 1142
rect 3094 1138 3098 1142
rect 3150 1138 3154 1142
rect 2942 1118 2946 1122
rect 2974 1118 2978 1122
rect 2990 1118 2994 1122
rect 3014 1118 3018 1122
rect 3118 1128 3122 1132
rect 3086 1118 3090 1122
rect 2958 1108 2962 1112
rect 3070 1108 3074 1112
rect 2934 1078 2938 1082
rect 3050 1103 3054 1107
rect 3057 1103 3061 1107
rect 2974 1088 2978 1092
rect 3070 1088 3074 1092
rect 3110 1088 3114 1092
rect 2894 1068 2898 1072
rect 3142 1108 3146 1112
rect 3134 1098 3138 1102
rect 3006 1068 3010 1072
rect 3022 1068 3026 1072
rect 2878 1058 2882 1062
rect 2886 1058 2890 1062
rect 2926 1058 2930 1062
rect 3014 1058 3018 1062
rect 3030 1058 3034 1062
rect 3054 1058 3058 1062
rect 3126 1058 3130 1062
rect 2870 1048 2874 1052
rect 2846 1018 2850 1022
rect 2838 968 2842 972
rect 2822 948 2826 952
rect 2782 938 2786 942
rect 2694 918 2698 922
rect 2742 918 2746 922
rect 2694 908 2698 912
rect 2902 1028 2906 1032
rect 2982 1038 2986 1042
rect 2990 1038 2994 1042
rect 2950 1028 2954 1032
rect 2974 1028 2978 1032
rect 2942 1018 2946 1022
rect 2950 1018 2954 1022
rect 2934 998 2938 1002
rect 2886 988 2890 992
rect 2862 978 2866 982
rect 2878 978 2882 982
rect 2910 968 2914 972
rect 2894 958 2898 962
rect 2870 948 2874 952
rect 2886 948 2890 952
rect 2854 938 2858 942
rect 2878 938 2882 942
rect 2910 948 2914 952
rect 2902 938 2906 942
rect 2918 938 2922 942
rect 2806 928 2810 932
rect 2878 928 2882 932
rect 2894 928 2898 932
rect 2766 918 2770 922
rect 2710 888 2714 892
rect 2750 888 2754 892
rect 2686 868 2690 872
rect 2718 858 2722 862
rect 2734 858 2738 862
rect 2742 848 2746 852
rect 2702 838 2706 842
rect 2726 838 2730 842
rect 2694 808 2698 812
rect 2686 798 2690 802
rect 2654 758 2658 762
rect 2670 758 2674 762
rect 2726 808 2730 812
rect 2702 788 2706 792
rect 2838 908 2842 912
rect 2862 918 2866 922
rect 2846 888 2850 892
rect 2766 868 2770 872
rect 2798 868 2802 872
rect 2886 868 2890 872
rect 2774 858 2778 862
rect 2830 858 2834 862
rect 2814 838 2818 842
rect 2822 828 2826 832
rect 2814 818 2818 822
rect 2750 768 2754 772
rect 2782 768 2786 772
rect 2838 848 2842 852
rect 2966 968 2970 972
rect 2990 958 2994 962
rect 2998 948 3002 952
rect 2950 938 2954 942
rect 2966 938 2970 942
rect 2974 938 2978 942
rect 2998 938 3002 942
rect 2974 918 2978 922
rect 2950 868 2954 872
rect 2966 868 2970 872
rect 2862 858 2866 862
rect 2854 848 2858 852
rect 2846 778 2850 782
rect 2734 758 2738 762
rect 2806 758 2810 762
rect 2662 748 2666 752
rect 2678 748 2682 752
rect 2726 748 2730 752
rect 2782 748 2786 752
rect 2622 738 2626 742
rect 2670 738 2674 742
rect 2694 738 2698 742
rect 2710 738 2714 742
rect 2734 738 2738 742
rect 2790 738 2794 742
rect 2614 728 2618 732
rect 2606 708 2610 712
rect 2662 728 2666 732
rect 2646 708 2650 712
rect 2582 678 2586 682
rect 2622 698 2626 702
rect 2654 688 2658 692
rect 2566 658 2570 662
rect 2574 608 2578 612
rect 2546 603 2550 607
rect 2553 603 2557 607
rect 2614 638 2618 642
rect 2606 588 2610 592
rect 2694 718 2698 722
rect 2678 708 2682 712
rect 2734 698 2738 702
rect 2742 698 2746 702
rect 2686 688 2690 692
rect 2718 688 2722 692
rect 2670 678 2674 682
rect 2654 648 2658 652
rect 2662 598 2666 602
rect 2806 728 2810 732
rect 2798 708 2802 712
rect 2782 688 2786 692
rect 2822 718 2826 722
rect 2894 788 2898 792
rect 2878 768 2882 772
rect 2862 748 2866 752
rect 2870 748 2874 752
rect 2854 738 2858 742
rect 2902 758 2906 762
rect 2886 748 2890 752
rect 2894 748 2898 752
rect 2846 708 2850 712
rect 2830 688 2834 692
rect 2862 718 2866 722
rect 2854 698 2858 702
rect 2798 668 2802 672
rect 2702 658 2706 662
rect 2782 658 2786 662
rect 2662 588 2666 592
rect 2630 578 2634 582
rect 2574 558 2578 562
rect 2598 558 2602 562
rect 2646 558 2650 562
rect 2542 538 2546 542
rect 2582 538 2586 542
rect 2534 528 2538 532
rect 2574 528 2578 532
rect 2526 518 2530 522
rect 2542 518 2546 522
rect 2566 498 2570 502
rect 2454 478 2458 482
rect 2470 478 2474 482
rect 2462 468 2466 472
rect 2494 468 2498 472
rect 2510 468 2514 472
rect 2542 468 2546 472
rect 2446 378 2450 382
rect 2446 368 2450 372
rect 2598 518 2602 522
rect 2630 538 2634 542
rect 2654 538 2658 542
rect 2614 528 2618 532
rect 2638 528 2642 532
rect 2590 508 2594 512
rect 2606 508 2610 512
rect 2630 508 2634 512
rect 2606 498 2610 502
rect 2582 468 2586 472
rect 2710 648 2714 652
rect 2750 648 2754 652
rect 2782 648 2786 652
rect 2822 648 2826 652
rect 2726 638 2730 642
rect 2726 578 2730 582
rect 2702 558 2706 562
rect 2670 538 2674 542
rect 2758 568 2762 572
rect 2734 558 2738 562
rect 2774 558 2778 562
rect 2830 638 2834 642
rect 2838 598 2842 602
rect 2814 568 2818 572
rect 2822 568 2826 572
rect 2830 568 2834 572
rect 2798 548 2802 552
rect 2734 538 2738 542
rect 2774 538 2778 542
rect 2806 538 2810 542
rect 2798 528 2802 532
rect 2678 508 2682 512
rect 2662 498 2666 502
rect 2670 498 2674 502
rect 2662 488 2666 492
rect 2654 468 2658 472
rect 2702 508 2706 512
rect 2686 488 2690 492
rect 2694 488 2698 492
rect 2598 458 2602 462
rect 2710 498 2714 502
rect 2790 498 2794 502
rect 2822 498 2826 502
rect 2854 578 2858 582
rect 2926 848 2930 852
rect 2958 818 2962 822
rect 2942 808 2946 812
rect 2982 868 2986 872
rect 3014 958 3018 962
rect 3094 1048 3098 1052
rect 3070 1008 3074 1012
rect 3062 988 3066 992
rect 3054 958 3058 962
rect 3038 948 3042 952
rect 3054 938 3058 942
rect 3030 908 3034 912
rect 3050 903 3054 907
rect 3057 903 3061 907
rect 3094 1038 3098 1042
rect 3102 968 3106 972
rect 3094 958 3098 962
rect 3094 938 3098 942
rect 3102 938 3106 942
rect 3086 918 3090 922
rect 3046 888 3050 892
rect 3022 868 3026 872
rect 3038 868 3042 872
rect 3102 928 3106 932
rect 3158 1088 3162 1092
rect 3190 1158 3194 1162
rect 3334 1348 3338 1352
rect 3318 1318 3322 1322
rect 3334 1308 3338 1312
rect 3294 1288 3298 1292
rect 3278 1268 3282 1272
rect 3302 1268 3306 1272
rect 3270 1248 3274 1252
rect 3318 1248 3322 1252
rect 3318 1228 3322 1232
rect 3254 1168 3258 1172
rect 3294 1198 3298 1202
rect 3278 1188 3282 1192
rect 3270 1158 3274 1162
rect 3190 1138 3194 1142
rect 3174 1098 3178 1102
rect 3190 1098 3194 1102
rect 3174 1078 3178 1082
rect 3254 1128 3258 1132
rect 3238 1108 3242 1112
rect 3262 1108 3266 1112
rect 3390 1588 3394 1592
rect 3438 1678 3442 1682
rect 3454 1658 3458 1662
rect 3430 1638 3434 1642
rect 3438 1638 3442 1642
rect 3454 1578 3458 1582
rect 3406 1548 3410 1552
rect 3374 1508 3378 1512
rect 3430 1538 3434 1542
rect 3446 1538 3450 1542
rect 3494 1728 3498 1732
rect 3478 1718 3482 1722
rect 3518 1708 3522 1712
rect 3478 1668 3482 1672
rect 3570 1803 3574 1807
rect 3577 1803 3581 1807
rect 3550 1798 3554 1802
rect 3534 1748 3538 1752
rect 3574 1748 3578 1752
rect 3550 1738 3554 1742
rect 3542 1728 3546 1732
rect 3574 1728 3578 1732
rect 3534 1708 3538 1712
rect 3542 1678 3546 1682
rect 3598 1788 3602 1792
rect 3622 1788 3626 1792
rect 3598 1758 3602 1762
rect 3630 1758 3634 1762
rect 3606 1748 3610 1752
rect 3622 1738 3626 1742
rect 3614 1728 3618 1732
rect 3590 1698 3594 1702
rect 3734 1808 3738 1812
rect 3678 1758 3682 1762
rect 3726 1748 3730 1752
rect 3678 1738 3682 1742
rect 3646 1708 3650 1712
rect 3654 1708 3658 1712
rect 3670 1708 3674 1712
rect 3662 1678 3666 1682
rect 3630 1668 3634 1672
rect 3470 1658 3474 1662
rect 3510 1658 3514 1662
rect 3494 1648 3498 1652
rect 3502 1598 3506 1602
rect 3494 1568 3498 1572
rect 3502 1568 3506 1572
rect 3494 1548 3498 1552
rect 3470 1538 3474 1542
rect 3454 1528 3458 1532
rect 3462 1528 3466 1532
rect 3382 1488 3386 1492
rect 3398 1488 3402 1492
rect 3406 1488 3410 1492
rect 3462 1478 3466 1482
rect 3398 1458 3402 1462
rect 3414 1428 3418 1432
rect 3366 1388 3370 1392
rect 3358 1368 3362 1372
rect 3374 1378 3378 1382
rect 3382 1348 3386 1352
rect 3366 1288 3370 1292
rect 3350 1278 3354 1282
rect 3486 1498 3490 1502
rect 3446 1458 3450 1462
rect 3446 1448 3450 1452
rect 3454 1418 3458 1422
rect 3430 1398 3434 1402
rect 3438 1398 3442 1402
rect 3430 1368 3434 1372
rect 3422 1348 3426 1352
rect 3430 1318 3434 1322
rect 3398 1298 3402 1302
rect 3406 1298 3410 1302
rect 3398 1288 3402 1292
rect 3422 1288 3426 1292
rect 3446 1288 3450 1292
rect 3366 1258 3370 1262
rect 3390 1258 3394 1262
rect 3406 1258 3410 1262
rect 3366 1238 3370 1242
rect 3430 1228 3434 1232
rect 3438 1228 3442 1232
rect 3350 1198 3354 1202
rect 3398 1198 3402 1202
rect 3342 1158 3346 1162
rect 3350 1158 3354 1162
rect 3382 1158 3386 1162
rect 3414 1158 3418 1162
rect 3278 1138 3282 1142
rect 3310 1138 3314 1142
rect 3294 1128 3298 1132
rect 3198 1068 3202 1072
rect 3238 1068 3242 1072
rect 3262 1068 3266 1072
rect 3182 1058 3186 1062
rect 3150 1048 3154 1052
rect 3142 1008 3146 1012
rect 3166 1008 3170 1012
rect 3150 968 3154 972
rect 3126 958 3130 962
rect 3174 968 3178 972
rect 3206 1058 3210 1062
rect 3214 1058 3218 1062
rect 3214 1038 3218 1042
rect 3206 1008 3210 1012
rect 3198 998 3202 1002
rect 3198 968 3202 972
rect 3126 938 3130 942
rect 3158 938 3162 942
rect 3174 938 3178 942
rect 3134 868 3138 872
rect 3174 868 3178 872
rect 3102 858 3106 862
rect 3126 858 3130 862
rect 3166 858 3170 862
rect 2982 848 2986 852
rect 3070 848 3074 852
rect 3102 848 3106 852
rect 3126 848 3130 852
rect 3158 848 3162 852
rect 3206 928 3210 932
rect 3270 1058 3274 1062
rect 3270 1018 3274 1022
rect 3222 998 3226 1002
rect 3246 998 3250 1002
rect 3262 978 3266 982
rect 3278 1008 3282 1012
rect 3230 948 3234 952
rect 3246 948 3250 952
rect 3262 948 3266 952
rect 3230 938 3234 942
rect 3222 928 3226 932
rect 3238 928 3242 932
rect 3198 888 3202 892
rect 3214 888 3218 892
rect 3238 888 3242 892
rect 3214 868 3218 872
rect 3222 868 3226 872
rect 3262 938 3266 942
rect 3278 928 3282 932
rect 3342 1128 3346 1132
rect 3366 1128 3370 1132
rect 3326 1118 3330 1122
rect 3302 1108 3306 1112
rect 3406 1138 3410 1142
rect 3382 1108 3386 1112
rect 3526 1648 3530 1652
rect 3518 1548 3522 1552
rect 3570 1603 3574 1607
rect 3577 1603 3581 1607
rect 3574 1578 3578 1582
rect 3654 1658 3658 1662
rect 3654 1628 3658 1632
rect 3638 1618 3642 1622
rect 3630 1568 3634 1572
rect 3694 1718 3698 1722
rect 3782 1928 3786 1932
rect 3766 1898 3770 1902
rect 3774 1898 3778 1902
rect 3766 1878 3770 1882
rect 3750 1858 3754 1862
rect 3766 1858 3770 1862
rect 3806 1988 3810 1992
rect 3838 2038 3842 2042
rect 3886 2048 3890 2052
rect 3926 2048 3930 2052
rect 3854 1998 3858 2002
rect 3862 1998 3866 2002
rect 3838 1988 3842 1992
rect 3814 1968 3818 1972
rect 3814 1958 3818 1962
rect 3830 1958 3834 1962
rect 3950 2048 3954 2052
rect 3966 2018 3970 2022
rect 3934 1998 3938 2002
rect 3934 1958 3938 1962
rect 3838 1948 3842 1952
rect 3870 1948 3874 1952
rect 3886 1948 3890 1952
rect 3902 1948 3906 1952
rect 3926 1948 3930 1952
rect 3822 1938 3826 1942
rect 3846 1938 3850 1942
rect 3790 1908 3794 1912
rect 3798 1898 3802 1902
rect 3830 1898 3834 1902
rect 3878 1938 3882 1942
rect 3918 1938 3922 1942
rect 3934 1938 3938 1942
rect 3990 2098 3994 2102
rect 4030 2138 4034 2142
rect 4006 2098 4010 2102
rect 4134 2208 4138 2212
rect 4134 2178 4138 2182
rect 4142 2178 4146 2182
rect 4046 2148 4050 2152
rect 4062 2148 4066 2152
rect 4078 2148 4082 2152
rect 4118 2148 4122 2152
rect 4158 2148 4162 2152
rect 4054 2138 4058 2142
rect 4070 2138 4074 2142
rect 4110 2138 4114 2142
rect 4126 2138 4130 2142
rect 4062 2118 4066 2122
rect 4082 2103 4086 2107
rect 4089 2103 4093 2107
rect 4070 2098 4074 2102
rect 3998 2078 4002 2082
rect 4014 2078 4018 2082
rect 4038 2078 4042 2082
rect 4134 2118 4138 2122
rect 4214 2348 4218 2352
rect 4222 2348 4226 2352
rect 4278 2348 4282 2352
rect 4206 2308 4210 2312
rect 4246 2328 4250 2332
rect 4262 2328 4266 2332
rect 4254 2318 4258 2322
rect 4246 2308 4250 2312
rect 4318 2328 4322 2332
rect 4334 2358 4338 2362
rect 4366 2358 4370 2362
rect 4406 2358 4410 2362
rect 4494 2428 4498 2432
rect 4566 2428 4570 2432
rect 4478 2398 4482 2402
rect 4526 2388 4530 2392
rect 4518 2378 4522 2382
rect 4502 2368 4506 2372
rect 4470 2358 4474 2362
rect 4366 2348 4370 2352
rect 4302 2308 4306 2312
rect 4326 2308 4330 2312
rect 4294 2288 4298 2292
rect 4302 2278 4306 2282
rect 4262 2268 4266 2272
rect 4190 2258 4194 2262
rect 4270 2258 4274 2262
rect 4254 2248 4258 2252
rect 4198 2238 4202 2242
rect 4214 2238 4218 2242
rect 4342 2268 4346 2272
rect 4302 2258 4306 2262
rect 4310 2258 4314 2262
rect 4326 2258 4330 2262
rect 4190 2228 4194 2232
rect 4222 2228 4226 2232
rect 4286 2228 4290 2232
rect 4294 2208 4298 2212
rect 4334 2248 4338 2252
rect 4342 2248 4346 2252
rect 4326 2238 4330 2242
rect 4342 2218 4346 2222
rect 4350 2208 4354 2212
rect 4334 2188 4338 2192
rect 4182 2178 4186 2182
rect 4254 2178 4258 2182
rect 4286 2178 4290 2182
rect 4182 2148 4186 2152
rect 4206 2148 4210 2152
rect 4230 2148 4234 2152
rect 4262 2148 4266 2152
rect 4294 2148 4298 2152
rect 4310 2148 4314 2152
rect 4318 2148 4322 2152
rect 4166 2138 4170 2142
rect 4182 2138 4186 2142
rect 4214 2138 4218 2142
rect 4270 2138 4274 2142
rect 4286 2138 4290 2142
rect 4166 2128 4170 2132
rect 4182 2128 4186 2132
rect 4198 2128 4202 2132
rect 4158 2088 4162 2092
rect 4190 2098 4194 2102
rect 4046 2068 4050 2072
rect 4150 2068 4154 2072
rect 4014 2058 4018 2062
rect 4022 2038 4026 2042
rect 4030 2038 4034 2042
rect 3998 2008 4002 2012
rect 3966 1958 3970 1962
rect 3958 1948 3962 1952
rect 3934 1928 3938 1932
rect 3958 1928 3962 1932
rect 3854 1898 3858 1902
rect 3870 1898 3874 1902
rect 3918 1898 3922 1902
rect 3838 1878 3842 1882
rect 3862 1878 3866 1882
rect 3886 1878 3890 1882
rect 3918 1878 3922 1882
rect 3806 1868 3810 1872
rect 4006 1948 4010 1952
rect 3990 1928 3994 1932
rect 3958 1908 3962 1912
rect 3982 1908 3986 1912
rect 3974 1898 3978 1902
rect 3942 1878 3946 1882
rect 3966 1878 3970 1882
rect 3798 1858 3802 1862
rect 3926 1858 3930 1862
rect 3894 1848 3898 1852
rect 3942 1848 3946 1852
rect 3838 1838 3842 1842
rect 3822 1828 3826 1832
rect 3782 1808 3786 1812
rect 3806 1808 3810 1812
rect 3766 1798 3770 1802
rect 3806 1788 3810 1792
rect 3758 1758 3762 1762
rect 3766 1758 3770 1762
rect 3790 1748 3794 1752
rect 3702 1708 3706 1712
rect 3686 1678 3690 1682
rect 3702 1678 3706 1682
rect 3686 1668 3690 1672
rect 3710 1668 3714 1672
rect 3678 1658 3682 1662
rect 3670 1648 3674 1652
rect 3678 1638 3682 1642
rect 3702 1638 3706 1642
rect 3758 1728 3762 1732
rect 3766 1718 3770 1722
rect 3726 1708 3730 1712
rect 3742 1708 3746 1712
rect 3766 1698 3770 1702
rect 3846 1828 3850 1832
rect 3846 1808 3850 1812
rect 3854 1808 3858 1812
rect 3830 1748 3834 1752
rect 3838 1748 3842 1752
rect 3830 1738 3834 1742
rect 3838 1738 3842 1742
rect 3814 1698 3818 1702
rect 3782 1678 3786 1682
rect 3806 1678 3810 1682
rect 3782 1668 3786 1672
rect 3718 1658 3722 1662
rect 3718 1648 3722 1652
rect 3742 1628 3746 1632
rect 3718 1578 3722 1582
rect 3590 1548 3594 1552
rect 3606 1548 3610 1552
rect 3622 1548 3626 1552
rect 3654 1548 3658 1552
rect 3774 1548 3778 1552
rect 3782 1548 3786 1552
rect 3534 1538 3538 1542
rect 3518 1468 3522 1472
rect 3566 1538 3570 1542
rect 3622 1538 3626 1542
rect 3630 1538 3634 1542
rect 3702 1538 3706 1542
rect 3550 1528 3554 1532
rect 3646 1528 3650 1532
rect 3566 1468 3570 1472
rect 3494 1448 3498 1452
rect 3510 1448 3514 1452
rect 3470 1398 3474 1402
rect 3470 1378 3474 1382
rect 3502 1388 3506 1392
rect 3502 1358 3506 1362
rect 3462 1268 3466 1272
rect 3486 1268 3490 1272
rect 3582 1448 3586 1452
rect 3550 1418 3554 1422
rect 3570 1403 3574 1407
rect 3577 1403 3581 1407
rect 3566 1378 3570 1382
rect 3590 1378 3594 1382
rect 3670 1518 3674 1522
rect 3702 1488 3706 1492
rect 3614 1478 3618 1482
rect 3678 1478 3682 1482
rect 3630 1468 3634 1472
rect 3654 1468 3658 1472
rect 3614 1458 3618 1462
rect 3614 1418 3618 1422
rect 3534 1358 3538 1362
rect 3598 1358 3602 1362
rect 3510 1348 3514 1352
rect 3558 1348 3562 1352
rect 3526 1338 3530 1342
rect 3542 1328 3546 1332
rect 3558 1318 3562 1322
rect 3534 1308 3538 1312
rect 3534 1268 3538 1272
rect 3534 1258 3538 1262
rect 3470 1248 3474 1252
rect 3486 1248 3490 1252
rect 3510 1248 3514 1252
rect 3550 1248 3554 1252
rect 3534 1228 3538 1232
rect 3454 1198 3458 1202
rect 3462 1188 3466 1192
rect 3478 1188 3482 1192
rect 3438 1168 3442 1172
rect 3454 1158 3458 1162
rect 3470 1168 3474 1172
rect 3318 1078 3322 1082
rect 3350 1078 3354 1082
rect 3358 1078 3362 1082
rect 3398 1078 3402 1082
rect 3422 1078 3426 1082
rect 3430 1078 3434 1082
rect 3334 1068 3338 1072
rect 3454 1138 3458 1142
rect 3470 1138 3474 1142
rect 3502 1168 3506 1172
rect 3526 1158 3530 1162
rect 3534 1158 3538 1162
rect 3502 1148 3506 1152
rect 3518 1148 3522 1152
rect 3510 1138 3514 1142
rect 3478 1128 3482 1132
rect 3502 1128 3506 1132
rect 3534 1128 3538 1132
rect 3454 1078 3458 1082
rect 3310 1058 3314 1062
rect 3334 1048 3338 1052
rect 3326 1018 3330 1022
rect 3326 978 3330 982
rect 3390 1068 3394 1072
rect 3486 1068 3490 1072
rect 3382 1058 3386 1062
rect 3406 1058 3410 1062
rect 3382 1048 3386 1052
rect 3350 1018 3354 1022
rect 3374 988 3378 992
rect 3342 978 3346 982
rect 3318 968 3322 972
rect 3350 958 3354 962
rect 3358 948 3362 952
rect 3430 1038 3434 1042
rect 3446 1048 3450 1052
rect 3454 1018 3458 1022
rect 3398 978 3402 982
rect 3438 978 3442 982
rect 3470 1008 3474 1012
rect 3534 1098 3538 1102
rect 3510 1078 3514 1082
rect 3502 1058 3506 1062
rect 3518 1048 3522 1052
rect 3494 1038 3498 1042
rect 3614 1328 3618 1332
rect 3606 1318 3610 1322
rect 3590 1308 3594 1312
rect 3566 1268 3570 1272
rect 3606 1298 3610 1302
rect 3606 1278 3610 1282
rect 3606 1268 3610 1272
rect 3566 1248 3570 1252
rect 3766 1498 3770 1502
rect 3790 1508 3794 1512
rect 3750 1488 3754 1492
rect 3766 1488 3770 1492
rect 3774 1488 3778 1492
rect 3718 1468 3722 1472
rect 3734 1468 3738 1472
rect 3670 1458 3674 1462
rect 3702 1458 3706 1462
rect 3710 1458 3714 1462
rect 3726 1458 3730 1462
rect 3670 1438 3674 1442
rect 3678 1378 3682 1382
rect 3710 1378 3714 1382
rect 3726 1368 3730 1372
rect 3742 1448 3746 1452
rect 3750 1428 3754 1432
rect 3758 1368 3762 1372
rect 3630 1348 3634 1352
rect 3734 1348 3738 1352
rect 3670 1338 3674 1342
rect 3806 1508 3810 1512
rect 3798 1478 3802 1482
rect 3774 1468 3778 1472
rect 3782 1468 3786 1472
rect 3830 1708 3834 1712
rect 3862 1798 3866 1802
rect 3878 1798 3882 1802
rect 3886 1788 3890 1792
rect 3870 1748 3874 1752
rect 3998 1918 4002 1922
rect 4022 1928 4026 1932
rect 4014 1908 4018 1912
rect 4094 2038 4098 2042
rect 4054 1988 4058 1992
rect 4166 2058 4170 2062
rect 4126 2028 4130 2032
rect 4110 2018 4114 2022
rect 4102 1998 4106 2002
rect 4078 1958 4082 1962
rect 4062 1948 4066 1952
rect 4046 1938 4050 1942
rect 4078 1938 4082 1942
rect 4118 1938 4122 1942
rect 4262 2118 4266 2122
rect 4294 2118 4298 2122
rect 4254 2108 4258 2112
rect 4222 2098 4226 2102
rect 4326 2128 4330 2132
rect 4310 2108 4314 2112
rect 4262 2088 4266 2092
rect 4254 2078 4258 2082
rect 4182 2048 4186 2052
rect 4190 2048 4194 2052
rect 4238 2048 4242 2052
rect 4206 2028 4210 2032
rect 4182 2018 4186 2022
rect 4190 1988 4194 1992
rect 4422 2348 4426 2352
rect 4494 2348 4498 2352
rect 4510 2348 4514 2352
rect 4406 2338 4410 2342
rect 4542 2378 4546 2382
rect 4542 2358 4546 2362
rect 4430 2328 4434 2332
rect 4462 2328 4466 2332
rect 4478 2328 4482 2332
rect 4382 2318 4386 2322
rect 4398 2318 4402 2322
rect 4470 2318 4474 2322
rect 4374 2308 4378 2312
rect 4390 2288 4394 2292
rect 4382 2278 4386 2282
rect 4390 2248 4394 2252
rect 4374 2178 4378 2182
rect 4342 2168 4346 2172
rect 4358 2168 4362 2172
rect 4350 2138 4354 2142
rect 4382 2138 4386 2142
rect 4470 2288 4474 2292
rect 4446 2268 4450 2272
rect 4454 2268 4458 2272
rect 4406 2258 4410 2262
rect 4446 2258 4450 2262
rect 4438 2218 4442 2222
rect 4430 2208 4434 2212
rect 4430 2168 4434 2172
rect 4494 2298 4498 2302
rect 4494 2258 4498 2262
rect 4486 2238 4490 2242
rect 4502 2238 4506 2242
rect 4494 2228 4498 2232
rect 4478 2208 4482 2212
rect 4454 2198 4458 2202
rect 4478 2198 4482 2202
rect 4534 2328 4538 2332
rect 4590 2408 4594 2412
rect 4582 2358 4586 2362
rect 4574 2338 4578 2342
rect 4558 2328 4562 2332
rect 4542 2318 4546 2322
rect 4558 2318 4562 2322
rect 4526 2248 4530 2252
rect 4526 2238 4530 2242
rect 4542 2238 4546 2242
rect 4510 2158 4514 2162
rect 4438 2148 4442 2152
rect 4430 2138 4434 2142
rect 4454 2138 4458 2142
rect 4398 2128 4402 2132
rect 4430 2128 4434 2132
rect 4470 2148 4474 2152
rect 4502 2148 4506 2152
rect 4438 2118 4442 2122
rect 4446 2118 4450 2122
rect 4462 2118 4466 2122
rect 4430 2088 4434 2092
rect 4270 2078 4274 2082
rect 4310 2078 4314 2082
rect 4374 2078 4378 2082
rect 4382 2078 4386 2082
rect 4286 2048 4290 2052
rect 4342 2068 4346 2072
rect 4358 2068 4362 2072
rect 4278 2018 4282 2022
rect 4302 2018 4306 2022
rect 4206 1978 4210 1982
rect 4150 1968 4154 1972
rect 4190 1968 4194 1972
rect 4246 1968 4250 1972
rect 4294 1968 4298 1972
rect 4302 1968 4306 1972
rect 4158 1958 4162 1962
rect 4134 1948 4138 1952
rect 4190 1948 4194 1952
rect 4230 1948 4234 1952
rect 4054 1928 4058 1932
rect 4070 1928 4074 1932
rect 4150 1928 4154 1932
rect 4166 1928 4170 1932
rect 4174 1928 4178 1932
rect 4046 1918 4050 1922
rect 4038 1898 4042 1902
rect 4142 1918 4146 1922
rect 4082 1903 4086 1907
rect 4089 1903 4093 1907
rect 4006 1878 4010 1882
rect 4022 1878 4026 1882
rect 4046 1878 4050 1882
rect 4086 1878 4090 1882
rect 4118 1878 4122 1882
rect 4134 1878 4138 1882
rect 4094 1858 4098 1862
rect 3998 1848 4002 1852
rect 4014 1848 4018 1852
rect 4038 1848 4042 1852
rect 4110 1848 4114 1852
rect 3934 1808 3938 1812
rect 3902 1768 3906 1772
rect 4030 1838 4034 1842
rect 4110 1818 4114 1822
rect 4030 1808 4034 1812
rect 3974 1798 3978 1802
rect 3998 1798 4002 1802
rect 3966 1788 3970 1792
rect 3942 1778 3946 1782
rect 3910 1748 3914 1752
rect 3918 1748 3922 1752
rect 4094 1788 4098 1792
rect 4054 1768 4058 1772
rect 4006 1748 4010 1752
rect 4110 1748 4114 1752
rect 3854 1738 3858 1742
rect 3870 1738 3874 1742
rect 3982 1738 3986 1742
rect 4134 1858 4138 1862
rect 4134 1748 4138 1752
rect 3846 1718 3850 1722
rect 3878 1728 3882 1732
rect 3926 1728 3930 1732
rect 3942 1728 3946 1732
rect 4046 1728 4050 1732
rect 4046 1718 4050 1722
rect 3878 1698 3882 1702
rect 3902 1678 3906 1682
rect 3838 1658 3842 1662
rect 3870 1658 3874 1662
rect 3886 1658 3890 1662
rect 3854 1648 3858 1652
rect 3838 1638 3842 1642
rect 3798 1458 3802 1462
rect 3814 1458 3818 1462
rect 3894 1568 3898 1572
rect 3846 1538 3850 1542
rect 3862 1538 3866 1542
rect 3830 1488 3834 1492
rect 3862 1498 3866 1502
rect 3878 1488 3882 1492
rect 3846 1468 3850 1472
rect 3774 1418 3778 1422
rect 3782 1398 3786 1402
rect 3782 1368 3786 1372
rect 3750 1338 3754 1342
rect 3774 1338 3778 1342
rect 3814 1418 3818 1422
rect 3814 1408 3818 1412
rect 3838 1358 3842 1362
rect 3870 1448 3874 1452
rect 3862 1378 3866 1382
rect 3878 1358 3882 1362
rect 3830 1348 3834 1352
rect 3862 1348 3866 1352
rect 3702 1328 3706 1332
rect 3638 1318 3642 1322
rect 3630 1308 3634 1312
rect 3622 1298 3626 1302
rect 3630 1278 3634 1282
rect 3694 1318 3698 1322
rect 3718 1318 3722 1322
rect 3686 1308 3690 1312
rect 3702 1308 3706 1312
rect 3678 1298 3682 1302
rect 3758 1328 3762 1332
rect 3662 1288 3666 1292
rect 3670 1288 3674 1292
rect 3686 1288 3690 1292
rect 3718 1288 3722 1292
rect 3734 1288 3738 1292
rect 3654 1268 3658 1272
rect 3742 1278 3746 1282
rect 3646 1258 3650 1262
rect 3670 1258 3674 1262
rect 3694 1258 3698 1262
rect 3622 1218 3626 1222
rect 3622 1208 3626 1212
rect 3570 1203 3574 1207
rect 3577 1203 3581 1207
rect 3582 1158 3586 1162
rect 3590 1158 3594 1162
rect 3566 1138 3570 1142
rect 3574 1128 3578 1132
rect 3582 1118 3586 1122
rect 3566 1098 3570 1102
rect 3726 1218 3730 1222
rect 3654 1208 3658 1212
rect 3678 1208 3682 1212
rect 3654 1198 3658 1202
rect 3678 1188 3682 1192
rect 3686 1158 3690 1162
rect 3646 1148 3650 1152
rect 3630 1138 3634 1142
rect 3614 1128 3618 1132
rect 3742 1218 3746 1222
rect 3758 1258 3762 1262
rect 3750 1208 3754 1212
rect 3734 1188 3738 1192
rect 3742 1148 3746 1152
rect 3686 1138 3690 1142
rect 3710 1138 3714 1142
rect 3782 1328 3786 1332
rect 3798 1318 3802 1322
rect 3830 1318 3834 1322
rect 3798 1308 3802 1312
rect 3782 1298 3786 1302
rect 3782 1288 3786 1292
rect 3774 1278 3778 1282
rect 3854 1338 3858 1342
rect 3846 1298 3850 1302
rect 3870 1298 3874 1302
rect 3838 1288 3842 1292
rect 3798 1278 3802 1282
rect 3822 1278 3826 1282
rect 3838 1268 3842 1272
rect 3870 1268 3874 1272
rect 3774 1258 3778 1262
rect 3766 1148 3770 1152
rect 3758 1138 3762 1142
rect 3678 1128 3682 1132
rect 3686 1128 3690 1132
rect 3670 1118 3674 1122
rect 3630 1108 3634 1112
rect 3662 1108 3666 1112
rect 3590 1078 3594 1082
rect 3598 1078 3602 1082
rect 3622 1078 3626 1082
rect 3638 1078 3642 1082
rect 3542 1058 3546 1062
rect 3526 1008 3530 1012
rect 3566 1068 3570 1072
rect 3582 1058 3586 1062
rect 3590 1058 3594 1062
rect 3570 1003 3574 1007
rect 3577 1003 3581 1007
rect 3494 998 3498 1002
rect 3526 998 3530 1002
rect 3558 998 3562 1002
rect 3486 988 3490 992
rect 3454 958 3458 962
rect 3406 948 3410 952
rect 3326 938 3330 942
rect 3342 938 3346 942
rect 3374 938 3378 942
rect 3558 968 3562 972
rect 3542 958 3546 962
rect 3422 948 3426 952
rect 3526 948 3530 952
rect 3534 948 3538 952
rect 3486 938 3490 942
rect 3518 938 3522 942
rect 3270 898 3274 902
rect 3294 898 3298 902
rect 3254 888 3258 892
rect 3286 888 3290 892
rect 3390 928 3394 932
rect 3334 918 3338 922
rect 3310 898 3314 902
rect 3302 878 3306 882
rect 3294 868 3298 872
rect 3270 858 3274 862
rect 3310 858 3314 862
rect 3286 848 3290 852
rect 3150 838 3154 842
rect 3158 838 3162 842
rect 3182 838 3186 842
rect 3206 838 3210 842
rect 3230 838 3234 842
rect 3014 828 3018 832
rect 3062 828 3066 832
rect 3022 818 3026 822
rect 2974 788 2978 792
rect 2990 788 2994 792
rect 2934 758 2938 762
rect 2958 758 2962 762
rect 2926 748 2930 752
rect 2990 748 2994 752
rect 2934 738 2938 742
rect 2918 728 2922 732
rect 2894 708 2898 712
rect 2910 708 2914 712
rect 2910 688 2914 692
rect 2870 668 2874 672
rect 2886 668 2890 672
rect 2934 668 2938 672
rect 2870 618 2874 622
rect 3014 778 3018 782
rect 3054 778 3058 782
rect 3038 748 3042 752
rect 3030 738 3034 742
rect 2990 728 2994 732
rect 3006 728 3010 732
rect 2926 658 2930 662
rect 2910 608 2914 612
rect 2910 598 2914 602
rect 2902 568 2906 572
rect 2878 548 2882 552
rect 2846 538 2850 542
rect 2870 538 2874 542
rect 2902 538 2906 542
rect 2982 698 2986 702
rect 3094 788 3098 792
rect 3110 758 3114 762
rect 3118 758 3122 762
rect 3134 758 3138 762
rect 3070 738 3074 742
rect 3102 738 3106 742
rect 3054 728 3058 732
rect 3050 703 3054 707
rect 3057 703 3061 707
rect 3022 688 3026 692
rect 3030 688 3034 692
rect 3006 678 3010 682
rect 2974 668 2978 672
rect 2934 638 2938 642
rect 2942 618 2946 622
rect 2950 608 2954 612
rect 2966 558 2970 562
rect 2958 548 2962 552
rect 2902 528 2906 532
rect 2886 518 2890 522
rect 2814 488 2818 492
rect 2870 488 2874 492
rect 2630 448 2634 452
rect 2670 448 2674 452
rect 2662 438 2666 442
rect 2534 428 2538 432
rect 2542 428 2546 432
rect 2622 428 2626 432
rect 2526 418 2530 422
rect 2478 408 2482 412
rect 2326 358 2330 362
rect 2350 358 2354 362
rect 2398 358 2402 362
rect 2414 358 2418 362
rect 2462 358 2466 362
rect 2302 348 2306 352
rect 2390 348 2394 352
rect 2438 348 2442 352
rect 2390 338 2394 342
rect 2294 288 2298 292
rect 2214 258 2218 262
rect 2278 258 2282 262
rect 2294 258 2298 262
rect 2238 248 2242 252
rect 2254 238 2258 242
rect 2206 208 2210 212
rect 2246 208 2250 212
rect 2126 178 2130 182
rect 2166 178 2170 182
rect 2190 178 2194 182
rect 2150 158 2154 162
rect 2214 158 2218 162
rect 2166 148 2170 152
rect 2182 148 2186 152
rect 2198 148 2202 152
rect 2238 148 2242 152
rect 2174 138 2178 142
rect 2150 128 2154 132
rect 2134 98 2138 102
rect 2118 78 2122 82
rect 2070 58 2074 62
rect 2086 58 2090 62
rect 2006 48 2010 52
rect 2014 48 2018 52
rect 2070 48 2074 52
rect 2158 88 2162 92
rect 2182 78 2186 82
rect 2190 78 2194 82
rect 2118 58 2122 62
rect 2134 58 2138 62
rect 2150 58 2154 62
rect 2222 128 2226 132
rect 2206 118 2210 122
rect 2222 108 2226 112
rect 2214 88 2218 92
rect 2262 228 2266 232
rect 2262 188 2266 192
rect 2286 198 2290 202
rect 2270 158 2274 162
rect 2270 98 2274 102
rect 2326 318 2330 322
rect 2318 308 2322 312
rect 2414 328 2418 332
rect 2366 318 2370 322
rect 2406 318 2410 322
rect 2446 318 2450 322
rect 2374 308 2378 312
rect 2358 298 2362 302
rect 2326 288 2330 292
rect 2342 278 2346 282
rect 2358 278 2362 282
rect 2326 258 2330 262
rect 2342 258 2346 262
rect 2350 248 2354 252
rect 2310 228 2314 232
rect 2318 228 2322 232
rect 2334 228 2338 232
rect 2358 208 2362 212
rect 2294 188 2298 192
rect 2358 178 2362 182
rect 2366 168 2370 172
rect 2350 158 2354 162
rect 2390 288 2394 292
rect 2390 278 2394 282
rect 2382 258 2386 262
rect 2414 288 2418 292
rect 2470 348 2474 352
rect 2502 358 2506 362
rect 2494 348 2498 352
rect 2546 403 2550 407
rect 2553 403 2557 407
rect 2558 378 2562 382
rect 2590 378 2594 382
rect 2574 348 2578 352
rect 2590 348 2594 352
rect 2462 338 2466 342
rect 2534 338 2538 342
rect 2486 328 2490 332
rect 2454 288 2458 292
rect 2510 318 2514 322
rect 2494 288 2498 292
rect 2486 278 2490 282
rect 2414 268 2418 272
rect 2454 268 2458 272
rect 2406 258 2410 262
rect 2422 258 2426 262
rect 2446 258 2450 262
rect 2390 248 2394 252
rect 2446 248 2450 252
rect 2438 208 2442 212
rect 2470 258 2474 262
rect 2534 278 2538 282
rect 2534 268 2538 272
rect 2646 408 2650 412
rect 2630 378 2634 382
rect 2622 348 2626 352
rect 2718 478 2722 482
rect 2758 478 2762 482
rect 2774 478 2778 482
rect 2822 478 2826 482
rect 2846 478 2850 482
rect 2894 488 2898 492
rect 2918 478 2922 482
rect 2710 468 2714 472
rect 2782 468 2786 472
rect 2830 468 2834 472
rect 2838 468 2842 472
rect 2862 468 2866 472
rect 2902 468 2906 472
rect 2758 458 2762 462
rect 2886 458 2890 462
rect 2718 448 2722 452
rect 2798 448 2802 452
rect 2734 438 2738 442
rect 2702 418 2706 422
rect 2678 398 2682 402
rect 2662 378 2666 382
rect 2654 368 2658 372
rect 2662 348 2666 352
rect 2710 368 2714 372
rect 2734 368 2738 372
rect 2686 348 2690 352
rect 2702 348 2706 352
rect 2806 428 2810 432
rect 2766 418 2770 422
rect 2750 408 2754 412
rect 2830 438 2834 442
rect 2878 438 2882 442
rect 3014 668 3018 672
rect 3062 668 3066 672
rect 3110 728 3114 732
rect 3094 708 3098 712
rect 3078 678 3082 682
rect 3102 668 3106 672
rect 3006 658 3010 662
rect 3070 658 3074 662
rect 3046 648 3050 652
rect 2990 618 2994 622
rect 3022 598 3026 602
rect 3014 588 3018 592
rect 2990 578 2994 582
rect 2998 578 3002 582
rect 2990 568 2994 572
rect 2982 528 2986 532
rect 2942 518 2946 522
rect 2974 518 2978 522
rect 2942 498 2946 502
rect 2934 468 2938 472
rect 2950 478 2954 482
rect 2974 468 2978 472
rect 2942 458 2946 462
rect 2966 458 2970 462
rect 2918 408 2922 412
rect 2814 388 2818 392
rect 2766 378 2770 382
rect 2742 358 2746 362
rect 2638 338 2642 342
rect 2694 338 2698 342
rect 2726 338 2730 342
rect 2742 338 2746 342
rect 2718 318 2722 322
rect 2726 318 2730 322
rect 2614 308 2618 312
rect 2630 308 2634 312
rect 2678 308 2682 312
rect 2710 308 2714 312
rect 2606 298 2610 302
rect 2662 288 2666 292
rect 2630 278 2634 282
rect 2598 268 2602 272
rect 2638 268 2642 272
rect 2462 198 2466 202
rect 2398 188 2402 192
rect 2502 248 2506 252
rect 2526 238 2530 242
rect 2510 228 2514 232
rect 2598 258 2602 262
rect 2614 258 2618 262
rect 2662 258 2666 262
rect 2566 248 2570 252
rect 2598 248 2602 252
rect 2622 248 2626 252
rect 2582 228 2586 232
rect 2546 203 2550 207
rect 2553 203 2557 207
rect 2590 188 2594 192
rect 2478 178 2482 182
rect 2574 168 2578 172
rect 2414 158 2418 162
rect 2310 148 2314 152
rect 2382 148 2386 152
rect 2398 148 2402 152
rect 2318 138 2322 142
rect 2294 128 2298 132
rect 2326 128 2330 132
rect 2382 138 2386 142
rect 2414 138 2418 142
rect 2422 138 2426 142
rect 2366 128 2370 132
rect 2294 88 2298 92
rect 2350 78 2354 82
rect 2406 108 2410 112
rect 2438 128 2442 132
rect 2470 148 2474 152
rect 2542 148 2546 152
rect 2470 128 2474 132
rect 2486 118 2490 122
rect 2686 268 2690 272
rect 2694 268 2698 272
rect 2782 358 2786 362
rect 2814 358 2818 362
rect 2830 358 2834 362
rect 2862 358 2866 362
rect 2822 348 2826 352
rect 2798 338 2802 342
rect 2814 338 2818 342
rect 2774 288 2778 292
rect 2750 278 2754 282
rect 2774 278 2778 282
rect 2790 318 2794 322
rect 2806 318 2810 322
rect 2838 318 2842 322
rect 2742 268 2746 272
rect 2782 268 2786 272
rect 2814 308 2818 312
rect 2878 348 2882 352
rect 2910 348 2914 352
rect 2854 338 2858 342
rect 2886 338 2890 342
rect 2862 268 2866 272
rect 2870 268 2874 272
rect 2894 268 2898 272
rect 2838 258 2842 262
rect 2870 258 2874 262
rect 2886 258 2890 262
rect 2718 248 2722 252
rect 2742 248 2746 252
rect 2638 238 2642 242
rect 2670 238 2674 242
rect 2686 238 2690 242
rect 2710 238 2714 242
rect 2662 218 2666 222
rect 2638 198 2642 202
rect 2630 188 2634 192
rect 2670 188 2674 192
rect 2662 178 2666 182
rect 2734 168 2738 172
rect 2686 158 2690 162
rect 2694 158 2698 162
rect 2758 168 2762 172
rect 2766 168 2770 172
rect 2614 148 2618 152
rect 2686 148 2690 152
rect 2702 148 2706 152
rect 2726 148 2730 152
rect 2758 148 2762 152
rect 2766 148 2770 152
rect 2822 248 2826 252
rect 2886 248 2890 252
rect 2902 248 2906 252
rect 2838 238 2842 242
rect 2798 218 2802 222
rect 2798 198 2802 202
rect 2982 448 2986 452
rect 2942 438 2946 442
rect 2934 338 2938 342
rect 2974 438 2978 442
rect 3006 568 3010 572
rect 3030 588 3034 592
rect 3022 568 3026 572
rect 3022 558 3026 562
rect 3046 558 3050 562
rect 3046 548 3050 552
rect 3102 658 3106 662
rect 3134 738 3138 742
rect 3150 738 3154 742
rect 3166 808 3170 812
rect 3254 808 3258 812
rect 3238 798 3242 802
rect 3214 788 3218 792
rect 3182 758 3186 762
rect 3190 758 3194 762
rect 3182 738 3186 742
rect 3150 728 3154 732
rect 3174 728 3178 732
rect 3142 708 3146 712
rect 3142 688 3146 692
rect 3134 668 3138 672
rect 3142 658 3146 662
rect 3078 638 3082 642
rect 3078 598 3082 602
rect 3038 538 3042 542
rect 3070 538 3074 542
rect 3050 503 3054 507
rect 3057 503 3061 507
rect 3126 638 3130 642
rect 3142 598 3146 602
rect 3094 578 3098 582
rect 3126 578 3130 582
rect 3102 558 3106 562
rect 3118 548 3122 552
rect 3094 538 3098 542
rect 3126 538 3130 542
rect 3030 478 3034 482
rect 3070 478 3074 482
rect 3014 468 3018 472
rect 3030 458 3034 462
rect 2966 428 2970 432
rect 2934 278 2938 282
rect 3014 428 3018 432
rect 3110 528 3114 532
rect 3158 698 3162 702
rect 3158 688 3162 692
rect 3166 678 3170 682
rect 3206 748 3210 752
rect 3238 768 3242 772
rect 3222 758 3226 762
rect 3206 728 3210 732
rect 3222 728 3226 732
rect 3214 698 3218 702
rect 3270 798 3274 802
rect 3262 748 3266 752
rect 3294 768 3298 772
rect 3302 758 3306 762
rect 3342 898 3346 902
rect 3326 868 3330 872
rect 3318 768 3322 772
rect 3270 738 3274 742
rect 3278 738 3282 742
rect 3414 928 3418 932
rect 3422 928 3426 932
rect 3462 928 3466 932
rect 3478 928 3482 932
rect 3494 928 3498 932
rect 3614 1068 3618 1072
rect 3742 1128 3746 1132
rect 3750 1128 3754 1132
rect 3710 1118 3714 1122
rect 3694 1098 3698 1102
rect 3710 1098 3714 1102
rect 3678 1068 3682 1072
rect 3702 1068 3706 1072
rect 3654 1058 3658 1062
rect 3694 1058 3698 1062
rect 3670 1048 3674 1052
rect 3702 1038 3706 1042
rect 3662 998 3666 1002
rect 3646 968 3650 972
rect 3678 968 3682 972
rect 3702 968 3706 972
rect 3622 958 3626 962
rect 3638 958 3642 962
rect 3686 958 3690 962
rect 3622 948 3626 952
rect 3646 948 3650 952
rect 3670 948 3674 952
rect 3678 948 3682 952
rect 3542 938 3546 942
rect 3558 938 3562 942
rect 3598 938 3602 942
rect 3630 938 3634 942
rect 3582 928 3586 932
rect 3358 878 3362 882
rect 3374 878 3378 882
rect 3390 878 3394 882
rect 3350 868 3354 872
rect 3422 918 3426 922
rect 3478 898 3482 902
rect 3462 888 3466 892
rect 3454 868 3458 872
rect 3614 918 3618 922
rect 3630 918 3634 922
rect 3654 928 3658 932
rect 3646 898 3650 902
rect 3534 888 3538 892
rect 3606 888 3610 892
rect 3646 888 3650 892
rect 3534 878 3538 882
rect 3542 878 3546 882
rect 3566 878 3570 882
rect 3662 878 3666 882
rect 3734 1078 3738 1082
rect 3766 1078 3770 1082
rect 3718 1058 3722 1062
rect 3742 1048 3746 1052
rect 3758 1048 3762 1052
rect 3726 1018 3730 1022
rect 3750 1018 3754 1022
rect 3742 1008 3746 1012
rect 3734 998 3738 1002
rect 3726 968 3730 972
rect 3734 968 3738 972
rect 3734 948 3738 952
rect 3750 998 3754 1002
rect 3806 1228 3810 1232
rect 3782 1188 3786 1192
rect 3790 1188 3794 1192
rect 3806 1188 3810 1192
rect 3790 1148 3794 1152
rect 3822 1158 3826 1162
rect 3798 1138 3802 1142
rect 3782 1128 3786 1132
rect 3782 1118 3786 1122
rect 3790 1098 3794 1102
rect 3878 1258 3882 1262
rect 3846 1248 3850 1252
rect 3958 1708 3962 1712
rect 3950 1698 3954 1702
rect 3926 1668 3930 1672
rect 4094 1718 4098 1722
rect 4054 1698 4058 1702
rect 3926 1658 3930 1662
rect 3958 1658 3962 1662
rect 3966 1658 3970 1662
rect 4082 1703 4086 1707
rect 4089 1703 4093 1707
rect 4206 1898 4210 1902
rect 4198 1878 4202 1882
rect 4214 1878 4218 1882
rect 4230 1878 4234 1882
rect 4494 2138 4498 2142
rect 4478 2128 4482 2132
rect 4486 2128 4490 2132
rect 4486 2098 4490 2102
rect 4574 2298 4578 2302
rect 4566 2248 4570 2252
rect 4574 2218 4578 2222
rect 4590 2148 4594 2152
rect 4550 2118 4554 2122
rect 4510 2078 4514 2082
rect 4598 2088 4602 2092
rect 4390 2068 4394 2072
rect 4438 2068 4442 2072
rect 4470 2068 4474 2072
rect 4510 2068 4514 2072
rect 4566 2068 4570 2072
rect 4374 2058 4378 2062
rect 4350 2048 4354 2052
rect 4454 2048 4458 2052
rect 4494 2058 4498 2062
rect 4406 2028 4410 2032
rect 4462 2028 4466 2032
rect 4326 2018 4330 2022
rect 4342 2018 4346 2022
rect 4342 1978 4346 1982
rect 4398 1978 4402 1982
rect 4318 1958 4322 1962
rect 4254 1918 4258 1922
rect 4294 1918 4298 1922
rect 4246 1908 4250 1912
rect 4294 1898 4298 1902
rect 4222 1868 4226 1872
rect 4238 1868 4242 1872
rect 4246 1868 4250 1872
rect 4254 1868 4258 1872
rect 4158 1858 4162 1862
rect 4262 1858 4266 1862
rect 4270 1858 4274 1862
rect 4278 1858 4282 1862
rect 4278 1848 4282 1852
rect 4158 1838 4162 1842
rect 4166 1768 4170 1772
rect 4222 1788 4226 1792
rect 4246 1788 4250 1792
rect 4222 1778 4226 1782
rect 4206 1758 4210 1762
rect 4174 1748 4178 1752
rect 4326 1878 4330 1882
rect 4318 1848 4322 1852
rect 4286 1838 4290 1842
rect 4310 1828 4314 1832
rect 4286 1788 4290 1792
rect 4318 1778 4322 1782
rect 4310 1768 4314 1772
rect 4278 1748 4282 1752
rect 4318 1748 4322 1752
rect 4174 1738 4178 1742
rect 4190 1738 4194 1742
rect 4246 1738 4250 1742
rect 4174 1718 4178 1722
rect 4070 1668 4074 1672
rect 4094 1668 4098 1672
rect 4150 1668 4154 1672
rect 3990 1658 3994 1662
rect 4022 1658 4026 1662
rect 4046 1658 4050 1662
rect 4078 1658 4082 1662
rect 4118 1658 4122 1662
rect 3982 1648 3986 1652
rect 4014 1648 4018 1652
rect 4054 1648 4058 1652
rect 3934 1638 3938 1642
rect 3950 1638 3954 1642
rect 3982 1588 3986 1592
rect 3926 1578 3930 1582
rect 4014 1568 4018 1572
rect 3942 1548 3946 1552
rect 3974 1548 3978 1552
rect 3990 1548 3994 1552
rect 4006 1548 4010 1552
rect 4046 1548 4050 1552
rect 3950 1538 3954 1542
rect 3966 1538 3970 1542
rect 3998 1538 4002 1542
rect 3910 1528 3914 1532
rect 3942 1528 3946 1532
rect 3902 1488 3906 1492
rect 3902 1478 3906 1482
rect 3918 1488 3922 1492
rect 3910 1468 3914 1472
rect 3918 1458 3922 1462
rect 4006 1528 4010 1532
rect 4006 1518 4010 1522
rect 3998 1508 4002 1512
rect 3990 1498 3994 1502
rect 3998 1488 4002 1492
rect 4022 1478 4026 1482
rect 4038 1518 4042 1522
rect 4038 1468 4042 1472
rect 4070 1578 4074 1582
rect 4118 1618 4122 1622
rect 4134 1618 4138 1622
rect 4126 1608 4130 1612
rect 4182 1688 4186 1692
rect 4150 1648 4154 1652
rect 4198 1698 4202 1702
rect 4198 1668 4202 1672
rect 4142 1598 4146 1602
rect 4166 1578 4170 1582
rect 4102 1548 4106 1552
rect 4134 1548 4138 1552
rect 4150 1548 4154 1552
rect 4070 1528 4074 1532
rect 4150 1528 4154 1532
rect 4246 1698 4250 1702
rect 4238 1688 4242 1692
rect 4246 1658 4250 1662
rect 4206 1648 4210 1652
rect 4230 1648 4234 1652
rect 4230 1618 4234 1622
rect 4294 1738 4298 1742
rect 4286 1728 4290 1732
rect 4278 1718 4282 1722
rect 4286 1718 4290 1722
rect 4326 1708 4330 1712
rect 4390 1968 4394 1972
rect 4422 2008 4426 2012
rect 4406 1958 4410 1962
rect 4350 1948 4354 1952
rect 4406 1948 4410 1952
rect 4358 1938 4362 1942
rect 4350 1898 4354 1902
rect 4382 1918 4386 1922
rect 4374 1908 4378 1912
rect 4366 1898 4370 1902
rect 4366 1868 4370 1872
rect 4414 1938 4418 1942
rect 4406 1928 4410 1932
rect 4494 1978 4498 1982
rect 4406 1908 4410 1912
rect 4422 1908 4426 1912
rect 4446 1918 4450 1922
rect 4438 1908 4442 1912
rect 4430 1898 4434 1902
rect 4398 1888 4402 1892
rect 4494 1938 4498 1942
rect 4470 1928 4474 1932
rect 4486 1928 4490 1932
rect 4454 1878 4458 1882
rect 4462 1878 4466 1882
rect 4558 2058 4562 2062
rect 4598 2058 4602 2062
rect 4542 2038 4546 2042
rect 4550 2038 4554 2042
rect 4534 2008 4538 2012
rect 4582 2008 4586 2012
rect 4558 1948 4562 1952
rect 4526 1938 4530 1942
rect 4518 1918 4522 1922
rect 4510 1908 4514 1912
rect 4510 1898 4514 1902
rect 4486 1888 4490 1892
rect 4526 1888 4530 1892
rect 4438 1868 4442 1872
rect 4398 1858 4402 1862
rect 4414 1848 4418 1852
rect 4366 1798 4370 1802
rect 4390 1778 4394 1782
rect 4398 1758 4402 1762
rect 4358 1748 4362 1752
rect 4374 1748 4378 1752
rect 4398 1748 4402 1752
rect 4350 1738 4354 1742
rect 4374 1728 4378 1732
rect 4406 1708 4410 1712
rect 4366 1698 4370 1702
rect 4334 1688 4338 1692
rect 4310 1678 4314 1682
rect 4382 1678 4386 1682
rect 4358 1668 4362 1672
rect 4294 1638 4298 1642
rect 4254 1588 4258 1592
rect 4238 1578 4242 1582
rect 4294 1578 4298 1582
rect 4198 1568 4202 1572
rect 4222 1568 4226 1572
rect 4286 1558 4290 1562
rect 4294 1558 4298 1562
rect 4182 1548 4186 1552
rect 4198 1548 4202 1552
rect 4206 1548 4210 1552
rect 4230 1548 4234 1552
rect 4238 1548 4242 1552
rect 4062 1508 4066 1512
rect 4126 1508 4130 1512
rect 4082 1503 4086 1507
rect 4089 1503 4093 1507
rect 4182 1518 4186 1522
rect 4134 1498 4138 1502
rect 4118 1488 4122 1492
rect 4206 1498 4210 1502
rect 4062 1468 4066 1472
rect 4110 1468 4114 1472
rect 4142 1468 4146 1472
rect 4166 1468 4170 1472
rect 3942 1458 3946 1462
rect 3958 1458 3962 1462
rect 3966 1458 3970 1462
rect 4006 1458 4010 1462
rect 4022 1458 4026 1462
rect 3990 1448 3994 1452
rect 4006 1448 4010 1452
rect 3926 1388 3930 1392
rect 3942 1388 3946 1392
rect 3926 1378 3930 1382
rect 3974 1368 3978 1372
rect 3942 1348 3946 1352
rect 3998 1358 4002 1362
rect 3990 1348 3994 1352
rect 3910 1338 3914 1342
rect 3966 1338 3970 1342
rect 3950 1328 3954 1332
rect 3958 1328 3962 1332
rect 4174 1458 4178 1462
rect 4254 1518 4258 1522
rect 4366 1658 4370 1662
rect 4374 1628 4378 1632
rect 4510 1878 4514 1882
rect 4478 1868 4482 1872
rect 4494 1868 4498 1872
rect 4502 1868 4506 1872
rect 4470 1848 4474 1852
rect 4486 1848 4490 1852
rect 4462 1838 4466 1842
rect 4446 1808 4450 1812
rect 4438 1798 4442 1802
rect 4430 1778 4434 1782
rect 4422 1748 4426 1752
rect 4454 1758 4458 1762
rect 4550 1928 4554 1932
rect 4566 1938 4570 1942
rect 4566 1928 4570 1932
rect 4582 1928 4586 1932
rect 4542 1878 4546 1882
rect 4558 1878 4562 1882
rect 4542 1868 4546 1872
rect 4566 1858 4570 1862
rect 4558 1838 4562 1842
rect 4558 1828 4562 1832
rect 4534 1758 4538 1762
rect 4486 1728 4490 1732
rect 4446 1718 4450 1722
rect 4462 1698 4466 1702
rect 4414 1688 4418 1692
rect 4422 1678 4426 1682
rect 4414 1668 4418 1672
rect 4446 1668 4450 1672
rect 4518 1748 4522 1752
rect 4582 1888 4586 1892
rect 4598 1868 4602 1872
rect 4574 1758 4578 1762
rect 4542 1738 4546 1742
rect 4502 1688 4506 1692
rect 4494 1668 4498 1672
rect 4526 1668 4530 1672
rect 4590 1748 4594 1752
rect 4590 1728 4594 1732
rect 4566 1718 4570 1722
rect 4486 1658 4490 1662
rect 4550 1658 4554 1662
rect 4414 1648 4418 1652
rect 4518 1648 4522 1652
rect 4542 1638 4546 1642
rect 4366 1588 4370 1592
rect 4326 1568 4330 1572
rect 4398 1568 4402 1572
rect 4422 1558 4426 1562
rect 4510 1598 4514 1602
rect 4318 1548 4322 1552
rect 4350 1548 4354 1552
rect 4406 1548 4410 1552
rect 4446 1548 4450 1552
rect 4478 1548 4482 1552
rect 4486 1548 4490 1552
rect 4278 1538 4282 1542
rect 4294 1538 4298 1542
rect 4286 1518 4290 1522
rect 4278 1508 4282 1512
rect 4238 1488 4242 1492
rect 4262 1488 4266 1492
rect 4294 1488 4298 1492
rect 4246 1478 4250 1482
rect 4262 1478 4266 1482
rect 4238 1468 4242 1472
rect 4254 1468 4258 1472
rect 4246 1458 4250 1462
rect 4262 1458 4266 1462
rect 4126 1448 4130 1452
rect 4150 1448 4154 1452
rect 4158 1448 4162 1452
rect 4174 1438 4178 1442
rect 4190 1428 4194 1432
rect 4030 1348 4034 1352
rect 4046 1348 4050 1352
rect 4054 1348 4058 1352
rect 4014 1318 4018 1322
rect 4046 1318 4050 1322
rect 3942 1308 3946 1312
rect 3950 1308 3954 1312
rect 4038 1308 4042 1312
rect 4062 1308 4066 1312
rect 3998 1298 4002 1302
rect 3942 1278 3946 1282
rect 4014 1278 4018 1282
rect 3950 1268 3954 1272
rect 3974 1268 3978 1272
rect 4030 1268 4034 1272
rect 3918 1258 3922 1262
rect 3934 1258 3938 1262
rect 3966 1258 3970 1262
rect 3918 1248 3922 1252
rect 3966 1248 3970 1252
rect 3902 1238 3906 1242
rect 3886 1228 3890 1232
rect 3926 1218 3930 1222
rect 3862 1208 3866 1212
rect 3894 1188 3898 1192
rect 3942 1188 3946 1192
rect 3910 1158 3914 1162
rect 3846 1148 3850 1152
rect 3886 1148 3890 1152
rect 3902 1148 3906 1152
rect 3830 1128 3834 1132
rect 3798 1078 3802 1082
rect 3814 1078 3818 1082
rect 3910 1138 3914 1142
rect 3870 1128 3874 1132
rect 3894 1128 3898 1132
rect 3846 1108 3850 1112
rect 3854 1108 3858 1112
rect 3854 1088 3858 1092
rect 3878 1078 3882 1082
rect 3790 1068 3794 1072
rect 3838 1068 3842 1072
rect 3878 1068 3882 1072
rect 3774 1058 3778 1062
rect 3918 1098 3922 1102
rect 3902 1078 3906 1082
rect 3926 1078 3930 1082
rect 3918 1068 3922 1072
rect 3862 1058 3866 1062
rect 3798 1048 3802 1052
rect 3830 1048 3834 1052
rect 3838 1048 3842 1052
rect 3806 998 3810 1002
rect 3782 968 3786 972
rect 3798 968 3802 972
rect 3766 958 3770 962
rect 3758 948 3762 952
rect 3686 938 3690 942
rect 3718 938 3722 942
rect 3750 938 3754 942
rect 3782 938 3786 942
rect 3798 938 3802 942
rect 3694 918 3698 922
rect 3694 908 3698 912
rect 3918 1048 3922 1052
rect 3942 1098 3946 1102
rect 3990 1238 3994 1242
rect 4022 1238 4026 1242
rect 3974 1208 3978 1212
rect 3966 1168 3970 1172
rect 3998 1158 4002 1162
rect 4006 1158 4010 1162
rect 4062 1268 4066 1272
rect 4054 1258 4058 1262
rect 4046 1248 4050 1252
rect 4054 1248 4058 1252
rect 4182 1408 4186 1412
rect 4094 1388 4098 1392
rect 4134 1358 4138 1362
rect 4198 1398 4202 1402
rect 4190 1388 4194 1392
rect 4166 1348 4170 1352
rect 4094 1328 4098 1332
rect 4082 1303 4086 1307
rect 4089 1303 4093 1307
rect 4126 1338 4130 1342
rect 4150 1328 4154 1332
rect 4174 1328 4178 1332
rect 4134 1318 4138 1322
rect 4118 1288 4122 1292
rect 4166 1298 4170 1302
rect 4158 1278 4162 1282
rect 4086 1268 4090 1272
rect 4134 1268 4138 1272
rect 4150 1268 4154 1272
rect 4078 1258 4082 1262
rect 4110 1258 4114 1262
rect 4102 1248 4106 1252
rect 4078 1238 4082 1242
rect 4070 1208 4074 1212
rect 4046 1198 4050 1202
rect 4062 1188 4066 1192
rect 4038 1148 4042 1152
rect 4014 1138 4018 1142
rect 3966 1118 3970 1122
rect 3990 1128 3994 1132
rect 4038 1108 4042 1112
rect 4030 1098 4034 1102
rect 3990 1088 3994 1092
rect 3958 1068 3962 1072
rect 3974 1068 3978 1072
rect 4014 1068 4018 1072
rect 3958 1058 3962 1062
rect 3990 1058 3994 1062
rect 4070 1168 4074 1172
rect 4054 1078 4058 1082
rect 4062 1058 4066 1062
rect 3942 1048 3946 1052
rect 3958 1048 3962 1052
rect 4006 1048 4010 1052
rect 4046 1048 4050 1052
rect 3926 1038 3930 1042
rect 3950 1018 3954 1022
rect 3830 958 3834 962
rect 3862 958 3866 962
rect 3878 958 3882 962
rect 3910 968 3914 972
rect 3934 968 3938 972
rect 3846 948 3850 952
rect 3886 948 3890 952
rect 3902 948 3906 952
rect 3950 948 3954 952
rect 3774 928 3778 932
rect 3814 928 3818 932
rect 3750 918 3754 922
rect 3782 898 3786 902
rect 3806 898 3810 902
rect 3710 888 3714 892
rect 3750 888 3754 892
rect 3774 888 3778 892
rect 3558 868 3562 872
rect 3638 868 3642 872
rect 3678 868 3682 872
rect 3694 868 3698 872
rect 3390 848 3394 852
rect 3414 848 3418 852
rect 3350 798 3354 802
rect 3342 748 3346 752
rect 3318 738 3322 742
rect 3246 728 3250 732
rect 3270 728 3274 732
rect 3286 728 3290 732
rect 3238 708 3242 712
rect 3230 698 3234 702
rect 3294 708 3298 712
rect 3270 678 3274 682
rect 3206 668 3210 672
rect 3222 668 3226 672
rect 3286 668 3290 672
rect 3166 658 3170 662
rect 3182 658 3186 662
rect 3182 638 3186 642
rect 3262 658 3266 662
rect 3222 618 3226 622
rect 3206 608 3210 612
rect 3190 598 3194 602
rect 3222 578 3226 582
rect 3238 578 3242 582
rect 3278 638 3282 642
rect 3342 728 3346 732
rect 3334 718 3338 722
rect 3342 718 3346 722
rect 3326 708 3330 712
rect 3358 748 3362 752
rect 3414 838 3418 842
rect 3406 798 3410 802
rect 3398 788 3402 792
rect 3374 768 3378 772
rect 3366 708 3370 712
rect 3382 748 3386 752
rect 3398 748 3402 752
rect 3390 738 3394 742
rect 3358 678 3362 682
rect 3366 678 3370 682
rect 3326 668 3330 672
rect 3318 658 3322 662
rect 3350 658 3354 662
rect 3310 618 3314 622
rect 3334 618 3338 622
rect 3334 608 3338 612
rect 3326 598 3330 602
rect 3302 588 3306 592
rect 3318 578 3322 582
rect 3190 558 3194 562
rect 3206 558 3210 562
rect 3190 548 3194 552
rect 3118 488 3122 492
rect 3086 468 3090 472
rect 3062 458 3066 462
rect 3038 448 3042 452
rect 3078 398 3082 402
rect 3030 358 3034 362
rect 2974 338 2978 342
rect 2990 338 2994 342
rect 2966 308 2970 312
rect 2982 278 2986 282
rect 3006 318 3010 322
rect 3038 328 3042 332
rect 3050 303 3054 307
rect 3057 303 3061 307
rect 3094 458 3098 462
rect 3126 478 3130 482
rect 3134 468 3138 472
rect 3110 448 3114 452
rect 3134 448 3138 452
rect 3102 408 3106 412
rect 3094 348 3098 352
rect 3086 328 3090 332
rect 3086 318 3090 322
rect 3110 308 3114 312
rect 3158 418 3162 422
rect 3182 528 3186 532
rect 3206 528 3210 532
rect 3190 518 3194 522
rect 3182 508 3186 512
rect 3270 558 3274 562
rect 3246 548 3250 552
rect 3270 548 3274 552
rect 3230 538 3234 542
rect 3254 538 3258 542
rect 3230 478 3234 482
rect 3246 478 3250 482
rect 3254 478 3258 482
rect 3174 468 3178 472
rect 3190 448 3194 452
rect 3166 408 3170 412
rect 3182 398 3186 402
rect 3150 378 3154 382
rect 3158 378 3162 382
rect 3142 358 3146 362
rect 3158 368 3162 372
rect 3198 418 3202 422
rect 3198 398 3202 402
rect 3198 378 3202 382
rect 3166 348 3170 352
rect 3150 328 3154 332
rect 3134 318 3138 322
rect 3134 298 3138 302
rect 3102 288 3106 292
rect 3038 278 3042 282
rect 3078 278 3082 282
rect 2942 268 2946 272
rect 3030 268 3034 272
rect 3086 268 3090 272
rect 2934 258 2938 262
rect 2926 248 2930 252
rect 2910 238 2914 242
rect 2934 218 2938 222
rect 2862 198 2866 202
rect 2886 188 2890 192
rect 2854 178 2858 182
rect 2790 158 2794 162
rect 2790 148 2794 152
rect 2846 148 2850 152
rect 2710 138 2714 142
rect 2774 138 2778 142
rect 2806 138 2810 142
rect 2590 128 2594 132
rect 2614 128 2618 132
rect 2638 128 2642 132
rect 2718 128 2722 132
rect 2518 118 2522 122
rect 2558 118 2562 122
rect 2598 118 2602 122
rect 2422 108 2426 112
rect 2454 108 2458 112
rect 2494 108 2498 112
rect 2574 108 2578 112
rect 2638 118 2642 122
rect 2638 98 2642 102
rect 2694 98 2698 102
rect 2430 88 2434 92
rect 2470 88 2474 92
rect 2630 88 2634 92
rect 2390 78 2394 82
rect 2502 78 2506 82
rect 2534 78 2538 82
rect 2622 78 2626 82
rect 2366 68 2370 72
rect 2406 68 2410 72
rect 2422 68 2426 72
rect 2526 68 2530 72
rect 2574 68 2578 72
rect 2590 68 2594 72
rect 2198 58 2202 62
rect 2238 58 2242 62
rect 2310 58 2314 62
rect 2326 58 2330 62
rect 2142 48 2146 52
rect 2190 48 2194 52
rect 2246 48 2250 52
rect 2254 48 2258 52
rect 2334 48 2338 52
rect 2454 48 2458 52
rect 2038 38 2042 42
rect 2102 38 2106 42
rect 2486 38 2490 42
rect 2734 98 2738 102
rect 2662 88 2666 92
rect 2646 78 2650 82
rect 2670 78 2674 82
rect 2678 78 2682 82
rect 2766 78 2770 82
rect 2878 168 2882 172
rect 2926 168 2930 172
rect 2918 158 2922 162
rect 2862 148 2866 152
rect 2950 248 2954 252
rect 2966 238 2970 242
rect 2982 188 2986 192
rect 2958 168 2962 172
rect 2974 168 2978 172
rect 2942 148 2946 152
rect 3118 268 3122 272
rect 2998 248 3002 252
rect 3014 238 3018 242
rect 2990 158 2994 162
rect 3022 198 3026 202
rect 3054 228 3058 232
rect 3118 228 3122 232
rect 3022 158 3026 162
rect 3086 218 3090 222
rect 3062 198 3066 202
rect 3126 198 3130 202
rect 3078 188 3082 192
rect 3190 298 3194 302
rect 3222 448 3226 452
rect 3302 548 3306 552
rect 3318 538 3322 542
rect 3294 518 3298 522
rect 3294 488 3298 492
rect 3318 478 3322 482
rect 3294 468 3298 472
rect 3254 458 3258 462
rect 3270 458 3274 462
rect 3302 458 3306 462
rect 3262 448 3266 452
rect 3302 448 3306 452
rect 3230 438 3234 442
rect 3238 408 3242 412
rect 3382 658 3386 662
rect 3374 568 3378 572
rect 3350 528 3354 532
rect 3502 848 3506 852
rect 3430 828 3434 832
rect 3438 818 3442 822
rect 3494 818 3498 822
rect 3422 758 3426 762
rect 3430 758 3434 762
rect 3462 758 3466 762
rect 3510 808 3514 812
rect 3550 828 3554 832
rect 3550 818 3554 822
rect 3542 798 3546 802
rect 3518 788 3522 792
rect 3510 748 3514 752
rect 3422 738 3426 742
rect 3438 738 3442 742
rect 3462 738 3466 742
rect 3438 708 3442 712
rect 3454 698 3458 702
rect 3422 668 3426 672
rect 3414 658 3418 662
rect 3398 638 3402 642
rect 3398 618 3402 622
rect 3470 728 3474 732
rect 3486 718 3490 722
rect 3478 698 3482 702
rect 3502 698 3506 702
rect 3526 718 3530 722
rect 3566 858 3570 862
rect 3590 858 3594 862
rect 3646 858 3650 862
rect 3582 848 3586 852
rect 3606 848 3610 852
rect 3654 848 3658 852
rect 3670 848 3674 852
rect 3590 808 3594 812
rect 3570 803 3574 807
rect 3577 803 3581 807
rect 3566 768 3570 772
rect 3654 828 3658 832
rect 3686 848 3690 852
rect 3686 798 3690 802
rect 3678 758 3682 762
rect 3598 748 3602 752
rect 3622 748 3626 752
rect 3694 748 3698 752
rect 3598 738 3602 742
rect 3534 698 3538 702
rect 3622 728 3626 732
rect 3638 728 3642 732
rect 3590 718 3594 722
rect 3614 718 3618 722
rect 3582 688 3586 692
rect 3614 708 3618 712
rect 3606 698 3610 702
rect 3670 718 3674 722
rect 3662 678 3666 682
rect 3478 668 3482 672
rect 3598 668 3602 672
rect 3670 668 3674 672
rect 3510 658 3514 662
rect 3486 648 3490 652
rect 3478 638 3482 642
rect 3446 588 3450 592
rect 3454 578 3458 582
rect 3414 558 3418 562
rect 3470 558 3474 562
rect 3494 558 3498 562
rect 3406 548 3410 552
rect 3358 518 3362 522
rect 3342 508 3346 512
rect 3358 488 3362 492
rect 3342 458 3346 462
rect 3310 438 3314 442
rect 3318 438 3322 442
rect 3302 398 3306 402
rect 3270 368 3274 372
rect 3262 358 3266 362
rect 3294 358 3298 362
rect 3238 348 3242 352
rect 3246 338 3250 342
rect 3206 298 3210 302
rect 3254 308 3258 312
rect 3246 298 3250 302
rect 3238 278 3242 282
rect 3150 268 3154 272
rect 3190 268 3194 272
rect 3222 268 3226 272
rect 3110 168 3114 172
rect 3158 168 3162 172
rect 3094 158 3098 162
rect 3134 148 3138 152
rect 2950 138 2954 142
rect 2998 138 3002 142
rect 3038 138 3042 142
rect 2854 128 2858 132
rect 2942 128 2946 132
rect 2806 108 2810 112
rect 2830 108 2834 112
rect 2790 68 2794 72
rect 2750 58 2754 62
rect 2782 58 2786 62
rect 2702 48 2706 52
rect 2814 68 2818 72
rect 2918 108 2922 112
rect 2878 98 2882 102
rect 2910 98 2914 102
rect 2926 98 2930 102
rect 2838 68 2842 72
rect 2854 68 2858 72
rect 2878 68 2882 72
rect 2974 98 2978 102
rect 3038 108 3042 112
rect 3050 103 3054 107
rect 3057 103 3061 107
rect 3126 138 3130 142
rect 3278 338 3282 342
rect 3302 328 3306 332
rect 3294 298 3298 302
rect 3198 258 3202 262
rect 3222 258 3226 262
rect 3222 248 3226 252
rect 3254 248 3258 252
rect 3246 198 3250 202
rect 3230 168 3234 172
rect 3190 158 3194 162
rect 3166 148 3170 152
rect 3174 148 3178 152
rect 3182 138 3186 142
rect 3134 108 3138 112
rect 3158 98 3162 102
rect 3086 88 3090 92
rect 3070 78 3074 82
rect 3102 78 3106 82
rect 3142 78 3146 82
rect 2958 68 2962 72
rect 2934 58 2938 62
rect 3342 378 3346 382
rect 3374 498 3378 502
rect 3398 538 3402 542
rect 3390 528 3394 532
rect 3398 498 3402 502
rect 3414 528 3418 532
rect 3406 488 3410 492
rect 3406 448 3410 452
rect 3478 548 3482 552
rect 3454 538 3458 542
rect 3422 498 3426 502
rect 3430 498 3434 502
rect 3462 488 3466 492
rect 3438 478 3442 482
rect 3454 478 3458 482
rect 3422 468 3426 472
rect 3430 468 3434 472
rect 3542 658 3546 662
rect 3550 618 3554 622
rect 3570 603 3574 607
rect 3577 603 3581 607
rect 3534 558 3538 562
rect 3542 558 3546 562
rect 3590 558 3594 562
rect 3486 538 3490 542
rect 3694 718 3698 722
rect 3774 878 3778 882
rect 3822 878 3826 882
rect 3846 928 3850 932
rect 3878 918 3882 922
rect 3846 898 3850 902
rect 3726 868 3730 872
rect 3734 868 3738 872
rect 3758 868 3762 872
rect 3806 868 3810 872
rect 3830 868 3834 872
rect 3798 858 3802 862
rect 3782 848 3786 852
rect 3718 818 3722 822
rect 3766 838 3770 842
rect 3782 828 3786 832
rect 3726 768 3730 772
rect 3750 758 3754 762
rect 3782 758 3786 762
rect 3822 858 3826 862
rect 3838 848 3842 852
rect 3822 838 3826 842
rect 3806 828 3810 832
rect 3742 748 3746 752
rect 3798 748 3802 752
rect 3726 738 3730 742
rect 3750 738 3754 742
rect 3798 738 3802 742
rect 3774 728 3778 732
rect 3830 788 3834 792
rect 3854 878 3858 882
rect 3862 878 3866 882
rect 3870 838 3874 842
rect 3862 828 3866 832
rect 3870 828 3874 832
rect 3838 758 3842 762
rect 3854 758 3858 762
rect 3822 748 3826 752
rect 3838 738 3842 742
rect 3798 708 3802 712
rect 3806 708 3810 712
rect 3830 708 3834 712
rect 3750 688 3754 692
rect 3814 688 3818 692
rect 3710 678 3714 682
rect 3718 668 3722 672
rect 3806 678 3810 682
rect 3766 668 3770 672
rect 3686 658 3690 662
rect 3606 648 3610 652
rect 3630 648 3634 652
rect 3670 648 3674 652
rect 3614 638 3618 642
rect 3614 558 3618 562
rect 3606 548 3610 552
rect 3542 538 3546 542
rect 3598 538 3602 542
rect 3582 528 3586 532
rect 3502 488 3506 492
rect 3542 508 3546 512
rect 3430 458 3434 462
rect 3438 458 3442 462
rect 3462 458 3466 462
rect 3486 458 3490 462
rect 3374 378 3378 382
rect 3390 378 3394 382
rect 3358 328 3362 332
rect 3398 368 3402 372
rect 3382 358 3386 362
rect 3406 358 3410 362
rect 3390 328 3394 332
rect 3366 318 3370 322
rect 3406 318 3410 322
rect 3398 308 3402 312
rect 3390 278 3394 282
rect 3350 268 3354 272
rect 3374 268 3378 272
rect 3342 258 3346 262
rect 3390 258 3394 262
rect 3318 238 3322 242
rect 3334 238 3338 242
rect 3302 218 3306 222
rect 3342 228 3346 232
rect 3286 168 3290 172
rect 3318 168 3322 172
rect 3334 168 3338 172
rect 3238 158 3242 162
rect 3262 158 3266 162
rect 3278 158 3282 162
rect 3294 158 3298 162
rect 3334 158 3338 162
rect 3198 148 3202 152
rect 3230 138 3234 142
rect 3374 228 3378 232
rect 3358 168 3362 172
rect 3350 148 3354 152
rect 3270 118 3274 122
rect 3222 108 3226 112
rect 3270 108 3274 112
rect 3294 118 3298 122
rect 3230 98 3234 102
rect 3270 98 3274 102
rect 3278 98 3282 102
rect 3166 78 3170 82
rect 3198 78 3202 82
rect 3206 78 3210 82
rect 3310 108 3314 112
rect 3278 88 3282 92
rect 3302 88 3306 92
rect 3262 78 3266 82
rect 2982 58 2986 62
rect 3030 58 3034 62
rect 3038 58 3042 62
rect 3070 58 3074 62
rect 3366 158 3370 162
rect 3454 448 3458 452
rect 3462 358 3466 362
rect 3446 348 3450 352
rect 3438 328 3442 332
rect 3454 318 3458 322
rect 3414 288 3418 292
rect 3438 288 3442 292
rect 3486 348 3490 352
rect 3558 458 3562 462
rect 3598 458 3602 462
rect 3630 498 3634 502
rect 3622 488 3626 492
rect 3622 468 3626 472
rect 3686 608 3690 612
rect 3678 598 3682 602
rect 3670 568 3674 572
rect 3718 648 3722 652
rect 3702 578 3706 582
rect 3702 568 3706 572
rect 3726 638 3730 642
rect 3734 638 3738 642
rect 3710 548 3714 552
rect 3662 528 3666 532
rect 3646 458 3650 462
rect 3678 458 3682 462
rect 3526 438 3530 442
rect 3518 368 3522 372
rect 3570 403 3574 407
rect 3577 403 3581 407
rect 3606 418 3610 422
rect 3598 398 3602 402
rect 3670 448 3674 452
rect 3686 448 3690 452
rect 3670 428 3674 432
rect 3766 608 3770 612
rect 3742 568 3746 572
rect 3718 528 3722 532
rect 3726 528 3730 532
rect 3742 488 3746 492
rect 3798 668 3802 672
rect 3798 658 3802 662
rect 3854 728 3858 732
rect 3846 718 3850 722
rect 3910 938 3914 942
rect 3894 928 3898 932
rect 3998 1028 4002 1032
rect 4006 1008 4010 1012
rect 3982 998 3986 1002
rect 4126 1228 4130 1232
rect 4110 1188 4114 1192
rect 4102 1168 4106 1172
rect 4118 1138 4122 1142
rect 4142 1248 4146 1252
rect 4142 1208 4146 1212
rect 4166 1258 4170 1262
rect 4182 1258 4186 1262
rect 4222 1428 4226 1432
rect 4310 1458 4314 1462
rect 4294 1448 4298 1452
rect 4230 1418 4234 1422
rect 4286 1418 4290 1422
rect 4238 1388 4242 1392
rect 4286 1388 4290 1392
rect 4246 1368 4250 1372
rect 4230 1358 4234 1362
rect 4270 1358 4274 1362
rect 4366 1538 4370 1542
rect 4350 1528 4354 1532
rect 4342 1478 4346 1482
rect 4334 1468 4338 1472
rect 4278 1348 4282 1352
rect 4206 1328 4210 1332
rect 4230 1338 4234 1342
rect 4230 1318 4234 1322
rect 4278 1338 4282 1342
rect 4278 1328 4282 1332
rect 4278 1318 4282 1322
rect 4238 1288 4242 1292
rect 4254 1288 4258 1292
rect 4166 1238 4170 1242
rect 4150 1198 4154 1202
rect 4150 1178 4154 1182
rect 4142 1158 4146 1162
rect 4190 1228 4194 1232
rect 4174 1218 4178 1222
rect 4198 1218 4202 1222
rect 4182 1178 4186 1182
rect 4262 1258 4266 1262
rect 4278 1248 4282 1252
rect 4294 1248 4298 1252
rect 4214 1228 4218 1232
rect 4286 1228 4290 1232
rect 4318 1338 4322 1342
rect 4342 1458 4346 1462
rect 4334 1438 4338 1442
rect 4358 1438 4362 1442
rect 4334 1368 4338 1372
rect 4390 1528 4394 1532
rect 4398 1498 4402 1502
rect 4590 1678 4594 1682
rect 4582 1668 4586 1672
rect 4470 1538 4474 1542
rect 4486 1538 4490 1542
rect 4454 1528 4458 1532
rect 4382 1478 4386 1482
rect 4374 1468 4378 1472
rect 4398 1468 4402 1472
rect 4438 1468 4442 1472
rect 4374 1458 4378 1462
rect 4414 1458 4418 1462
rect 4382 1448 4386 1452
rect 4422 1448 4426 1452
rect 4430 1448 4434 1452
rect 4494 1478 4498 1482
rect 4462 1468 4466 1472
rect 4486 1468 4490 1472
rect 4470 1458 4474 1462
rect 4502 1458 4506 1462
rect 4454 1438 4458 1442
rect 4534 1538 4538 1542
rect 4558 1528 4562 1532
rect 4566 1528 4570 1532
rect 4550 1488 4554 1492
rect 4542 1468 4546 1472
rect 4550 1468 4554 1472
rect 4582 1468 4586 1472
rect 4478 1448 4482 1452
rect 4510 1448 4514 1452
rect 4462 1408 4466 1412
rect 4510 1438 4514 1442
rect 4390 1378 4394 1382
rect 4446 1378 4450 1382
rect 4374 1368 4378 1372
rect 4326 1328 4330 1332
rect 4326 1308 4330 1312
rect 4318 1298 4322 1302
rect 4350 1358 4354 1362
rect 4342 1338 4346 1342
rect 4334 1298 4338 1302
rect 4494 1368 4498 1372
rect 4406 1358 4410 1362
rect 4486 1358 4490 1362
rect 4470 1348 4474 1352
rect 4430 1338 4434 1342
rect 4454 1338 4458 1342
rect 4542 1458 4546 1462
rect 4582 1458 4586 1462
rect 4550 1448 4554 1452
rect 4566 1438 4570 1442
rect 4550 1428 4554 1432
rect 4518 1388 4522 1392
rect 4518 1358 4522 1362
rect 4494 1348 4498 1352
rect 4510 1338 4514 1342
rect 4398 1328 4402 1332
rect 4366 1308 4370 1312
rect 4350 1278 4354 1282
rect 4334 1228 4338 1232
rect 4302 1218 4306 1222
rect 4214 1208 4218 1212
rect 4206 1178 4210 1182
rect 4222 1178 4226 1182
rect 4166 1148 4170 1152
rect 4190 1148 4194 1152
rect 4150 1138 4154 1142
rect 4110 1128 4114 1132
rect 4118 1128 4122 1132
rect 4134 1128 4138 1132
rect 4150 1128 4154 1132
rect 4174 1128 4178 1132
rect 4082 1103 4086 1107
rect 4089 1103 4093 1107
rect 4078 1078 4082 1082
rect 4110 1078 4114 1082
rect 4094 1068 4098 1072
rect 4126 1098 4130 1102
rect 4294 1198 4298 1202
rect 4254 1168 4258 1172
rect 4222 1138 4226 1142
rect 4230 1128 4234 1132
rect 4134 1078 4138 1082
rect 4166 1078 4170 1082
rect 4190 1078 4194 1082
rect 4198 1078 4202 1082
rect 4158 1068 4162 1072
rect 4182 1068 4186 1072
rect 4102 1038 4106 1042
rect 4070 998 4074 1002
rect 4070 958 4074 962
rect 3974 948 3978 952
rect 3942 878 3946 882
rect 3950 878 3954 882
rect 3998 948 4002 952
rect 4094 948 4098 952
rect 4014 938 4018 942
rect 4054 938 4058 942
rect 4022 928 4026 932
rect 4030 928 4034 932
rect 3998 888 4002 892
rect 3982 878 3986 882
rect 3894 858 3898 862
rect 3942 858 3946 862
rect 3966 858 3970 862
rect 3990 858 3994 862
rect 3918 848 3922 852
rect 3958 848 3962 852
rect 3982 848 3986 852
rect 3886 838 3890 842
rect 3942 838 3946 842
rect 3966 838 3970 842
rect 3910 788 3914 792
rect 3886 758 3890 762
rect 3990 828 3994 832
rect 3974 788 3978 792
rect 4046 918 4050 922
rect 4038 908 4042 912
rect 4046 898 4050 902
rect 4022 878 4026 882
rect 4038 838 4042 842
rect 4014 828 4018 832
rect 4062 858 4066 862
rect 4094 938 4098 942
rect 4082 903 4086 907
rect 4089 903 4093 907
rect 4198 1058 4202 1062
rect 4198 1028 4202 1032
rect 4270 1158 4274 1162
rect 4406 1288 4410 1292
rect 4374 1278 4378 1282
rect 4438 1268 4442 1272
rect 4366 1258 4370 1262
rect 4374 1258 4378 1262
rect 4390 1258 4394 1262
rect 4310 1178 4314 1182
rect 4350 1178 4354 1182
rect 4382 1248 4386 1252
rect 4422 1248 4426 1252
rect 4406 1238 4410 1242
rect 4478 1298 4482 1302
rect 4462 1268 4466 1272
rect 4494 1278 4498 1282
rect 4486 1268 4490 1272
rect 4574 1388 4578 1392
rect 4574 1358 4578 1362
rect 4558 1348 4562 1352
rect 4582 1328 4586 1332
rect 4598 1338 4602 1342
rect 4590 1288 4594 1292
rect 4518 1278 4522 1282
rect 4534 1278 4538 1282
rect 4550 1268 4554 1272
rect 4462 1248 4466 1252
rect 4494 1248 4498 1252
rect 4390 1218 4394 1222
rect 4398 1218 4402 1222
rect 4398 1198 4402 1202
rect 4374 1188 4378 1192
rect 4390 1188 4394 1192
rect 4286 1148 4290 1152
rect 4310 1148 4314 1152
rect 4262 1138 4266 1142
rect 4278 1138 4282 1142
rect 4254 1098 4258 1102
rect 4270 1088 4274 1092
rect 4310 1138 4314 1142
rect 4334 1138 4338 1142
rect 4326 1128 4330 1132
rect 4302 1098 4306 1102
rect 4334 1098 4338 1102
rect 4254 1068 4258 1072
rect 4278 1078 4282 1082
rect 4182 1018 4186 1022
rect 4134 1008 4138 1012
rect 4134 958 4138 962
rect 4118 948 4122 952
rect 4134 948 4138 952
rect 4150 948 4154 952
rect 4118 928 4122 932
rect 4126 878 4130 882
rect 4110 868 4114 872
rect 4094 858 4098 862
rect 4062 848 4066 852
rect 4046 808 4050 812
rect 4206 1008 4210 1012
rect 4166 948 4170 952
rect 4190 948 4194 952
rect 4206 918 4210 922
rect 4326 1088 4330 1092
rect 4350 1088 4354 1092
rect 4294 1068 4298 1072
rect 4334 1078 4338 1082
rect 4334 1058 4338 1062
rect 4310 1048 4314 1052
rect 4262 1028 4266 1032
rect 4286 1028 4290 1032
rect 4302 1028 4306 1032
rect 4246 998 4250 1002
rect 4254 998 4258 1002
rect 4230 978 4234 982
rect 4286 968 4290 972
rect 4318 958 4322 962
rect 4238 948 4242 952
rect 4254 948 4258 952
rect 4246 938 4250 942
rect 4230 918 4234 922
rect 4174 878 4178 882
rect 4190 878 4194 882
rect 4198 878 4202 882
rect 4214 878 4218 882
rect 4174 868 4178 872
rect 4158 848 4162 852
rect 4134 798 4138 802
rect 4046 788 4050 792
rect 4006 768 4010 772
rect 4014 758 4018 762
rect 4222 868 4226 872
rect 4238 898 4242 902
rect 4246 888 4250 892
rect 4238 868 4242 872
rect 4230 858 4234 862
rect 4190 848 4194 852
rect 4222 848 4226 852
rect 4198 838 4202 842
rect 4214 838 4218 842
rect 4246 838 4250 842
rect 4238 828 4242 832
rect 4334 1048 4338 1052
rect 4294 948 4298 952
rect 4326 948 4330 952
rect 4286 938 4290 942
rect 4310 938 4314 942
rect 4302 928 4306 932
rect 4350 1018 4354 1022
rect 4382 1108 4386 1112
rect 4366 1068 4370 1072
rect 4398 1148 4402 1152
rect 4446 1178 4450 1182
rect 4518 1248 4522 1252
rect 4502 1218 4506 1222
rect 4510 1208 4514 1212
rect 4558 1258 4562 1262
rect 4542 1238 4546 1242
rect 4582 1188 4586 1192
rect 4566 1168 4570 1172
rect 4462 1158 4466 1162
rect 4518 1158 4522 1162
rect 4534 1158 4538 1162
rect 4558 1158 4562 1162
rect 4422 1148 4426 1152
rect 4430 1148 4434 1152
rect 4398 1108 4402 1112
rect 4430 1098 4434 1102
rect 4414 1078 4418 1082
rect 4398 1068 4402 1072
rect 4422 1068 4426 1072
rect 4438 1058 4442 1062
rect 4478 1138 4482 1142
rect 4486 1138 4490 1142
rect 4454 1088 4458 1092
rect 4502 1108 4506 1112
rect 4494 1098 4498 1102
rect 4486 1088 4490 1092
rect 4454 1078 4458 1082
rect 4462 1068 4466 1072
rect 4478 1068 4482 1072
rect 4486 1058 4490 1062
rect 4390 1048 4394 1052
rect 4406 1048 4410 1052
rect 4438 1048 4442 1052
rect 4446 1048 4450 1052
rect 4382 1028 4386 1032
rect 4438 1018 4442 1022
rect 4374 1008 4378 1012
rect 4382 1008 4386 1012
rect 4382 988 4386 992
rect 4358 958 4362 962
rect 4398 958 4402 962
rect 4430 958 4434 962
rect 4350 948 4354 952
rect 4334 908 4338 912
rect 4262 898 4266 902
rect 4270 898 4274 902
rect 4326 878 4330 882
rect 4278 868 4282 872
rect 4294 868 4298 872
rect 4270 858 4274 862
rect 4278 858 4282 862
rect 4206 818 4210 822
rect 4254 818 4258 822
rect 4166 778 4170 782
rect 4198 778 4202 782
rect 4110 758 4114 762
rect 4166 758 4170 762
rect 3958 748 3962 752
rect 4006 748 4010 752
rect 4022 748 4026 752
rect 3910 738 3914 742
rect 3926 738 3930 742
rect 4030 738 4034 742
rect 4062 738 4066 742
rect 4110 738 4114 742
rect 4142 738 4146 742
rect 4046 728 4050 732
rect 3902 678 3906 682
rect 3886 668 3890 672
rect 3950 668 3954 672
rect 3958 668 3962 672
rect 3814 648 3818 652
rect 3838 648 3842 652
rect 3862 638 3866 642
rect 3822 618 3826 622
rect 3854 618 3858 622
rect 3790 598 3794 602
rect 3902 648 3906 652
rect 3918 638 3922 642
rect 3934 608 3938 612
rect 3870 598 3874 602
rect 3854 578 3858 582
rect 3878 578 3882 582
rect 3926 578 3930 582
rect 3838 568 3842 572
rect 3766 558 3770 562
rect 3790 558 3794 562
rect 3830 558 3834 562
rect 3814 548 3818 552
rect 3782 538 3786 542
rect 3798 528 3802 532
rect 3838 548 3842 552
rect 3822 538 3826 542
rect 3854 568 3858 572
rect 3870 558 3874 562
rect 3902 558 3906 562
rect 3854 548 3858 552
rect 3846 538 3850 542
rect 3758 508 3762 512
rect 3806 508 3810 512
rect 3758 478 3762 482
rect 3806 478 3810 482
rect 3814 468 3818 472
rect 3710 458 3714 462
rect 3742 458 3746 462
rect 3878 528 3882 532
rect 3886 528 3890 532
rect 3894 498 3898 502
rect 3854 488 3858 492
rect 3878 488 3882 492
rect 3886 488 3890 492
rect 3830 478 3834 482
rect 3862 478 3866 482
rect 3846 468 3850 472
rect 3854 468 3858 472
rect 3878 468 3882 472
rect 3782 448 3786 452
rect 3798 438 3802 442
rect 3718 428 3722 432
rect 3702 418 3706 422
rect 3766 418 3770 422
rect 3678 398 3682 402
rect 3606 368 3610 372
rect 3534 358 3538 362
rect 3558 358 3562 362
rect 3518 348 3522 352
rect 3502 328 3506 332
rect 3446 278 3450 282
rect 3470 278 3474 282
rect 3494 278 3498 282
rect 3406 268 3410 272
rect 3422 268 3426 272
rect 3550 328 3554 332
rect 3510 288 3514 292
rect 3526 288 3530 292
rect 3454 268 3458 272
rect 3502 268 3506 272
rect 3566 308 3570 312
rect 3566 298 3570 302
rect 3574 298 3578 302
rect 3542 278 3546 282
rect 3550 278 3554 282
rect 3414 238 3418 242
rect 3470 238 3474 242
rect 3486 218 3490 222
rect 3510 218 3514 222
rect 3518 208 3522 212
rect 3438 198 3442 202
rect 3486 198 3490 202
rect 3494 198 3498 202
rect 3454 158 3458 162
rect 3374 118 3378 122
rect 3382 108 3386 112
rect 3326 78 3330 82
rect 3342 78 3346 82
rect 3366 68 3370 72
rect 3398 88 3402 92
rect 3390 78 3394 82
rect 3342 58 3346 62
rect 3382 58 3386 62
rect 3422 138 3426 142
rect 3478 148 3482 152
rect 3462 138 3466 142
rect 3470 118 3474 122
rect 3438 108 3442 112
rect 3430 98 3434 102
rect 3446 98 3450 102
rect 3558 238 3562 242
rect 3598 278 3602 282
rect 3638 358 3642 362
rect 3630 348 3634 352
rect 3654 348 3658 352
rect 3622 328 3626 332
rect 3614 288 3618 292
rect 3590 258 3594 262
rect 3662 328 3666 332
rect 3646 278 3650 282
rect 3654 278 3658 282
rect 3662 278 3666 282
rect 3590 238 3594 242
rect 3614 238 3618 242
rect 3574 228 3578 232
rect 3570 203 3574 207
rect 3577 203 3581 207
rect 3550 178 3554 182
rect 3510 148 3514 152
rect 3526 148 3530 152
rect 3534 148 3538 152
rect 3542 138 3546 142
rect 3534 128 3538 132
rect 3518 108 3522 112
rect 3526 108 3530 112
rect 3574 138 3578 142
rect 3550 128 3554 132
rect 3558 128 3562 132
rect 3606 118 3610 122
rect 3590 98 3594 102
rect 3662 218 3666 222
rect 3622 198 3626 202
rect 3630 178 3634 182
rect 3654 178 3658 182
rect 3598 88 3602 92
rect 3422 78 3426 82
rect 3438 78 3442 82
rect 3646 158 3650 162
rect 3686 368 3690 372
rect 4126 728 4130 732
rect 4182 748 4186 752
rect 4190 738 4194 742
rect 4126 718 4130 722
rect 4158 718 4162 722
rect 4102 708 4106 712
rect 4082 703 4086 707
rect 4089 703 4093 707
rect 4110 698 4114 702
rect 3990 688 3994 692
rect 4030 678 4034 682
rect 4046 678 4050 682
rect 4070 678 4074 682
rect 4038 668 4042 672
rect 3982 658 3986 662
rect 3998 658 4002 662
rect 4102 668 4106 672
rect 4054 658 4058 662
rect 3998 648 4002 652
rect 4014 648 4018 652
rect 4038 648 4042 652
rect 3998 618 4002 622
rect 4022 618 4026 622
rect 3974 608 3978 612
rect 4014 608 4018 612
rect 3958 558 3962 562
rect 3966 558 3970 562
rect 3934 538 3938 542
rect 3950 538 3954 542
rect 3918 528 3922 532
rect 3926 528 3930 532
rect 3910 498 3914 502
rect 3910 478 3914 482
rect 3934 518 3938 522
rect 3942 508 3946 512
rect 3950 508 3954 512
rect 3918 458 3922 462
rect 3942 458 3946 462
rect 3958 458 3962 462
rect 3950 448 3954 452
rect 3958 448 3962 452
rect 3822 438 3826 442
rect 3830 438 3834 442
rect 3846 438 3850 442
rect 3934 438 3938 442
rect 3734 408 3738 412
rect 3814 408 3818 412
rect 3934 408 3938 412
rect 3942 408 3946 412
rect 3806 368 3810 372
rect 3926 368 3930 372
rect 3718 358 3722 362
rect 3766 358 3770 362
rect 3694 348 3698 352
rect 3726 348 3730 352
rect 3734 348 3738 352
rect 3678 328 3682 332
rect 3694 298 3698 302
rect 3742 338 3746 342
rect 3710 328 3714 332
rect 3710 308 3714 312
rect 3774 348 3778 352
rect 3750 298 3754 302
rect 3702 278 3706 282
rect 3718 278 3722 282
rect 3686 268 3690 272
rect 3742 268 3746 272
rect 3678 258 3682 262
rect 3710 258 3714 262
rect 3718 258 3722 262
rect 3678 208 3682 212
rect 3670 188 3674 192
rect 3742 228 3746 232
rect 3734 188 3738 192
rect 3686 158 3690 162
rect 3694 158 3698 162
rect 3710 158 3714 162
rect 3702 148 3706 152
rect 3718 138 3722 142
rect 3734 138 3738 142
rect 3710 128 3714 132
rect 3694 118 3698 122
rect 3670 98 3674 102
rect 3622 78 3626 82
rect 3438 68 3442 72
rect 3462 68 3466 72
rect 3478 68 3482 72
rect 3502 68 3506 72
rect 3550 68 3554 72
rect 3598 68 3602 72
rect 3630 68 3634 72
rect 3638 68 3642 72
rect 3670 68 3674 72
rect 3430 58 3434 62
rect 3454 58 3458 62
rect 3478 58 3482 62
rect 3494 58 3498 62
rect 3526 58 3530 62
rect 3574 58 3578 62
rect 2910 48 2914 52
rect 2958 48 2962 52
rect 2974 48 2978 52
rect 3006 48 3010 52
rect 3014 48 3018 52
rect 3054 48 3058 52
rect 3126 48 3130 52
rect 3174 48 3178 52
rect 3214 48 3218 52
rect 3238 48 3242 52
rect 3254 48 3258 52
rect 3278 48 3282 52
rect 3286 48 3290 52
rect 3310 48 3314 52
rect 3406 48 3410 52
rect 3606 48 3610 52
rect 3414 38 3418 42
rect 3654 38 3658 42
rect 3118 28 3122 32
rect 3342 28 3346 32
rect 3078 18 3082 22
rect 1522 3 1526 7
rect 1529 3 1533 7
rect 3702 78 3706 82
rect 3718 68 3722 72
rect 3702 58 3706 62
rect 3694 48 3698 52
rect 3838 338 3842 342
rect 3790 328 3794 332
rect 3814 328 3818 332
rect 3838 328 3842 332
rect 3822 318 3826 322
rect 3814 308 3818 312
rect 3830 288 3834 292
rect 3958 408 3962 412
rect 3950 398 3954 402
rect 3894 348 3898 352
rect 3854 328 3858 332
rect 3854 318 3858 322
rect 3862 288 3866 292
rect 3830 268 3834 272
rect 3846 268 3850 272
rect 3862 268 3866 272
rect 3782 238 3786 242
rect 3774 208 3778 212
rect 3758 188 3762 192
rect 3822 258 3826 262
rect 3854 248 3858 252
rect 3878 298 3882 302
rect 4062 588 4066 592
rect 3982 548 3986 552
rect 4030 548 4034 552
rect 4046 548 4050 552
rect 4062 548 4066 552
rect 4086 548 4090 552
rect 3974 528 3978 532
rect 3990 528 3994 532
rect 3990 518 3994 522
rect 3998 518 4002 522
rect 3974 498 3978 502
rect 3982 488 3986 492
rect 4102 648 4106 652
rect 4166 698 4170 702
rect 4158 678 4162 682
rect 4190 708 4194 712
rect 4238 808 4242 812
rect 4214 778 4218 782
rect 4262 778 4266 782
rect 4238 768 4242 772
rect 4238 758 4242 762
rect 4214 748 4218 752
rect 4246 738 4250 742
rect 4238 728 4242 732
rect 4238 688 4242 692
rect 4254 688 4258 692
rect 4206 678 4210 682
rect 4262 678 4266 682
rect 4174 668 4178 672
rect 4182 668 4186 672
rect 4118 638 4122 642
rect 4190 658 4194 662
rect 4142 608 4146 612
rect 4230 668 4234 672
rect 4254 668 4258 672
rect 4206 638 4210 642
rect 4166 608 4170 612
rect 4182 608 4186 612
rect 4150 578 4154 582
rect 4118 548 4122 552
rect 4126 548 4130 552
rect 4038 538 4042 542
rect 4054 538 4058 542
rect 4094 538 4098 542
rect 4126 538 4130 542
rect 4022 528 4026 532
rect 4006 498 4010 502
rect 3998 488 4002 492
rect 4062 498 4066 502
rect 4054 488 4058 492
rect 4062 478 4066 482
rect 4158 548 4162 552
rect 4190 588 4194 592
rect 4134 528 4138 532
rect 4142 528 4146 532
rect 4158 528 4162 532
rect 4082 503 4086 507
rect 4089 503 4093 507
rect 4102 488 4106 492
rect 3998 468 4002 472
rect 4006 468 4010 472
rect 4022 468 4026 472
rect 4038 468 4042 472
rect 4054 468 4058 472
rect 4022 438 4026 442
rect 3974 398 3978 402
rect 4006 398 4010 402
rect 4038 398 4042 402
rect 4046 398 4050 402
rect 4070 378 4074 382
rect 4022 368 4026 372
rect 4062 368 4066 372
rect 3966 358 3970 362
rect 4014 358 4018 362
rect 3974 348 3978 352
rect 3982 348 3986 352
rect 3990 348 3994 352
rect 3950 338 3954 342
rect 3918 328 3922 332
rect 3942 328 3946 332
rect 3910 318 3914 322
rect 3910 308 3914 312
rect 3894 288 3898 292
rect 3982 328 3986 332
rect 4006 328 4010 332
rect 3990 318 3994 322
rect 3998 308 4002 312
rect 3950 288 3954 292
rect 3966 288 3970 292
rect 3942 278 3946 282
rect 3958 278 3962 282
rect 3966 278 3970 282
rect 3926 258 3930 262
rect 3942 258 3946 262
rect 3950 258 3954 262
rect 3838 238 3842 242
rect 3870 238 3874 242
rect 3974 238 3978 242
rect 3798 198 3802 202
rect 3782 188 3786 192
rect 3774 148 3778 152
rect 3758 138 3762 142
rect 3814 168 3818 172
rect 3798 158 3802 162
rect 3862 218 3866 222
rect 3902 218 3906 222
rect 3958 218 3962 222
rect 3854 198 3858 202
rect 3846 158 3850 162
rect 3790 148 3794 152
rect 3822 148 3826 152
rect 3830 138 3834 142
rect 3838 138 3842 142
rect 3774 128 3778 132
rect 3750 108 3754 112
rect 3750 78 3754 82
rect 3766 78 3770 82
rect 3854 148 3858 152
rect 3870 148 3874 152
rect 3894 148 3898 152
rect 3886 138 3890 142
rect 3910 208 3914 212
rect 3934 178 3938 182
rect 4022 348 4026 352
rect 4046 348 4050 352
rect 4046 338 4050 342
rect 4062 338 4066 342
rect 4150 498 4154 502
rect 4158 498 4162 502
rect 4174 498 4178 502
rect 4126 478 4130 482
rect 4110 468 4114 472
rect 4118 468 4122 472
rect 4142 468 4146 472
rect 4174 488 4178 492
rect 4198 568 4202 572
rect 4374 898 4378 902
rect 4318 868 4322 872
rect 4366 868 4370 872
rect 4414 948 4418 952
rect 4454 1008 4458 1012
rect 4470 978 4474 982
rect 4446 968 4450 972
rect 4454 968 4458 972
rect 4470 958 4474 962
rect 4406 928 4410 932
rect 4390 908 4394 912
rect 4414 898 4418 902
rect 4510 1048 4514 1052
rect 4494 988 4498 992
rect 4510 958 4514 962
rect 4454 938 4458 942
rect 4478 938 4482 942
rect 4478 908 4482 912
rect 4502 928 4506 932
rect 4558 1128 4562 1132
rect 4534 1068 4538 1072
rect 4534 1058 4538 1062
rect 4526 1038 4530 1042
rect 4542 1038 4546 1042
rect 4526 968 4530 972
rect 4526 918 4530 922
rect 4486 898 4490 902
rect 4518 898 4522 902
rect 4478 878 4482 882
rect 4430 868 4434 872
rect 4414 858 4418 862
rect 4302 848 4306 852
rect 4294 838 4298 842
rect 4286 788 4290 792
rect 4326 828 4330 832
rect 4318 788 4322 792
rect 4382 848 4386 852
rect 4422 838 4426 842
rect 4470 858 4474 862
rect 4502 858 4506 862
rect 4518 858 4522 862
rect 4454 848 4458 852
rect 4510 848 4514 852
rect 4430 818 4434 822
rect 4438 818 4442 822
rect 4374 808 4378 812
rect 4382 778 4386 782
rect 4414 768 4418 772
rect 4422 768 4426 772
rect 4286 738 4290 742
rect 4294 728 4298 732
rect 4294 718 4298 722
rect 4318 738 4322 742
rect 4310 698 4314 702
rect 4358 738 4362 742
rect 4382 738 4386 742
rect 4390 738 4394 742
rect 4406 738 4410 742
rect 4342 728 4346 732
rect 4350 728 4354 732
rect 4398 728 4402 732
rect 4382 718 4386 722
rect 4374 698 4378 702
rect 4366 688 4370 692
rect 4286 678 4290 682
rect 4294 678 4298 682
rect 4278 658 4282 662
rect 4214 598 4218 602
rect 4246 648 4250 652
rect 4230 618 4234 622
rect 4270 638 4274 642
rect 4342 668 4346 672
rect 4366 668 4370 672
rect 4374 668 4378 672
rect 4310 658 4314 662
rect 4318 648 4322 652
rect 4310 638 4314 642
rect 4222 578 4226 582
rect 4238 578 4242 582
rect 4198 528 4202 532
rect 4198 478 4202 482
rect 4206 448 4210 452
rect 4118 358 4122 362
rect 4102 338 4106 342
rect 4022 308 4026 312
rect 4030 298 4034 302
rect 4038 288 4042 292
rect 3998 258 4002 262
rect 4014 258 4018 262
rect 4038 258 4042 262
rect 3990 168 3994 172
rect 4006 168 4010 172
rect 3934 158 3938 162
rect 3950 158 3954 162
rect 3910 138 3914 142
rect 3782 108 3786 112
rect 3798 108 3802 112
rect 3886 108 3890 112
rect 3902 108 3906 112
rect 3878 88 3882 92
rect 3790 78 3794 82
rect 3862 78 3866 82
rect 3838 68 3842 72
rect 4022 218 4026 222
rect 4070 328 4074 332
rect 4094 328 4098 332
rect 4082 303 4086 307
rect 4089 303 4093 307
rect 4070 298 4074 302
rect 4054 278 4058 282
rect 4110 318 4114 322
rect 4190 438 4194 442
rect 4174 408 4178 412
rect 4150 368 4154 372
rect 4166 368 4170 372
rect 4214 408 4218 412
rect 4206 398 4210 402
rect 4278 568 4282 572
rect 4302 568 4306 572
rect 4254 548 4258 552
rect 4246 528 4250 532
rect 4286 548 4290 552
rect 4294 528 4298 532
rect 4246 518 4250 522
rect 4262 518 4266 522
rect 4238 488 4242 492
rect 4254 478 4258 482
rect 4294 508 4298 512
rect 4350 638 4354 642
rect 4334 628 4338 632
rect 4350 628 4354 632
rect 4318 588 4322 592
rect 4414 698 4418 702
rect 4518 838 4522 842
rect 4534 828 4538 832
rect 4550 1028 4554 1032
rect 4598 1168 4602 1172
rect 4590 1118 4594 1122
rect 4598 1028 4602 1032
rect 4550 958 4554 962
rect 4558 948 4562 952
rect 4550 938 4554 942
rect 4574 918 4578 922
rect 4550 878 4554 882
rect 4566 878 4570 882
rect 4582 878 4586 882
rect 4470 768 4474 772
rect 4518 768 4522 772
rect 4542 768 4546 772
rect 4454 758 4458 762
rect 4438 738 4442 742
rect 4430 728 4434 732
rect 4406 658 4410 662
rect 4422 658 4426 662
rect 4398 618 4402 622
rect 4382 608 4386 612
rect 4326 578 4330 582
rect 4390 578 4394 582
rect 4446 678 4450 682
rect 4470 738 4474 742
rect 4462 708 4466 712
rect 4438 648 4442 652
rect 4454 648 4458 652
rect 4430 638 4434 642
rect 4414 628 4418 632
rect 4406 568 4410 572
rect 4382 548 4386 552
rect 4318 528 4322 532
rect 4374 528 4378 532
rect 4366 508 4370 512
rect 4478 718 4482 722
rect 4494 728 4498 732
rect 4510 718 4514 722
rect 4486 708 4490 712
rect 4494 668 4498 672
rect 4486 658 4490 662
rect 4478 648 4482 652
rect 4470 618 4474 622
rect 4454 588 4458 592
rect 4462 568 4466 572
rect 4406 548 4410 552
rect 4438 548 4442 552
rect 4446 518 4450 522
rect 4430 508 4434 512
rect 4502 658 4506 662
rect 4494 638 4498 642
rect 4486 588 4490 592
rect 4502 578 4506 582
rect 4534 748 4538 752
rect 4526 728 4530 732
rect 4542 728 4546 732
rect 4534 718 4538 722
rect 4542 708 4546 712
rect 4590 838 4594 842
rect 4574 818 4578 822
rect 4574 718 4578 722
rect 4598 708 4602 712
rect 4550 698 4554 702
rect 4566 678 4570 682
rect 4526 668 4530 672
rect 4526 658 4530 662
rect 4574 618 4578 622
rect 4574 608 4578 612
rect 4558 598 4562 602
rect 4550 568 4554 572
rect 4558 568 4562 572
rect 4526 558 4530 562
rect 4518 548 4522 552
rect 4550 548 4554 552
rect 4582 548 4586 552
rect 4478 538 4482 542
rect 4462 528 4466 532
rect 4470 508 4474 512
rect 4398 498 4402 502
rect 4414 498 4418 502
rect 4366 488 4370 492
rect 4382 488 4386 492
rect 4414 488 4418 492
rect 4462 488 4466 492
rect 4310 478 4314 482
rect 4326 478 4330 482
rect 4350 478 4354 482
rect 4302 458 4306 462
rect 4238 448 4242 452
rect 4278 448 4282 452
rect 4230 378 4234 382
rect 4238 358 4242 362
rect 4262 408 4266 412
rect 4334 468 4338 472
rect 4318 458 4322 462
rect 4318 438 4322 442
rect 4334 428 4338 432
rect 4310 418 4314 422
rect 4398 468 4402 472
rect 4510 528 4514 532
rect 4502 488 4506 492
rect 4518 478 4522 482
rect 4350 458 4354 462
rect 4398 458 4402 462
rect 4470 458 4474 462
rect 4494 458 4498 462
rect 4518 458 4522 462
rect 4366 438 4370 442
rect 4390 408 4394 412
rect 4278 388 4282 392
rect 4302 358 4306 362
rect 4318 358 4322 362
rect 4222 348 4226 352
rect 4246 348 4250 352
rect 4254 348 4258 352
rect 4270 348 4274 352
rect 4278 348 4282 352
rect 4310 348 4314 352
rect 4350 348 4354 352
rect 4382 348 4386 352
rect 4142 338 4146 342
rect 4126 298 4130 302
rect 4102 288 4106 292
rect 4110 288 4114 292
rect 4110 268 4114 272
rect 4078 248 4082 252
rect 4062 238 4066 242
rect 4054 208 4058 212
rect 4062 208 4066 212
rect 4054 188 4058 192
rect 4046 178 4050 182
rect 4030 148 4034 152
rect 3942 138 3946 142
rect 3966 138 3970 142
rect 3982 138 3986 142
rect 3990 138 3994 142
rect 4022 138 4026 142
rect 4102 258 4106 262
rect 4134 258 4138 262
rect 4086 198 4090 202
rect 4166 248 4170 252
rect 4158 238 4162 242
rect 4126 228 4130 232
rect 4150 228 4154 232
rect 4166 228 4170 232
rect 4118 188 4122 192
rect 4094 158 4098 162
rect 4110 158 4114 162
rect 4142 188 4146 192
rect 4142 168 4146 172
rect 4134 148 4138 152
rect 4150 148 4154 152
rect 4190 338 4194 342
rect 4182 328 4186 332
rect 4214 328 4218 332
rect 4230 328 4234 332
rect 4246 328 4250 332
rect 4286 328 4290 332
rect 4310 328 4314 332
rect 4190 318 4194 322
rect 4198 318 4202 322
rect 4198 308 4202 312
rect 4246 308 4250 312
rect 4182 278 4186 282
rect 4206 278 4210 282
rect 4222 278 4226 282
rect 4222 258 4226 262
rect 4182 228 4186 232
rect 4238 238 4242 242
rect 4214 208 4218 212
rect 4174 158 4178 162
rect 4190 158 4194 162
rect 4198 158 4202 162
rect 4206 148 4210 152
rect 4118 138 4122 142
rect 4158 138 4162 142
rect 3926 128 3930 132
rect 3950 128 3954 132
rect 3982 128 3986 132
rect 4014 128 4018 132
rect 3894 78 3898 82
rect 3918 78 3922 82
rect 3926 78 3930 82
rect 3958 78 3962 82
rect 3918 68 3922 72
rect 4118 128 4122 132
rect 4102 108 4106 112
rect 4082 103 4086 107
rect 4089 103 4093 107
rect 4046 98 4050 102
rect 4070 98 4074 102
rect 3998 68 4002 72
rect 4038 68 4042 72
rect 3782 58 3786 62
rect 3806 58 3810 62
rect 3862 58 3866 62
rect 3910 58 3914 62
rect 3926 58 3930 62
rect 3942 58 3946 62
rect 3798 48 3802 52
rect 3806 48 3810 52
rect 3830 48 3834 52
rect 3854 48 3858 52
rect 3942 48 3946 52
rect 3774 28 3778 32
rect 3846 28 3850 32
rect 4030 58 4034 62
rect 3974 48 3978 52
rect 3990 48 3994 52
rect 4070 88 4074 92
rect 4222 198 4226 202
rect 4286 318 4290 322
rect 4294 288 4298 292
rect 4270 258 4274 262
rect 4254 238 4258 242
rect 4254 208 4258 212
rect 4246 198 4250 202
rect 4294 168 4298 172
rect 4358 318 4362 322
rect 4342 298 4346 302
rect 4350 298 4354 302
rect 4374 308 4378 312
rect 4390 328 4394 332
rect 4422 448 4426 452
rect 4438 438 4442 442
rect 4574 538 4578 542
rect 4534 528 4538 532
rect 4558 528 4562 532
rect 4550 498 4554 502
rect 4542 478 4546 482
rect 4574 478 4578 482
rect 4534 458 4538 462
rect 4558 458 4562 462
rect 4534 448 4538 452
rect 4478 438 4482 442
rect 4558 438 4562 442
rect 4518 408 4522 412
rect 4438 368 4442 372
rect 4502 368 4506 372
rect 4566 358 4570 362
rect 4406 348 4410 352
rect 4446 348 4450 352
rect 4494 348 4498 352
rect 4526 348 4530 352
rect 4550 348 4554 352
rect 4566 348 4570 352
rect 4534 338 4538 342
rect 4422 328 4426 332
rect 4478 328 4482 332
rect 4486 328 4490 332
rect 4414 308 4418 312
rect 4414 298 4418 302
rect 4446 298 4450 302
rect 4470 298 4474 302
rect 4518 298 4522 302
rect 4318 288 4322 292
rect 4350 288 4354 292
rect 4358 288 4362 292
rect 4318 258 4322 262
rect 4350 258 4354 262
rect 4382 258 4386 262
rect 4390 258 4394 262
rect 4406 258 4410 262
rect 4342 218 4346 222
rect 4302 158 4306 162
rect 4318 158 4322 162
rect 4230 148 4234 152
rect 4358 248 4362 252
rect 4478 288 4482 292
rect 4518 288 4522 292
rect 4486 278 4490 282
rect 4510 278 4514 282
rect 4502 268 4506 272
rect 4542 328 4546 332
rect 4558 308 4562 312
rect 4422 258 4426 262
rect 4414 228 4418 232
rect 4406 218 4410 222
rect 4382 178 4386 182
rect 4366 158 4370 162
rect 4454 238 4458 242
rect 4494 218 4498 222
rect 4446 188 4450 192
rect 4366 148 4370 152
rect 4398 148 4402 152
rect 4438 148 4442 152
rect 4270 138 4274 142
rect 4294 138 4298 142
rect 4190 108 4194 112
rect 4230 108 4234 112
rect 4238 108 4242 112
rect 4270 108 4274 112
rect 4342 138 4346 142
rect 4342 128 4346 132
rect 4358 128 4362 132
rect 4318 118 4322 122
rect 4326 108 4330 112
rect 4302 98 4306 102
rect 4158 88 4162 92
rect 4206 88 4210 92
rect 4286 88 4290 92
rect 4310 88 4314 92
rect 4414 138 4418 142
rect 4406 128 4410 132
rect 4454 158 4458 162
rect 4470 158 4474 162
rect 4470 138 4474 142
rect 4430 128 4434 132
rect 4422 118 4426 122
rect 4478 108 4482 112
rect 4430 98 4434 102
rect 4190 78 4194 82
rect 4246 78 4250 82
rect 4294 78 4298 82
rect 4334 78 4338 82
rect 4374 78 4378 82
rect 4054 68 4058 72
rect 4126 68 4130 72
rect 4182 68 4186 72
rect 4262 68 4266 72
rect 4134 58 4138 62
rect 4158 58 4162 62
rect 4046 38 4050 42
rect 4318 68 4322 72
rect 4366 68 4370 72
rect 4070 48 4074 52
rect 4182 48 4186 52
rect 4222 48 4226 52
rect 4278 48 4282 52
rect 4342 48 4346 52
rect 4390 68 4394 72
rect 4422 58 4426 62
rect 4382 48 4386 52
rect 4454 88 4458 92
rect 4446 78 4450 82
rect 4470 78 4474 82
rect 4438 68 4442 72
rect 4470 58 4474 62
rect 4478 58 4482 62
rect 4518 208 4522 212
rect 4542 198 4546 202
rect 4510 168 4514 172
rect 4542 158 4546 162
rect 4510 148 4514 152
rect 4542 138 4546 142
rect 4526 128 4530 132
rect 4526 118 4530 122
rect 4534 88 4538 92
rect 4550 68 4554 72
rect 4566 58 4570 62
rect 4494 48 4498 52
rect 4502 48 4506 52
rect 4574 48 4578 52
rect 4374 38 4378 42
rect 4406 38 4410 42
rect 4550 38 4554 42
rect 4574 38 4578 42
rect 4046 28 4050 32
rect 4054 28 4058 32
rect 4150 28 4154 32
rect 4494 28 4498 32
rect 3726 18 3730 22
rect 3950 18 3954 22
rect 4046 18 4050 22
rect 4166 18 4170 22
rect 3678 8 3682 12
rect 4262 8 4266 12
rect 2546 3 2550 7
rect 2553 3 2557 7
rect 3570 3 3574 7
rect 3577 3 3581 7
<< metal3 >>
rect 496 4403 498 4407
rect 502 4403 505 4407
rect 510 4403 512 4407
rect 1520 4403 1522 4407
rect 1526 4403 1529 4407
rect 1534 4403 1536 4407
rect 2544 4403 2546 4407
rect 2550 4403 2553 4407
rect 2558 4403 2560 4407
rect 3568 4403 3570 4407
rect 3574 4403 3577 4407
rect 3582 4403 3584 4407
rect 3634 4398 3686 4401
rect 3690 4398 3702 4401
rect 3754 4398 3758 4401
rect 3794 4398 3806 4401
rect 3826 4398 3830 4401
rect 3906 4398 3918 4401
rect 3954 4398 3966 4401
rect 3994 4398 4006 4401
rect 4010 4398 4014 4401
rect 4058 4398 4062 4401
rect 4130 4398 4158 4401
rect 4322 4398 4342 4401
rect 4378 4398 4430 4401
rect 1998 4392 2001 4398
rect 3942 4392 3945 4398
rect 4022 4392 4025 4398
rect 3986 4388 3998 4391
rect 4370 4388 4382 4391
rect 1586 4378 2022 4381
rect 3862 4381 3865 4388
rect 3862 4378 3934 4381
rect 4046 4381 4049 4388
rect 4046 4378 4118 4381
rect 4234 4378 4502 4381
rect 3766 4372 3769 4378
rect 1730 4368 1910 4371
rect 3422 4368 3478 4371
rect 3498 4368 3502 4371
rect 3598 4368 3670 4371
rect 4026 4368 4038 4371
rect 4042 4368 4190 4371
rect 4198 4371 4201 4378
rect 4198 4368 4278 4371
rect 4418 4368 4566 4371
rect 34 4358 190 4361
rect 774 4361 777 4368
rect 762 4358 777 4361
rect 794 4358 798 4361
rect 1510 4361 1513 4368
rect 3422 4362 3425 4368
rect 3598 4362 3601 4368
rect 1510 4358 1534 4361
rect 1706 4358 1734 4361
rect 1762 4358 1766 4361
rect 2150 4358 2158 4361
rect 2162 4358 2182 4361
rect 2186 4358 2238 4361
rect 2242 4358 2334 4361
rect 2426 4358 2462 4361
rect 2466 4358 2670 4361
rect 2674 4358 2678 4361
rect 2682 4358 2694 4361
rect 2978 4358 2990 4361
rect 2994 4358 3014 4361
rect 3314 4358 3334 4361
rect 3418 4358 3422 4361
rect 3442 4358 3486 4361
rect 3626 4358 3638 4361
rect 3722 4358 3750 4361
rect 3918 4358 3921 4368
rect 3942 4361 3945 4368
rect 3930 4358 3945 4361
rect 3974 4361 3977 4368
rect 3970 4358 3977 4361
rect 4146 4358 4150 4361
rect 4218 4358 4222 4361
rect 4346 4358 4358 4361
rect 4442 4358 4446 4361
rect -26 4351 -22 4352
rect -26 4348 6 4351
rect 74 4348 110 4351
rect 410 4348 462 4351
rect 546 4348 614 4351
rect 618 4348 638 4351
rect 726 4351 729 4358
rect 706 4348 729 4351
rect 746 4348 782 4351
rect 786 4348 798 4351
rect 942 4351 945 4358
rect 922 4348 974 4351
rect 1738 4348 1761 4351
rect 1758 4342 1761 4348
rect 1882 4348 1902 4351
rect 2018 4348 2158 4351
rect 2290 4348 2526 4351
rect 2530 4348 2606 4351
rect 2834 4348 3070 4351
rect 3254 4351 3257 4358
rect 3254 4348 3278 4351
rect 3414 4348 3422 4351
rect 3426 4348 3438 4351
rect 3470 4348 3478 4351
rect 3482 4348 3494 4351
rect 3510 4348 3518 4351
rect 3522 4348 3550 4351
rect 3562 4348 3694 4351
rect 3746 4348 3758 4351
rect 3782 4348 3790 4351
rect 3794 4348 3798 4351
rect 3814 4351 3817 4358
rect 4062 4352 4065 4358
rect 3814 4348 3822 4351
rect 3874 4348 3886 4351
rect 3938 4348 3945 4351
rect 3970 4348 3974 4351
rect 3978 4348 3998 4351
rect 4114 4348 4142 4351
rect 4170 4348 4182 4351
rect 4226 4348 4238 4351
rect 4326 4351 4329 4358
rect 4290 4348 4329 4351
rect 4362 4348 4390 4351
rect 4450 4348 4478 4351
rect 4490 4348 4494 4351
rect 4530 4348 4534 4351
rect 3942 4342 3945 4348
rect 4398 4342 4401 4348
rect 4510 4342 4513 4348
rect 4582 4342 4585 4348
rect 34 4338 54 4341
rect 106 4338 286 4341
rect 362 4338 582 4341
rect 586 4338 654 4341
rect 730 4338 942 4341
rect 946 4338 982 4341
rect 1086 4338 1134 4341
rect 1290 4338 1318 4341
rect 1506 4338 1710 4341
rect 2170 4338 2302 4341
rect 2658 4338 2678 4341
rect 2730 4338 2825 4341
rect 2890 4338 2942 4341
rect 2946 4338 2974 4341
rect 3234 4338 3238 4341
rect 3362 4338 3366 4341
rect 3474 4338 3486 4341
rect 3498 4338 3638 4341
rect 3642 4338 3686 4341
rect 3706 4338 3798 4341
rect 3802 4338 3894 4341
rect 3946 4338 3958 4341
rect 3970 4338 3990 4341
rect 4010 4338 4110 4341
rect 4114 4338 4198 4341
rect 4282 4338 4302 4341
rect 4330 4338 4334 4341
rect 4354 4338 4358 4341
rect 4410 4338 4414 4341
rect 4458 4338 4462 4341
rect 1086 4332 1089 4338
rect 82 4328 129 4331
rect 194 4328 270 4331
rect 594 4328 614 4331
rect 786 4328 790 4331
rect 802 4328 862 4331
rect 866 4328 873 4331
rect 938 4328 1086 4331
rect 1570 4328 1766 4331
rect 1770 4328 1798 4331
rect 1890 4328 1966 4331
rect 1970 4328 2078 4331
rect 2134 4331 2137 4338
rect 2422 4332 2425 4338
rect 2134 4328 2174 4331
rect 2210 4328 2214 4331
rect 2242 4328 2310 4331
rect 2598 4331 2601 4338
rect 2598 4328 2662 4331
rect 2822 4331 2825 4338
rect 3262 4332 3265 4338
rect 2822 4328 2966 4331
rect 3370 4328 3494 4331
rect 3506 4328 3646 4331
rect 3666 4328 3702 4331
rect 3730 4328 3806 4331
rect 3842 4328 3982 4331
rect 4058 4328 4086 4331
rect 4090 4328 4102 4331
rect 4122 4328 4126 4331
rect 4146 4328 4350 4331
rect 4362 4328 4390 4331
rect 4410 4328 4422 4331
rect 4434 4328 4558 4331
rect 126 4322 129 4328
rect 606 4318 614 4321
rect 618 4318 670 4321
rect 682 4318 686 4321
rect 738 4318 766 4321
rect 770 4318 838 4321
rect 926 4321 929 4328
rect 926 4318 958 4321
rect 1394 4318 1510 4321
rect 1698 4318 1766 4321
rect 1798 4321 1801 4328
rect 2406 4321 2409 4328
rect 2814 4322 2817 4328
rect 1798 4318 2201 4321
rect 2406 4318 2662 4321
rect 2674 4318 2809 4321
rect 3250 4318 3302 4321
rect 3450 4318 3614 4321
rect 3634 4318 3678 4321
rect 3690 4318 3806 4321
rect 3810 4318 3822 4321
rect 3962 4318 3990 4321
rect 3994 4318 4046 4321
rect 4066 4318 4078 4321
rect 4082 4318 4102 4321
rect 4146 4318 4166 4321
rect 4178 4318 4182 4321
rect 4202 4318 4270 4321
rect 4394 4318 4550 4321
rect 338 4308 350 4311
rect 682 4308 710 4311
rect 850 4308 934 4311
rect 2198 4311 2201 4318
rect 2198 4308 2710 4311
rect 2806 4311 2809 4318
rect 4054 4312 4057 4318
rect 2806 4308 2918 4311
rect 2938 4308 3038 4311
rect 3242 4308 3478 4311
rect 3482 4308 3542 4311
rect 3546 4308 3654 4311
rect 3714 4308 3718 4311
rect 3762 4308 3977 4311
rect 4138 4308 4302 4311
rect 4314 4308 4478 4311
rect 4490 4308 4518 4311
rect 4538 4308 4550 4311
rect 1000 4303 1002 4307
rect 1006 4303 1009 4307
rect 1014 4303 1016 4307
rect 2024 4303 2026 4307
rect 2030 4303 2033 4307
rect 2038 4303 2040 4307
rect 3048 4303 3050 4307
rect 3054 4303 3057 4307
rect 3062 4303 3064 4307
rect 3974 4302 3977 4308
rect 4080 4303 4082 4307
rect 4086 4303 4089 4307
rect 4094 4303 4096 4307
rect 354 4298 358 4301
rect 410 4298 438 4301
rect 2082 4298 2134 4301
rect 2466 4298 2774 4301
rect 2954 4298 2982 4301
rect 3090 4298 3262 4301
rect 3274 4298 3278 4301
rect 3338 4298 3446 4301
rect 3522 4298 3598 4301
rect 3602 4298 3670 4301
rect 3690 4298 3742 4301
rect 3754 4298 3782 4301
rect 3818 4298 3830 4301
rect 3882 4298 3918 4301
rect 3978 4298 4046 4301
rect 4106 4298 4134 4301
rect 4154 4298 4238 4301
rect 4250 4298 4422 4301
rect 4450 4298 4454 4301
rect 234 4288 414 4291
rect 418 4288 534 4291
rect 538 4288 630 4291
rect 634 4288 646 4291
rect 738 4288 846 4291
rect 962 4288 966 4291
rect 1914 4288 2022 4291
rect 2082 4288 2086 4291
rect 2098 4288 2118 4291
rect 2274 4288 2438 4291
rect 2442 4288 2454 4291
rect 2706 4288 2870 4291
rect 2914 4288 2990 4291
rect 2994 4288 3094 4291
rect 3234 4288 3358 4291
rect 3486 4291 3489 4298
rect 3394 4288 3489 4291
rect 3498 4288 3598 4291
rect 3622 4288 3630 4291
rect 3634 4288 3670 4291
rect 3682 4288 3774 4291
rect 3778 4288 3878 4291
rect 3890 4288 3902 4291
rect 3990 4288 3998 4291
rect 4002 4288 4038 4291
rect 4098 4288 4102 4291
rect 4118 4288 4126 4291
rect 4130 4288 4238 4291
rect 4302 4288 4310 4291
rect 4314 4288 4358 4291
rect 4366 4288 4374 4291
rect 4378 4288 4406 4291
rect 4522 4288 4574 4291
rect 354 4278 382 4281
rect 386 4278 454 4281
rect 810 4278 894 4281
rect 898 4278 918 4281
rect 922 4278 990 4281
rect 1002 4278 1046 4281
rect 1066 4278 1102 4281
rect 1154 4278 1270 4281
rect 1426 4278 1478 4281
rect 1722 4278 1846 4281
rect 1954 4278 2494 4281
rect 2498 4278 2718 4281
rect 2930 4278 2958 4281
rect 2962 4278 3126 4281
rect 3130 4278 3142 4281
rect 3330 4278 3398 4281
rect 3402 4278 3430 4281
rect 3442 4278 3654 4281
rect 3658 4278 3838 4281
rect 3842 4278 4102 4281
rect 4106 4278 4262 4281
rect 4266 4278 4430 4281
rect 4442 4278 4454 4281
rect 4466 4278 4502 4281
rect 4530 4278 4534 4281
rect 34 4268 54 4271
rect 146 4268 193 4271
rect 258 4268 294 4271
rect 298 4268 302 4271
rect 306 4268 534 4271
rect 546 4268 582 4271
rect 662 4271 665 4278
rect 618 4268 665 4271
rect 866 4268 870 4271
rect 938 4268 966 4271
rect 1042 4268 1118 4271
rect 1138 4268 1158 4271
rect 1186 4268 1222 4271
rect 1230 4268 1238 4271
rect 1242 4268 1254 4271
rect 1506 4268 1558 4271
rect 1574 4268 1593 4271
rect 110 4261 113 4268
rect 50 4258 113 4261
rect 190 4262 193 4268
rect 1574 4262 1577 4268
rect 1590 4262 1593 4268
rect 1818 4268 1822 4271
rect 1970 4268 2030 4271
rect 2114 4268 2230 4271
rect 2290 4268 2294 4271
rect 2330 4268 2334 4271
rect 2338 4268 2478 4271
rect 2482 4268 2526 4271
rect 2538 4268 2638 4271
rect 2842 4268 2846 4271
rect 2858 4268 2910 4271
rect 2938 4268 3014 4271
rect 3082 4268 3174 4271
rect 3370 4268 3454 4271
rect 3490 4268 3622 4271
rect 3626 4268 3654 4271
rect 3746 4268 3918 4271
rect 3994 4268 4294 4271
rect 4298 4268 4489 4271
rect 4498 4268 4526 4271
rect 302 4258 430 4261
rect 434 4258 590 4261
rect 834 4258 870 4261
rect 878 4258 902 4261
rect 962 4258 1030 4261
rect 1050 4258 1094 4261
rect 1106 4258 1134 4261
rect 1138 4258 1145 4261
rect 1202 4258 1206 4261
rect 1242 4258 1270 4261
rect 1350 4258 1358 4261
rect 1370 4258 1409 4261
rect 1490 4258 1510 4261
rect 1750 4261 1753 4268
rect 1594 4258 1886 4261
rect 2002 4258 2006 4261
rect 2302 4258 2318 4261
rect 2350 4258 2377 4261
rect 2410 4258 2414 4261
rect 2450 4258 2662 4261
rect 2686 4261 2689 4268
rect 2686 4258 2702 4261
rect 2766 4261 2769 4268
rect 2766 4258 2782 4261
rect 2830 4261 2833 4268
rect 2830 4258 2878 4261
rect 2954 4258 3102 4261
rect 3290 4258 3310 4261
rect 3362 4258 3406 4261
rect 3506 4258 3638 4261
rect 3666 4258 3710 4261
rect 3738 4258 3742 4261
rect 3746 4258 3750 4261
rect 3762 4258 3766 4261
rect 3778 4258 3782 4261
rect 3794 4258 3798 4261
rect 3818 4258 3822 4261
rect 3866 4258 3870 4261
rect 3958 4261 3961 4268
rect 3958 4258 3998 4261
rect 4010 4258 4014 4261
rect 4098 4258 4110 4261
rect 4130 4258 4150 4261
rect 4162 4258 4206 4261
rect 4258 4258 4286 4261
rect 4306 4258 4334 4261
rect 4354 4258 4470 4261
rect 4474 4258 4478 4261
rect 4486 4261 4489 4268
rect 4566 4262 4569 4268
rect 4486 4258 4534 4261
rect 302 4252 305 4258
rect 878 4252 881 4258
rect 1350 4252 1353 4258
rect 1406 4252 1409 4258
rect 2166 4252 2169 4258
rect 2302 4252 2305 4258
rect 2350 4252 2353 4258
rect 2374 4252 2377 4258
rect -26 4251 -22 4252
rect -26 4248 6 4251
rect 34 4248 206 4251
rect 266 4248 302 4251
rect 378 4248 518 4251
rect 538 4248 678 4251
rect 682 4248 710 4251
rect 810 4248 814 4251
rect 1058 4248 1126 4251
rect 1210 4248 1246 4251
rect 1978 4248 2150 4251
rect 2274 4248 2278 4251
rect 2442 4248 2502 4251
rect 2522 4248 2574 4251
rect 2602 4248 2630 4251
rect 2650 4248 2654 4251
rect 2674 4248 2750 4251
rect 2754 4248 2814 4251
rect 2818 4248 2846 4251
rect 2954 4248 2969 4251
rect 2986 4248 3046 4251
rect 3298 4248 3334 4251
rect 3358 4248 3374 4251
rect 3382 4248 3478 4251
rect 3506 4248 3534 4251
rect 3610 4248 3654 4251
rect 3658 4248 3678 4251
rect 3706 4248 3790 4251
rect 3910 4251 3913 4258
rect 3794 4248 4022 4251
rect 4074 4248 4166 4251
rect 4194 4248 4238 4251
rect 4274 4248 4278 4251
rect 4298 4248 4302 4251
rect 4354 4248 4382 4251
rect 4466 4248 4478 4251
rect 942 4242 945 4248
rect 370 4238 510 4241
rect 586 4238 670 4241
rect 674 4238 702 4241
rect 754 4238 806 4241
rect 962 4238 966 4241
rect 1122 4238 1150 4241
rect 1254 4241 1257 4248
rect 1254 4238 1462 4241
rect 1482 4238 1606 4241
rect 1786 4238 1806 4241
rect 1986 4238 1990 4241
rect 2206 4241 2209 4248
rect 2966 4242 2969 4248
rect 3358 4242 3361 4248
rect 3382 4242 3385 4248
rect 2186 4238 2209 4241
rect 2250 4238 2310 4241
rect 2458 4238 2478 4241
rect 2490 4238 2526 4241
rect 2546 4238 2598 4241
rect 2666 4238 2694 4241
rect 2794 4238 2846 4241
rect 3306 4238 3326 4241
rect 3402 4238 3422 4241
rect 3534 4241 3537 4248
rect 3534 4238 3966 4241
rect 3970 4238 4134 4241
rect 4138 4238 4190 4241
rect 4354 4238 4358 4241
rect 4482 4238 4510 4241
rect 434 4228 454 4231
rect 466 4228 470 4231
rect 482 4228 598 4231
rect 634 4228 790 4231
rect 858 4228 1246 4231
rect 1250 4228 1278 4231
rect 1666 4228 1702 4231
rect 1898 4228 2078 4231
rect 2170 4228 2254 4231
rect 2258 4228 2286 4231
rect 2290 4228 2390 4231
rect 2418 4228 2486 4231
rect 2494 4228 2614 4231
rect 2682 4228 2742 4231
rect 2746 4228 2790 4231
rect 2842 4228 2918 4231
rect 2922 4228 2942 4231
rect 3282 4228 3422 4231
rect 3426 4228 3462 4231
rect 3478 4231 3481 4238
rect 3478 4228 3622 4231
rect 3626 4228 3750 4231
rect 3826 4228 3830 4231
rect 3850 4228 3894 4231
rect 3922 4228 3974 4231
rect 4082 4228 4126 4231
rect 4258 4228 4302 4231
rect 4322 4228 4326 4231
rect 4410 4228 4486 4231
rect 4490 4228 4574 4231
rect 790 4221 793 4228
rect 2494 4222 2497 4228
rect 790 4218 886 4221
rect 914 4218 1086 4221
rect 1114 4218 1222 4221
rect 1498 4218 1518 4221
rect 1522 4218 1678 4221
rect 1818 4218 1966 4221
rect 2018 4218 2038 4221
rect 2122 4218 2246 4221
rect 2250 4218 2257 4221
rect 2594 4218 2806 4221
rect 2850 4218 3054 4221
rect 3266 4218 3310 4221
rect 3378 4218 3510 4221
rect 3714 4218 3718 4221
rect 3762 4218 4454 4221
rect 4570 4218 4590 4221
rect 270 4212 273 4218
rect 842 4208 1238 4211
rect 1826 4208 1998 4211
rect 2034 4208 2206 4211
rect 2218 4208 2318 4211
rect 2338 4208 2534 4211
rect 2666 4208 2678 4211
rect 2722 4208 2798 4211
rect 2802 4208 2894 4211
rect 2930 4208 3326 4211
rect 3450 4208 3510 4211
rect 3818 4208 3854 4211
rect 3882 4208 4014 4211
rect 4018 4208 4102 4211
rect 4106 4208 4142 4211
rect 4266 4208 4302 4211
rect 4306 4208 4398 4211
rect 4442 4208 4518 4211
rect 4522 4208 4542 4211
rect 4546 4208 4550 4211
rect 496 4203 498 4207
rect 502 4203 505 4207
rect 510 4203 512 4207
rect 1520 4203 1522 4207
rect 1526 4203 1529 4207
rect 1534 4203 1536 4207
rect 2544 4203 2546 4207
rect 2550 4203 2553 4207
rect 2558 4203 2560 4207
rect 3568 4203 3570 4207
rect 3574 4203 3577 4207
rect 3582 4203 3584 4207
rect 178 4198 230 4201
rect 626 4198 838 4201
rect 1098 4198 1214 4201
rect 1842 4198 2102 4201
rect 2186 4198 2262 4201
rect 2266 4198 2294 4201
rect 2330 4198 2537 4201
rect 2714 4198 2950 4201
rect 3762 4198 3878 4201
rect 3946 4198 3966 4201
rect 3978 4198 4246 4201
rect 4250 4198 4278 4201
rect 4282 4198 4294 4201
rect 4298 4198 4390 4201
rect 258 4188 366 4191
rect 446 4191 449 4198
rect 446 4188 542 4191
rect 706 4188 870 4191
rect 942 4188 950 4191
rect 954 4188 1126 4191
rect 1138 4188 1166 4191
rect 1790 4188 1798 4191
rect 1802 4188 1942 4191
rect 2134 4188 2142 4191
rect 2146 4188 2238 4191
rect 2282 4188 2286 4191
rect 2294 4191 2297 4198
rect 2294 4188 2382 4191
rect 2418 4188 2462 4191
rect 2534 4191 2537 4198
rect 2534 4188 2678 4191
rect 2770 4188 2774 4191
rect 2794 4188 3158 4191
rect 3246 4191 3249 4198
rect 3246 4188 3358 4191
rect 3890 4188 4118 4191
rect 4122 4188 4142 4191
rect 4434 4188 4502 4191
rect 138 4178 430 4181
rect 694 4181 697 4188
rect 694 4178 710 4181
rect 882 4178 1038 4181
rect 1050 4178 1094 4181
rect 1794 4178 1814 4181
rect 1938 4178 2094 4181
rect 2098 4178 2238 4181
rect 2246 4181 2249 4188
rect 2246 4178 2326 4181
rect 2390 4178 2398 4181
rect 2402 4178 2502 4181
rect 2618 4178 2798 4181
rect 2810 4178 3118 4181
rect 3250 4178 3278 4181
rect 3282 4178 3302 4181
rect 3306 4178 3494 4181
rect 3874 4178 3974 4181
rect 4002 4178 4038 4181
rect 4042 4178 4174 4181
rect 4178 4178 4230 4181
rect 4234 4178 4334 4181
rect 4338 4178 4414 4181
rect 4418 4178 4430 4181
rect 258 4168 326 4171
rect 698 4168 806 4171
rect 810 4168 958 4171
rect 970 4168 1254 4171
rect 1286 4171 1289 4178
rect 1286 4168 1494 4171
rect 1926 4171 1929 4178
rect 1926 4168 2006 4171
rect 2010 4168 2046 4171
rect 2050 4168 2182 4171
rect 2210 4168 2414 4171
rect 2458 4168 2486 4171
rect 2490 4168 2510 4171
rect 2514 4168 2678 4171
rect 2834 4168 2990 4171
rect 3146 4168 3230 4171
rect 3234 4168 3286 4171
rect 3350 4168 3638 4171
rect 3642 4168 3678 4171
rect 3698 4168 3870 4171
rect 3966 4168 4022 4171
rect 4146 4168 4158 4171
rect 4162 4168 4182 4171
rect 4338 4168 4406 4171
rect 4630 4171 4634 4172
rect 4562 4168 4634 4171
rect 114 4158 174 4161
rect 218 4158 246 4161
rect 322 4158 382 4161
rect 562 4158 566 4161
rect 610 4158 702 4161
rect 722 4158 726 4161
rect 794 4158 817 4161
rect 930 4158 1070 4161
rect 1146 4158 1238 4161
rect 1262 4161 1265 4168
rect 2430 4162 2433 4168
rect 2686 4162 2689 4168
rect 3270 4162 3273 4168
rect 3350 4162 3353 4168
rect 1262 4158 1302 4161
rect 1322 4158 1334 4161
rect 1442 4158 1446 4161
rect 1626 4158 1750 4161
rect 1754 4158 1790 4161
rect 1810 4158 2206 4161
rect 2218 4158 2222 4161
rect 2410 4158 2422 4161
rect 2530 4158 2534 4161
rect 2538 4158 2606 4161
rect 2874 4158 2934 4161
rect 2938 4158 2942 4161
rect 3418 4158 3446 4161
rect 3450 4158 3526 4161
rect 3530 4158 3662 4161
rect 3762 4158 3830 4161
rect 3910 4161 3913 4168
rect 3950 4161 3953 4168
rect 3910 4158 3953 4161
rect 3966 4162 3969 4168
rect 4042 4158 4062 4161
rect 4114 4158 4118 4161
rect 4134 4161 4137 4168
rect 4134 4158 4142 4161
rect 4162 4158 4206 4161
rect 4254 4161 4257 4168
rect 4254 4158 4262 4161
rect 4286 4161 4289 4168
rect 4286 4158 4310 4161
rect 4370 4158 4382 4161
rect 4446 4161 4449 4168
rect 4402 4158 4449 4161
rect 4462 4158 4510 4161
rect 814 4152 817 4158
rect 2334 4152 2337 4158
rect -26 4151 -22 4152
rect -26 4148 6 4151
rect 90 4148 446 4151
rect 634 4148 638 4151
rect 706 4148 734 4151
rect 738 4148 774 4151
rect 778 4148 798 4151
rect 858 4148 870 4151
rect 1018 4148 1062 4151
rect 1082 4148 1126 4151
rect 1410 4148 1670 4151
rect 1674 4148 1694 4151
rect 1702 4148 1718 4151
rect 1850 4148 1854 4151
rect 1866 4148 1926 4151
rect 1930 4148 1942 4151
rect 2018 4148 2022 4151
rect 2026 4148 2070 4151
rect 2074 4148 2110 4151
rect 2114 4148 2158 4151
rect 2222 4148 2254 4151
rect 2346 4148 2350 4151
rect 2442 4148 2462 4151
rect 2486 4151 2489 4158
rect 2486 4148 2502 4151
rect 2586 4148 2726 4151
rect 2798 4151 2801 4158
rect 2846 4151 2849 4158
rect 2798 4148 2849 4151
rect 2862 4151 2865 4158
rect 2862 4148 2878 4151
rect 2906 4148 2942 4151
rect 2946 4148 3022 4151
rect 3138 4148 3150 4151
rect 3226 4148 3302 4151
rect 3330 4148 3350 4151
rect 3498 4148 3558 4151
rect 3674 4148 3766 4151
rect 3818 4148 3982 4151
rect 3986 4148 4006 4151
rect 4066 4148 4198 4151
rect 4202 4148 4214 4151
rect 4218 4148 4358 4151
rect 4362 4148 4438 4151
rect 4462 4151 4465 4158
rect 4450 4148 4465 4151
rect 4474 4148 4478 4151
rect 4530 4148 4558 4151
rect 4598 4151 4601 4158
rect 4630 4151 4634 4152
rect 4594 4148 4634 4151
rect 34 4138 54 4141
rect 234 4138 270 4141
rect 290 4138 302 4141
rect 314 4138 334 4141
rect 338 4138 542 4141
rect 546 4138 670 4141
rect 674 4138 726 4141
rect 730 4138 750 4141
rect 810 4138 854 4141
rect 898 4138 910 4141
rect 1050 4138 1054 4141
rect 1074 4138 1086 4141
rect 1210 4138 1318 4141
rect 1402 4138 1430 4141
rect 1702 4141 1705 4148
rect 1438 4138 1705 4141
rect 1766 4141 1769 4148
rect 2222 4142 2225 4148
rect 1714 4138 1769 4141
rect 1778 4138 1822 4141
rect 1826 4138 1838 4141
rect 1842 4138 1886 4141
rect 1914 4138 1918 4141
rect 1970 4138 2086 4141
rect 2314 4138 2366 4141
rect 2578 4138 2598 4141
rect 2766 4141 2769 4148
rect 2766 4138 2814 4141
rect 2818 4138 2998 4141
rect 3042 4138 3190 4141
rect 3194 4138 3214 4141
rect 3274 4138 3286 4141
rect 3306 4138 3374 4141
rect 3434 4138 3438 4141
rect 3458 4138 3470 4141
rect 3474 4138 3502 4141
rect 3738 4138 3758 4141
rect 3762 4138 3854 4141
rect 3858 4138 3918 4141
rect 3922 4138 3950 4141
rect 3954 4138 4254 4141
rect 4258 4138 4270 4141
rect 4274 4138 4318 4141
rect 4330 4138 4377 4141
rect 4386 4138 4422 4141
rect 4434 4138 4454 4141
rect 1438 4132 1441 4138
rect 202 4128 222 4131
rect 242 4128 246 4131
rect 298 4128 326 4131
rect 354 4128 398 4131
rect 498 4128 558 4131
rect 562 4128 638 4131
rect 642 4128 654 4131
rect 826 4128 990 4131
rect 1026 4128 1070 4131
rect 1074 4128 1182 4131
rect 1250 4128 1302 4131
rect 1474 4128 1518 4131
rect 1522 4128 1566 4131
rect 1774 4131 1777 4138
rect 1762 4128 1777 4131
rect 1970 4128 1974 4131
rect 2082 4128 2086 4131
rect 2090 4128 2118 4131
rect 2146 4128 2182 4131
rect 2250 4128 2254 4131
rect 2354 4128 2630 4131
rect 2682 4128 2846 4131
rect 2878 4128 2894 4131
rect 2914 4128 3038 4131
rect 3170 4128 3198 4131
rect 3202 4128 3230 4131
rect 3234 4128 3302 4131
rect 3314 4128 3422 4131
rect 3426 4128 3574 4131
rect 3578 4128 3710 4131
rect 3770 4128 3894 4131
rect 3898 4128 3918 4131
rect 3930 4128 4262 4131
rect 4298 4128 4334 4131
rect 4338 4128 4366 4131
rect 4374 4131 4377 4138
rect 4374 4128 4489 4131
rect 182 4121 185 4128
rect 286 4121 289 4128
rect 182 4118 289 4121
rect 434 4118 574 4121
rect 578 4118 606 4121
rect 610 4118 718 4121
rect 722 4118 726 4121
rect 818 4118 878 4121
rect 946 4118 974 4121
rect 978 4118 1030 4121
rect 1042 4118 1126 4121
rect 1130 4118 1158 4121
rect 1326 4121 1329 4128
rect 1326 4118 1694 4121
rect 1742 4121 1745 4128
rect 2878 4122 2881 4128
rect 1742 4118 1977 4121
rect 1986 4118 2142 4121
rect 2178 4118 2262 4121
rect 2354 4118 2358 4121
rect 2362 4118 2582 4121
rect 2602 4118 2654 4121
rect 2666 4118 2806 4121
rect 2882 4118 3078 4121
rect 3430 4118 3438 4121
rect 3442 4118 3486 4121
rect 3506 4118 3582 4121
rect 3586 4118 3678 4121
rect 3686 4118 3814 4121
rect 3926 4121 3929 4128
rect 4486 4122 4489 4128
rect 3866 4118 3929 4121
rect 4034 4118 4054 4121
rect 4058 4118 4126 4121
rect 4130 4118 4174 4121
rect 4178 4118 4438 4121
rect 4442 4118 4478 4121
rect 4562 4118 4598 4121
rect 1974 4112 1977 4118
rect 3686 4112 3689 4118
rect 210 4108 318 4111
rect 386 4108 534 4111
rect 602 4108 686 4111
rect 690 4108 822 4111
rect 962 4108 990 4111
rect 1418 4108 1430 4111
rect 1690 4108 1718 4111
rect 1722 4108 1790 4111
rect 2226 4108 2238 4111
rect 2274 4108 2398 4111
rect 2426 4108 2478 4111
rect 2506 4108 2518 4111
rect 2522 4108 2686 4111
rect 2690 4108 2718 4111
rect 2754 4108 2910 4111
rect 3074 4108 3302 4111
rect 3338 4108 3550 4111
rect 3826 4108 3918 4111
rect 3930 4108 3942 4111
rect 3946 4108 4038 4111
rect 4106 4108 4134 4111
rect 4186 4108 4206 4111
rect 4226 4108 4302 4111
rect 4306 4108 4374 4111
rect 4442 4108 4470 4111
rect 4474 4108 4558 4111
rect 4562 4108 4590 4111
rect 1000 4103 1002 4107
rect 1006 4103 1009 4107
rect 1014 4103 1016 4107
rect 2024 4103 2026 4107
rect 2030 4103 2033 4107
rect 2038 4103 2040 4107
rect 3048 4103 3050 4107
rect 3054 4103 3057 4107
rect 3062 4103 3064 4107
rect 4080 4103 4082 4107
rect 4086 4103 4089 4107
rect 4094 4103 4096 4107
rect 114 4098 142 4101
rect 186 4098 294 4101
rect 338 4098 470 4101
rect 722 4098 758 4101
rect 834 4098 966 4101
rect 1266 4098 1286 4101
rect 1490 4098 1550 4101
rect 1642 4098 1654 4101
rect 1706 4098 1742 4101
rect 2306 4098 2350 4101
rect 2362 4098 2382 4101
rect 2386 4098 2558 4101
rect 2658 4098 2854 4101
rect 2946 4098 2966 4101
rect 3074 4098 3102 4101
rect 3362 4098 3558 4101
rect 3578 4098 3662 4101
rect 3666 4098 3782 4101
rect 3818 4098 3990 4101
rect 4106 4098 4150 4101
rect 4218 4098 4238 4101
rect 4298 4098 4318 4101
rect 4458 4098 4510 4101
rect 4514 4098 4542 4101
rect 226 4088 350 4091
rect 450 4088 470 4091
rect 474 4088 702 4091
rect 770 4088 782 4091
rect 786 4088 830 4091
rect 1202 4088 1270 4091
rect 1282 4088 1326 4091
rect 1330 4088 1414 4091
rect 1546 4088 1638 4091
rect 1770 4088 2910 4091
rect 3602 4088 3630 4091
rect 3650 4088 3686 4091
rect 3734 4088 3798 4091
rect 3850 4088 3982 4091
rect 4114 4088 4126 4091
rect 4138 4088 4390 4091
rect 4394 4088 4422 4091
rect 4474 4088 4534 4091
rect 178 4078 182 4081
rect 198 4078 230 4081
rect 322 4078 382 4081
rect 530 4078 606 4081
rect 718 4081 721 4088
rect 690 4078 721 4081
rect 754 4078 766 4081
rect 770 4078 798 4081
rect 826 4078 846 4081
rect 890 4078 894 4081
rect 982 4081 985 4088
rect 962 4078 985 4081
rect 1002 4078 1089 4081
rect 1306 4078 1518 4081
rect 1618 4078 1678 4081
rect 1770 4078 1782 4081
rect 1786 4078 1814 4081
rect 1818 4078 1846 4081
rect 2002 4078 2110 4081
rect 2122 4078 2182 4081
rect 2186 4078 2230 4081
rect 2234 4078 2254 4081
rect 2258 4078 2342 4081
rect 2450 4078 2462 4081
rect 2474 4078 2526 4081
rect 2658 4078 2734 4081
rect 2890 4078 3038 4081
rect 3174 4081 3177 4088
rect 3090 4078 3177 4081
rect 3234 4078 3262 4081
rect 3366 4081 3369 4088
rect 3734 4082 3737 4088
rect 3266 4078 3446 4081
rect 3450 4078 3478 4081
rect 3482 4078 3510 4081
rect 3514 4078 3566 4081
rect 3666 4078 3678 4081
rect 3682 4078 3734 4081
rect 3786 4078 3814 4081
rect 3874 4078 3910 4081
rect 3922 4078 4110 4081
rect 4114 4078 4118 4081
rect 4130 4078 4398 4081
rect 4402 4078 4430 4081
rect 4474 4078 4478 4081
rect 4482 4078 4510 4081
rect 4514 4078 4521 4081
rect 4538 4078 4542 4081
rect 198 4072 201 4078
rect 1086 4072 1089 4078
rect 186 4068 198 4071
rect 218 4068 238 4071
rect 242 4068 310 4071
rect 338 4068 374 4071
rect 538 4068 830 4071
rect 834 4068 838 4071
rect 850 4068 902 4071
rect 906 4068 934 4071
rect 978 4068 990 4071
rect 1090 4068 1134 4071
rect 1530 4068 1662 4071
rect 1714 4068 1774 4071
rect 1810 4068 1838 4071
rect 1846 4071 1849 4078
rect 2054 4072 2057 4078
rect 2638 4072 2641 4078
rect 1846 4068 1870 4071
rect 2066 4068 2190 4071
rect 2338 4068 2358 4071
rect 2450 4068 2590 4071
rect 2598 4068 2622 4071
rect 2666 4068 2750 4071
rect 2990 4068 3238 4071
rect 3242 4068 3262 4071
rect 3306 4068 3329 4071
rect 3434 4068 3454 4071
rect 3530 4068 3646 4071
rect 3650 4068 3750 4071
rect 3754 4068 3766 4071
rect 3770 4068 3798 4071
rect 3890 4068 3998 4071
rect 4010 4068 4046 4071
rect 4170 4068 4198 4071
rect 4234 4068 4238 4071
rect 4266 4068 4286 4071
rect 4290 4068 4318 4071
rect 4322 4068 4326 4071
rect 4362 4068 4366 4071
rect 4370 4068 4502 4071
rect 4506 4068 4550 4071
rect 4554 4068 4566 4071
rect 1502 4062 1505 4068
rect 2598 4062 2601 4068
rect 2990 4062 2993 4068
rect 3326 4062 3329 4068
rect 4134 4062 4137 4068
rect 4142 4062 4145 4068
rect 194 4058 206 4061
rect 210 4058 230 4061
rect 242 4058 366 4061
rect 370 4058 478 4061
rect 578 4058 598 4061
rect 670 4058 782 4061
rect 834 4058 918 4061
rect 946 4058 950 4061
rect 1066 4058 1302 4061
rect 1418 4058 1486 4061
rect 1490 4058 1494 4061
rect 1614 4058 1742 4061
rect 1746 4058 1782 4061
rect 1794 4058 1854 4061
rect 1866 4058 1881 4061
rect 1922 4058 1958 4061
rect 1962 4058 2006 4061
rect 2074 4058 2286 4061
rect 2338 4058 2342 4061
rect 2346 4058 2398 4061
rect 2402 4058 2438 4061
rect 2458 4058 2486 4061
rect 2778 4058 2814 4061
rect 2826 4058 2830 4061
rect 2890 4058 2894 4061
rect 2922 4058 2990 4061
rect 3074 4058 3126 4061
rect 3130 4058 3182 4061
rect 3210 4058 3225 4061
rect 3258 4058 3278 4061
rect 3394 4058 3446 4061
rect 3450 4058 3502 4061
rect 3570 4058 3582 4061
rect 3586 4058 3614 4061
rect 3674 4058 3838 4061
rect 3842 4058 3894 4061
rect 3978 4058 4078 4061
rect 4218 4058 4254 4061
rect 4274 4058 4294 4061
rect 4298 4058 4318 4061
rect 4490 4058 4510 4061
rect 4514 4058 4574 4061
rect 250 4048 334 4051
rect 346 4048 358 4051
rect 490 4048 630 4051
rect 670 4051 673 4058
rect 1614 4052 1617 4058
rect 1878 4052 1881 4058
rect 2710 4052 2713 4058
rect 3222 4052 3225 4058
rect 666 4048 673 4051
rect 762 4048 766 4051
rect 786 4048 790 4051
rect 810 4048 862 4051
rect 930 4048 1046 4051
rect 1498 4048 1505 4051
rect 1954 4048 1974 4051
rect 2078 4048 2086 4051
rect 2090 4048 2110 4051
rect 2138 4048 2150 4051
rect 2154 4048 2206 4051
rect 2330 4048 2414 4051
rect 2422 4048 2430 4051
rect 2434 4048 2494 4051
rect 2514 4048 2518 4051
rect 2618 4048 2622 4051
rect 2634 4048 2694 4051
rect 2762 4048 2782 4051
rect 2786 4048 2862 4051
rect 2866 4048 2894 4051
rect 3266 4048 3318 4051
rect 3546 4048 3598 4051
rect 3602 4048 3646 4051
rect 3666 4048 3750 4051
rect 3778 4048 3790 4051
rect 3810 4048 3870 4051
rect 3934 4051 3937 4058
rect 3934 4048 4014 4051
rect 4034 4048 4094 4051
rect 4266 4048 4273 4051
rect 462 4041 465 4048
rect 1502 4042 1505 4048
rect 426 4038 465 4041
rect 714 4038 846 4041
rect 858 4038 886 4041
rect 890 4038 1094 4041
rect 1106 4038 1294 4041
rect 1466 4038 1494 4041
rect 1826 4038 1926 4041
rect 1934 4041 1937 4048
rect 1934 4038 1950 4041
rect 1954 4038 1998 4041
rect 2002 4038 2006 4041
rect 2114 4038 2134 4041
rect 2210 4038 2222 4041
rect 2306 4038 2358 4041
rect 2378 4038 2390 4041
rect 2418 4038 2430 4041
rect 2518 4041 2521 4048
rect 2590 4041 2593 4048
rect 2518 4038 2593 4041
rect 2746 4038 2782 4041
rect 2810 4038 2838 4041
rect 2842 4038 2910 4041
rect 3046 4041 3049 4048
rect 4270 4042 4273 4048
rect 4322 4048 4366 4051
rect 4370 4048 4406 4051
rect 4454 4051 4457 4058
rect 4426 4048 4457 4051
rect 4498 4048 4510 4051
rect 4530 4048 4566 4051
rect 4630 4051 4634 4052
rect 4570 4048 4634 4051
rect 2938 4038 3049 4041
rect 3202 4038 3222 4041
rect 3226 4038 3310 4041
rect 3578 4038 3590 4041
rect 3634 4038 3710 4041
rect 3714 4038 3902 4041
rect 3906 4038 3934 4041
rect 3962 4038 3998 4041
rect 4002 4038 4046 4041
rect 4286 4041 4289 4048
rect 4286 4038 4350 4041
rect 4354 4038 4374 4041
rect 4378 4038 4446 4041
rect 4470 4041 4473 4048
rect 4470 4038 4534 4041
rect 4542 4038 4598 4041
rect 4542 4032 4545 4038
rect 314 4028 326 4031
rect 330 4028 406 4031
rect 410 4028 526 4031
rect 530 4028 534 4031
rect 538 4028 558 4031
rect 770 4028 1110 4031
rect 1306 4028 1846 4031
rect 1850 4028 2294 4031
rect 2298 4028 2678 4031
rect 2722 4028 2750 4031
rect 3706 4028 3726 4031
rect 3730 4028 3734 4031
rect 3834 4028 3918 4031
rect 3922 4028 3950 4031
rect 3986 4028 4222 4031
rect 4562 4028 4598 4031
rect 42 4018 70 4021
rect 114 4018 254 4021
rect 258 4018 342 4021
rect 346 4018 358 4021
rect 378 4018 566 4021
rect 734 4021 737 4028
rect 734 4018 1102 4021
rect 1114 4018 1390 4021
rect 1394 4018 1486 4021
rect 1610 4018 1822 4021
rect 1930 4018 2126 4021
rect 2130 4018 2206 4021
rect 2210 4018 2222 4021
rect 2474 4018 2582 4021
rect 2586 4018 2702 4021
rect 2810 4018 2926 4021
rect 3738 4018 3814 4021
rect 3866 4018 3926 4021
rect 3930 4018 3966 4021
rect 3994 4018 3998 4021
rect 4122 4018 4158 4021
rect 250 4008 270 4011
rect 274 4008 286 4011
rect 322 4008 486 4011
rect 706 4008 910 4011
rect 1786 4008 1982 4011
rect 2114 4008 2446 4011
rect 2626 4008 2702 4011
rect 2802 4008 3030 4011
rect 3626 4008 3958 4011
rect 3962 4008 4062 4011
rect 4154 4008 4166 4011
rect 496 4003 498 4007
rect 502 4003 505 4007
rect 510 4003 512 4007
rect 1398 4002 1401 4008
rect 1520 4003 1522 4007
rect 1526 4003 1529 4007
rect 1534 4003 1536 4007
rect 2544 4003 2546 4007
rect 2550 4003 2553 4007
rect 2558 4003 2560 4007
rect 3568 4003 3570 4007
rect 3574 4003 3577 4007
rect 3582 4003 3584 4007
rect 794 3998 1030 4001
rect 1546 3998 1918 4001
rect 1922 3998 2534 4001
rect 2570 3998 2670 4001
rect 2674 3998 2750 4001
rect 2754 3998 2830 4001
rect 2898 3998 3214 4001
rect 3810 3998 4030 4001
rect 4074 3998 4390 4001
rect 178 3988 254 3991
rect 258 3988 302 3991
rect 306 3988 350 3991
rect 490 3988 510 3991
rect 626 3988 702 3991
rect 858 3988 1038 3991
rect 1322 3988 1649 3991
rect 1770 3988 1774 3991
rect 1814 3988 1822 3991
rect 1826 3988 1958 3991
rect 1986 3988 1990 3991
rect 2122 3988 2918 3991
rect 3002 3988 3038 3991
rect 3042 3988 3086 3991
rect 3090 3988 3094 3991
rect 3274 3988 3414 3991
rect 3514 3988 3750 3991
rect 3754 3988 4006 3991
rect 4010 3988 4062 3991
rect 4434 3988 4521 3991
rect 1646 3982 1649 3988
rect 170 3978 174 3981
rect 458 3978 486 3981
rect 898 3978 1542 3981
rect 1650 3978 1918 3981
rect 2086 3978 2214 3981
rect 2218 3978 2422 3981
rect 2426 3978 2454 3981
rect 2622 3978 2790 3981
rect 2834 3978 3406 3981
rect 3414 3981 3417 3988
rect 4518 3982 4521 3988
rect 3414 3978 3462 3981
rect 3554 3978 3566 3981
rect 3618 3978 3694 3981
rect 3698 3978 3790 3981
rect 3802 3978 3838 3981
rect 3970 3978 4022 3981
rect 4026 3978 4166 3981
rect 4218 3978 4350 3981
rect 4354 3978 4494 3981
rect -26 3971 -22 3972
rect -26 3968 6 3971
rect 350 3971 353 3978
rect 274 3968 353 3971
rect 394 3968 446 3971
rect 634 3968 646 3971
rect 650 3968 833 3971
rect 842 3968 1662 3971
rect 2086 3971 2089 3978
rect 2622 3972 2625 3978
rect 1666 3968 2089 3971
rect 2098 3968 2110 3971
rect 2154 3968 2318 3971
rect 2354 3968 2598 3971
rect 2690 3968 2822 3971
rect 2834 3968 3022 3971
rect 3026 3968 3110 3971
rect 3338 3968 3406 3971
rect 3426 3968 3446 3971
rect 3594 3968 3758 3971
rect 3762 3968 3942 3971
rect 4250 3968 4358 3971
rect 4434 3968 4462 3971
rect 4542 3971 4545 3978
rect 4530 3968 4545 3971
rect 338 3958 486 3961
rect 830 3961 833 3968
rect 830 3958 838 3961
rect 842 3958 894 3961
rect 898 3958 950 3961
rect 1418 3958 1518 3961
rect 1538 3958 1782 3961
rect 1810 3958 1814 3961
rect 1906 3958 1910 3961
rect 1970 3958 1982 3961
rect 2018 3958 2174 3961
rect 2194 3958 2198 3961
rect 2210 3958 2238 3961
rect 2282 3958 2630 3961
rect 2650 3958 2697 3961
rect -26 3948 -22 3952
rect 58 3948 126 3951
rect 298 3948 342 3951
rect 426 3948 550 3951
rect 554 3948 790 3951
rect 818 3948 830 3951
rect 954 3948 1054 3951
rect 1058 3948 1158 3951
rect 1266 3948 1270 3951
rect 1298 3948 1342 3951
rect 1374 3951 1377 3958
rect 2694 3952 2697 3958
rect 2810 3958 2862 3961
rect 2866 3958 2886 3961
rect 3142 3961 3145 3968
rect 2890 3958 3145 3961
rect 3362 3958 3550 3961
rect 3610 3958 3622 3961
rect 3730 3958 3806 3961
rect 3850 3958 3854 3961
rect 3882 3958 3894 3961
rect 3982 3961 3985 3968
rect 4022 3961 4025 3968
rect 3982 3958 4142 3961
rect 4250 3958 4254 3961
rect 4450 3958 4470 3961
rect 4482 3958 4534 3961
rect 4538 3958 4582 3961
rect 4594 3958 4598 3961
rect 4630 3961 4634 3962
rect 4602 3958 4634 3961
rect 1374 3948 1406 3951
rect 1526 3948 1662 3951
rect 1666 3948 1998 3951
rect 2002 3948 2006 3951
rect 2098 3948 2134 3951
rect 2186 3948 2190 3951
rect 2362 3948 2382 3951
rect 2530 3948 2534 3951
rect 2538 3948 2550 3951
rect 2734 3951 2737 3958
rect 3902 3952 3905 3958
rect 2734 3948 2782 3951
rect 2930 3948 2934 3951
rect -26 3941 -23 3948
rect -26 3938 70 3941
rect 206 3941 209 3948
rect 262 3941 265 3948
rect 206 3938 265 3941
rect 290 3938 294 3941
rect 298 3938 358 3941
rect 374 3941 377 3948
rect 374 3938 398 3941
rect 414 3941 417 3948
rect 402 3938 417 3941
rect 522 3938 617 3941
rect 642 3938 766 3941
rect 802 3938 806 3941
rect 1526 3941 1529 3948
rect 1042 3938 1529 3941
rect 1786 3938 1806 3941
rect 1810 3938 1814 3941
rect 1850 3938 1854 3941
rect 1858 3938 1894 3941
rect 1906 3938 2326 3941
rect 2330 3938 2342 3941
rect 2554 3938 2614 3941
rect 2618 3938 2766 3941
rect 2838 3941 2841 3948
rect 3274 3948 3286 3951
rect 3322 3948 3334 3951
rect 3338 3948 3382 3951
rect 3410 3948 3441 3951
rect 3438 3942 3441 3948
rect 3470 3948 3582 3951
rect 3590 3948 3606 3951
rect 3658 3948 3718 3951
rect 3730 3948 3854 3951
rect 3874 3948 3878 3951
rect 3890 3948 3894 3951
rect 3926 3951 3929 3958
rect 3906 3948 3929 3951
rect 3978 3948 3982 3951
rect 3994 3948 4054 3951
rect 4130 3948 4190 3951
rect 4194 3948 4230 3951
rect 4234 3948 4270 3951
rect 4410 3948 4414 3951
rect 4490 3948 4545 3951
rect 4554 3948 4558 3951
rect 4562 3948 4566 3951
rect 3470 3942 3473 3948
rect 3590 3942 3593 3948
rect 3622 3942 3625 3948
rect 2818 3938 2841 3941
rect 3126 3938 3206 3941
rect 3226 3938 3230 3941
rect 3378 3938 3430 3941
rect 3662 3938 3686 3941
rect 3746 3938 3782 3941
rect 3818 3938 3822 3941
rect 3858 3938 3926 3941
rect 3950 3941 3953 3948
rect 4366 3942 4369 3948
rect 4438 3942 4441 3948
rect 4470 3942 4473 3948
rect 3934 3938 3953 3941
rect 3970 3938 4046 3941
rect 4186 3938 4222 3941
rect 4226 3938 4230 3941
rect 4234 3938 4246 3941
rect 4250 3938 4302 3941
rect 4394 3938 4414 3941
rect 4542 3941 4545 3948
rect 4582 3941 4585 3948
rect 4630 3941 4634 3942
rect 4542 3938 4634 3941
rect 614 3932 617 3938
rect 3126 3932 3129 3938
rect 3662 3932 3665 3938
rect 3838 3932 3841 3938
rect 50 3928 78 3931
rect 82 3928 102 3931
rect 210 3928 326 3931
rect 378 3928 462 3931
rect 482 3928 598 3931
rect 730 3928 806 3931
rect 1306 3928 1694 3931
rect 1842 3928 1878 3931
rect 1890 3928 1950 3931
rect 1970 3928 1974 3931
rect 2082 3928 2086 3931
rect 2178 3928 2190 3931
rect 2378 3928 2382 3931
rect 2498 3928 2622 3931
rect 2666 3928 2718 3931
rect 2726 3928 2742 3931
rect 2746 3928 2758 3931
rect 2778 3928 2798 3931
rect 2834 3928 2854 3931
rect 3322 3928 3358 3931
rect 3362 3928 3526 3931
rect 3530 3928 3550 3931
rect 3554 3928 3590 3931
rect 3778 3928 3825 3931
rect 3882 3928 3894 3931
rect 3934 3931 3937 3938
rect 3922 3928 3937 3931
rect 3962 3928 3974 3931
rect 4194 3928 4238 3931
rect 4242 3928 4286 3931
rect 4290 3928 4294 3931
rect 4354 3928 4382 3931
rect 4394 3928 4502 3931
rect 4506 3928 4558 3931
rect 314 3918 326 3921
rect 338 3918 382 3921
rect 450 3918 454 3921
rect 598 3921 601 3928
rect 598 3918 630 3921
rect 754 3918 854 3921
rect 1186 3918 1510 3921
rect 1882 3918 2086 3921
rect 2374 3918 2382 3921
rect 2386 3918 2630 3921
rect 2634 3918 2670 3921
rect 2726 3921 2729 3928
rect 3822 3922 3825 3928
rect 2674 3918 2729 3921
rect 2738 3918 3198 3921
rect 3458 3918 3518 3921
rect 3522 3918 3630 3921
rect 3650 3918 3814 3921
rect 3834 3918 3934 3921
rect 4042 3918 4238 3921
rect 4298 3918 4302 3921
rect 4402 3918 4454 3921
rect 274 3908 414 3911
rect 490 3908 582 3911
rect 1226 3908 1310 3911
rect 1506 3908 1542 3911
rect 1738 3908 1766 3911
rect 1922 3908 1998 3911
rect 2234 3908 2270 3911
rect 2410 3908 2686 3911
rect 2706 3908 2718 3911
rect 2850 3908 2918 3911
rect 3586 3908 3710 3911
rect 3714 3908 3870 3911
rect 3914 3908 4070 3911
rect 4106 3908 4174 3911
rect 4218 3908 4518 3911
rect 4522 3908 4534 3911
rect 1000 3903 1002 3907
rect 1006 3903 1009 3907
rect 1014 3903 1016 3907
rect 2024 3903 2026 3907
rect 2030 3903 2033 3907
rect 2038 3903 2040 3907
rect 3048 3903 3050 3907
rect 3054 3903 3057 3907
rect 3062 3903 3064 3907
rect 4080 3903 4082 3907
rect 4086 3903 4089 3907
rect 4094 3903 4096 3907
rect 362 3898 510 3901
rect 514 3898 558 3901
rect 634 3898 774 3901
rect 778 3898 838 3901
rect 842 3898 854 3901
rect 1114 3898 1126 3901
rect 2154 3898 2302 3901
rect 2498 3898 2574 3901
rect 2586 3898 2710 3901
rect 2722 3898 2814 3901
rect 2826 3898 2886 3901
rect 2890 3898 2910 3901
rect 2914 3898 3006 3901
rect 3130 3898 3142 3901
rect 3394 3898 3582 3901
rect 3594 3898 3774 3901
rect 3802 3898 3974 3901
rect 3978 3898 4006 3901
rect 4226 3898 4350 3901
rect 574 3892 577 3898
rect 1502 3892 1505 3898
rect 466 3888 574 3891
rect 610 3888 694 3891
rect 714 3888 766 3891
rect 938 3888 942 3891
rect 1274 3888 1494 3891
rect 2018 3888 2406 3891
rect 2442 3888 2574 3891
rect 2578 3888 2606 3891
rect 2650 3888 2921 3891
rect 3010 3888 3030 3891
rect 3034 3888 3110 3891
rect 3818 3888 3878 3891
rect 4054 3888 4062 3891
rect 4066 3888 4102 3891
rect 4234 3888 4430 3891
rect 4434 3888 4441 3891
rect 4450 3888 4486 3891
rect 4490 3888 4550 3891
rect 98 3878 214 3881
rect 218 3878 422 3881
rect 562 3878 638 3881
rect 722 3878 726 3881
rect 730 3878 806 3881
rect 810 3878 926 3881
rect 1154 3878 1190 3881
rect 1314 3878 1526 3881
rect 1594 3878 1718 3881
rect 1866 3878 1953 3881
rect 2002 3878 2086 3881
rect 2090 3878 2118 3881
rect 2122 3878 2182 3881
rect 2386 3878 2390 3881
rect 2394 3878 2430 3881
rect 2490 3878 2494 3881
rect 2514 3878 2710 3881
rect 2730 3878 2902 3881
rect 2918 3881 2921 3888
rect 3142 3881 3145 3888
rect 2918 3878 3145 3881
rect 3258 3878 3430 3881
rect 3434 3878 3438 3881
rect 3442 3878 3494 3881
rect 3570 3878 3678 3881
rect 3762 3878 3782 3881
rect 3938 3878 3998 3881
rect 4002 3878 4038 3881
rect 4042 3878 4078 3881
rect 4274 3878 4310 3881
rect 4322 3878 4374 3881
rect 4426 3878 4534 3881
rect 334 3870 342 3871
rect 78 3861 81 3868
rect 338 3868 342 3870
rect 346 3868 366 3871
rect 546 3868 574 3871
rect 686 3871 689 3878
rect 578 3868 689 3871
rect 722 3868 910 3871
rect 914 3868 950 3871
rect 1070 3871 1073 3878
rect 986 3868 1073 3871
rect 1170 3868 1262 3871
rect 1266 3868 1286 3871
rect 1338 3868 1382 3871
rect 1498 3868 1622 3871
rect 1726 3871 1729 3878
rect 1726 3868 1910 3871
rect 1950 3871 1953 3878
rect 2246 3872 2249 3878
rect 1950 3868 2014 3871
rect 2034 3868 2086 3871
rect 2106 3868 2150 3871
rect 2178 3868 2214 3871
rect 2450 3868 2494 3871
rect 2506 3868 2702 3871
rect 2754 3868 2838 3871
rect 2874 3868 2878 3871
rect 2910 3871 2913 3878
rect 2910 3868 2942 3871
rect 3386 3868 3422 3871
rect 3498 3868 3566 3871
rect 3706 3870 3782 3871
rect 3706 3868 3742 3870
rect 78 3858 158 3861
rect 302 3858 350 3861
rect 354 3858 374 3861
rect 386 3858 630 3861
rect 770 3858 790 3861
rect 842 3858 846 3861
rect 1218 3858 1326 3861
rect 1474 3858 1566 3861
rect 1686 3858 1790 3861
rect 1938 3858 2046 3861
rect 2130 3858 2142 3861
rect 2178 3858 2278 3861
rect 2370 3858 2454 3861
rect 2466 3858 2598 3861
rect 2666 3858 2678 3861
rect 2706 3858 2718 3861
rect 2722 3858 2742 3861
rect 2850 3858 2894 3861
rect 2906 3858 2982 3861
rect 3022 3861 3025 3868
rect 3038 3861 3041 3868
rect 3022 3858 3041 3861
rect 3102 3861 3105 3868
rect 3118 3861 3121 3868
rect 3746 3868 3782 3870
rect 3846 3871 3849 3878
rect 3794 3868 3849 3871
rect 3918 3872 3921 3878
rect 3930 3868 3934 3871
rect 3954 3868 4022 3871
rect 4050 3868 4054 3871
rect 4146 3868 4206 3871
rect 4266 3868 4302 3871
rect 4306 3868 4326 3871
rect 4410 3868 4470 3871
rect 4474 3868 4481 3871
rect 4506 3868 4550 3871
rect 3102 3858 3121 3861
rect 3306 3858 3414 3861
rect 3418 3858 3462 3861
rect 3514 3858 3518 3861
rect 3594 3858 3694 3861
rect 3722 3858 3822 3861
rect 3890 3858 3918 3861
rect 3946 3858 3982 3861
rect 4066 3858 4158 3861
rect 4222 3861 4225 3868
rect 4222 3858 4262 3861
rect 4290 3858 4334 3861
rect 4354 3858 4366 3861
rect 4378 3858 4382 3861
rect 4402 3858 4430 3861
rect 4434 3858 4446 3861
rect 4530 3858 4558 3861
rect 302 3852 305 3858
rect -26 3851 -22 3852
rect -26 3848 6 3851
rect 666 3848 710 3851
rect 834 3848 854 3851
rect 902 3851 905 3858
rect 1406 3852 1409 3858
rect 1686 3852 1689 3858
rect 3294 3852 3297 3858
rect 902 3848 926 3851
rect 1182 3848 1198 3851
rect 1210 3848 1222 3851
rect 1778 3848 1854 3851
rect 1866 3848 1966 3851
rect 1994 3848 2054 3851
rect 2058 3848 2158 3851
rect 2162 3848 2214 3851
rect 2218 3848 2246 3851
rect 2374 3848 2414 3851
rect 2418 3848 2470 3851
rect 2474 3848 2502 3851
rect 2514 3848 2542 3851
rect 2562 3848 2566 3851
rect 2642 3848 2774 3851
rect 2858 3848 2870 3851
rect 2906 3848 3046 3851
rect 3074 3848 3078 3851
rect 3434 3848 3590 3851
rect 3682 3848 3758 3851
rect 3866 3848 3870 3851
rect 3874 3848 3886 3851
rect 4074 3848 4118 3851
rect 4218 3848 4230 3851
rect 4234 3848 4374 3851
rect 4458 3848 4526 3851
rect 4630 3851 4634 3852
rect 4554 3848 4634 3851
rect 218 3838 390 3841
rect 394 3838 510 3841
rect 814 3841 817 3848
rect 1182 3842 1185 3848
rect 2374 3842 2377 3848
rect 814 3838 870 3841
rect 1034 3838 1038 3841
rect 1042 3838 1110 3841
rect 1354 3838 1374 3841
rect 1378 3838 1422 3841
rect 1426 3838 1478 3841
rect 1754 3838 1830 3841
rect 1954 3838 1958 3841
rect 2002 3838 2006 3841
rect 2010 3838 2086 3841
rect 2090 3838 2118 3841
rect 2122 3838 2166 3841
rect 2234 3838 2238 3841
rect 2322 3838 2326 3841
rect 2426 3838 2470 3841
rect 2490 3838 2598 3841
rect 2606 3838 2678 3841
rect 2682 3838 2790 3841
rect 2794 3838 2830 3841
rect 2834 3838 2870 3841
rect 3018 3838 3062 3841
rect 3678 3841 3681 3848
rect 3354 3838 3681 3841
rect 3714 3838 3862 3841
rect 3866 3838 4030 3841
rect 4178 3838 4406 3841
rect 4442 3838 4462 3841
rect 1962 3828 1974 3831
rect 1986 3828 2278 3831
rect 2290 3828 2398 3831
rect 2402 3828 2518 3831
rect 2534 3828 2542 3831
rect 2606 3831 2609 3838
rect 2546 3828 2609 3831
rect 2618 3828 2646 3831
rect 2850 3828 3006 3831
rect 3010 3828 3086 3831
rect 3562 3828 3766 3831
rect 3770 3828 3806 3831
rect 3810 3828 3838 3831
rect 3986 3828 4134 3831
rect 4194 3828 4246 3831
rect 4274 3828 4438 3831
rect 970 3818 974 3821
rect 2114 3818 2230 3821
rect 2234 3818 2358 3821
rect 2378 3818 3382 3821
rect 3610 3818 4334 3821
rect 2130 3808 2150 3811
rect 2354 3808 2414 3811
rect 2418 3808 2486 3811
rect 2626 3808 2758 3811
rect 2802 3808 3174 3811
rect 3930 3808 4198 3811
rect 4202 3808 4230 3811
rect 4346 3808 4486 3811
rect 4490 3808 4598 3811
rect 496 3803 498 3807
rect 502 3803 505 3807
rect 510 3803 512 3807
rect 1520 3803 1522 3807
rect 1526 3803 1529 3807
rect 1534 3803 1536 3807
rect 1918 3802 1921 3808
rect 2544 3803 2546 3807
rect 2550 3803 2553 3807
rect 2558 3803 2560 3807
rect 3568 3803 3570 3807
rect 3574 3803 3577 3807
rect 3582 3803 3584 3807
rect 274 3798 430 3801
rect 434 3798 478 3801
rect 906 3798 1270 3801
rect 1282 3798 1438 3801
rect 2058 3798 2302 3801
rect 2314 3798 2534 3801
rect 2674 3798 2830 3801
rect 2858 3798 3006 3801
rect 4466 3798 4478 3801
rect 4546 3798 4582 3801
rect 238 3792 241 3798
rect 614 3792 617 3798
rect 322 3788 326 3791
rect 1106 3788 1134 3791
rect 1810 3788 1870 3791
rect 1874 3788 1926 3791
rect 2122 3788 2126 3791
rect 2162 3788 2366 3791
rect 2378 3788 2422 3791
rect 2426 3788 2702 3791
rect 2706 3788 2742 3791
rect 2746 3788 2766 3791
rect 2818 3788 2862 3791
rect 2882 3788 3278 3791
rect 3970 3788 4006 3791
rect 4010 3788 4054 3791
rect 4058 3788 4198 3791
rect 4202 3788 4206 3791
rect 1398 3782 1401 3788
rect 634 3778 678 3781
rect 1122 3778 1134 3781
rect 1386 3778 1398 3781
rect 1694 3781 1697 3788
rect 1482 3778 1697 3781
rect 2106 3778 2134 3781
rect 2374 3781 2377 3788
rect 2330 3778 2377 3781
rect 2714 3778 2862 3781
rect 2866 3778 3014 3781
rect 3234 3778 3606 3781
rect 3610 3778 3670 3781
rect 3674 3778 3790 3781
rect 3898 3778 3974 3781
rect 3854 3772 3857 3778
rect 506 3768 566 3771
rect 570 3768 1022 3771
rect 1298 3768 1326 3771
rect 1394 3768 1430 3771
rect 1442 3768 1502 3771
rect 1858 3768 1918 3771
rect 1970 3768 2158 3771
rect 2274 3768 2310 3771
rect 2346 3768 2350 3771
rect 2370 3768 2518 3771
rect 2538 3768 2598 3771
rect 2602 3768 2606 3771
rect 2762 3768 2806 3771
rect 2962 3768 3017 3771
rect 3026 3768 3414 3771
rect 3914 3768 3934 3771
rect 4138 3768 4254 3771
rect 4362 3768 4438 3771
rect 4630 3771 4634 3772
rect 4442 3768 4634 3771
rect 34 3758 174 3761
rect 650 3758 750 3761
rect 1290 3758 1358 3761
rect 1362 3758 1470 3761
rect 1490 3758 1558 3761
rect 1562 3758 1606 3761
rect 1690 3758 1878 3761
rect 1986 3758 2006 3761
rect 2074 3758 2126 3761
rect 2130 3758 2166 3761
rect 2258 3758 2278 3761
rect 2282 3758 2385 3761
rect 2530 3758 2534 3761
rect 2722 3758 2774 3761
rect 2810 3758 2886 3761
rect 2938 3758 2982 3761
rect 2986 3758 3006 3761
rect 3014 3761 3017 3768
rect 4294 3762 4297 3768
rect 3014 3758 3126 3761
rect 3270 3758 3278 3761
rect 3282 3758 3326 3761
rect 3346 3758 3398 3761
rect 3406 3758 3438 3761
rect 3842 3758 3926 3761
rect 4074 3758 4102 3761
rect 4322 3758 4326 3761
rect 4402 3758 4518 3761
rect -26 3751 -22 3752
rect -26 3748 6 3751
rect 18 3748 118 3751
rect 714 3748 726 3751
rect 790 3751 793 3758
rect 1062 3752 1065 3758
rect 2382 3752 2385 3758
rect 3406 3752 3409 3758
rect 762 3748 793 3751
rect 1146 3748 1214 3751
rect 1354 3748 1550 3751
rect 1674 3748 1750 3751
rect 34 3738 54 3741
rect 258 3738 366 3741
rect 370 3738 406 3741
rect 426 3738 558 3741
rect 562 3738 614 3741
rect 770 3738 774 3741
rect 934 3741 937 3748
rect 1770 3748 1902 3751
rect 1930 3748 1950 3751
rect 1954 3748 1990 3751
rect 2266 3748 2270 3751
rect 2274 3748 2310 3751
rect 2386 3748 2422 3751
rect 2514 3748 2534 3751
rect 2594 3748 2694 3751
rect 2722 3748 2846 3751
rect 3018 3748 3094 3751
rect 3122 3748 3142 3751
rect 3154 3748 3166 3751
rect 3170 3748 3198 3751
rect 3202 3748 3246 3751
rect 3250 3748 3262 3751
rect 3518 3751 3521 3758
rect 3458 3748 3521 3751
rect 3634 3748 3742 3751
rect 3806 3751 3809 3758
rect 4262 3752 4265 3758
rect 3746 3748 3809 3751
rect 3834 3748 3910 3751
rect 4026 3748 4046 3751
rect 4058 3748 4078 3751
rect 4274 3748 4310 3751
rect 4334 3751 4337 3758
rect 4314 3748 4337 3751
rect 4366 3751 4369 3758
rect 4354 3748 4369 3751
rect 4398 3751 4401 3758
rect 4386 3748 4422 3751
rect 4514 3748 4534 3751
rect 4630 3751 4634 3752
rect 4602 3748 4634 3751
rect 2054 3742 2057 3748
rect 874 3738 937 3741
rect 1170 3738 1190 3741
rect 1194 3738 1278 3741
rect 1282 3738 1382 3741
rect 1386 3738 1398 3741
rect 1402 3738 1406 3741
rect 1422 3738 1446 3741
rect 1578 3738 1678 3741
rect 1762 3738 1854 3741
rect 1858 3738 1878 3741
rect 1882 3738 1934 3741
rect 1938 3738 1982 3741
rect 2074 3738 2222 3741
rect 2226 3738 2398 3741
rect 2498 3738 2518 3741
rect 2538 3738 2542 3741
rect 2578 3738 2790 3741
rect 2878 3741 2881 3748
rect 2834 3738 2881 3741
rect 2934 3741 2937 3748
rect 2922 3738 2937 3741
rect 3002 3738 3014 3741
rect 3090 3738 3118 3741
rect 3274 3738 3406 3741
rect 3410 3738 3430 3741
rect 3434 3738 3462 3741
rect 3810 3738 3822 3741
rect 3954 3738 3982 3741
rect 3986 3738 4014 3741
rect 4090 3738 4198 3741
rect 4250 3738 4262 3741
rect 4266 3738 4302 3741
rect 4306 3738 4326 3741
rect 4362 3738 4390 3741
rect 4434 3738 4446 3741
rect 4490 3738 4502 3741
rect 1422 3732 1425 3738
rect 90 3728 102 3731
rect 106 3728 118 3731
rect 162 3728 446 3731
rect 450 3728 518 3731
rect 522 3728 553 3731
rect 770 3728 910 3731
rect 1314 3728 1366 3731
rect 1506 3728 1814 3731
rect 1858 3728 1894 3731
rect 2218 3728 2358 3731
rect 2666 3728 2822 3731
rect 2890 3728 2910 3731
rect 2946 3728 3038 3731
rect 3130 3728 3254 3731
rect 3362 3728 3534 3731
rect 3778 3728 3798 3731
rect 3802 3728 3822 3731
rect 3842 3728 3878 3731
rect 3894 3731 3897 3738
rect 3882 3728 3958 3731
rect 3962 3728 3998 3731
rect 4002 3728 4038 3731
rect 4290 3728 4398 3731
rect 4402 3728 4438 3731
rect 4458 3728 4470 3731
rect 4474 3728 4542 3731
rect 4546 3728 4550 3731
rect 4554 3728 4566 3731
rect 550 3722 553 3728
rect 126 3718 134 3721
rect 138 3718 270 3721
rect 554 3718 662 3721
rect 706 3718 734 3721
rect 1026 3718 1198 3721
rect 1218 3718 1262 3721
rect 1298 3718 1478 3721
rect 1830 3721 1833 3728
rect 1830 3718 2318 3721
rect 2322 3718 2334 3721
rect 2446 3721 2449 3728
rect 2798 3722 2801 3728
rect 2446 3718 2793 3721
rect 2926 3721 2929 3728
rect 2926 3718 2998 3721
rect 3226 3718 3438 3721
rect 3738 3718 3782 3721
rect 3786 3718 3798 3721
rect 3814 3718 3886 3721
rect 3890 3718 4310 3721
rect 4402 3718 4414 3721
rect 4418 3718 4462 3721
rect 4466 3718 4534 3721
rect 4538 3718 4566 3721
rect 4570 3718 4582 3721
rect 2342 3712 2345 3718
rect 1026 3708 1158 3711
rect 1234 3708 1838 3711
rect 1850 3708 1934 3711
rect 2146 3708 2238 3711
rect 2290 3708 2334 3711
rect 2354 3708 2606 3711
rect 2738 3708 2742 3711
rect 2790 3711 2793 3718
rect 3814 3712 3817 3718
rect 2790 3708 2862 3711
rect 2906 3708 2926 3711
rect 3114 3708 3262 3711
rect 3394 3708 3398 3711
rect 3714 3708 3758 3711
rect 3762 3708 3782 3711
rect 4114 3708 4126 3711
rect 4130 3708 4158 3711
rect 1000 3703 1002 3707
rect 1006 3703 1009 3707
rect 1014 3703 1016 3707
rect 2024 3703 2026 3707
rect 2030 3703 2033 3707
rect 2038 3703 2040 3707
rect 3048 3703 3050 3707
rect 3054 3703 3057 3707
rect 3062 3703 3064 3707
rect 4080 3703 4082 3707
rect 4086 3703 4089 3707
rect 4094 3703 4096 3707
rect 1162 3698 1454 3701
rect 1522 3698 1726 3701
rect 1730 3698 1798 3701
rect 1810 3698 1934 3701
rect 1962 3698 1990 3701
rect 2090 3698 2182 3701
rect 2186 3698 2262 3701
rect 2274 3698 2566 3701
rect 2574 3698 2806 3701
rect 2874 3698 2942 3701
rect 3098 3698 3238 3701
rect 4122 3698 4478 3701
rect 1110 3692 1113 3698
rect 362 3688 590 3691
rect 594 3688 670 3691
rect 810 3688 814 3691
rect 990 3688 1038 3691
rect 1178 3688 1182 3691
rect 1306 3688 1750 3691
rect 1842 3688 2022 3691
rect 2574 3691 2577 3698
rect 3494 3692 3497 3698
rect 2458 3688 2577 3691
rect 2626 3688 2694 3691
rect 2722 3688 2726 3691
rect 2746 3688 2902 3691
rect 3018 3688 3169 3691
rect 3178 3688 3486 3691
rect 3962 3688 4190 3691
rect 4258 3688 4326 3691
rect 4330 3688 4382 3691
rect 38 3681 41 3688
rect 990 3682 993 3688
rect 2326 3682 2329 3688
rect 38 3678 86 3681
rect 90 3678 134 3681
rect 170 3678 262 3681
rect 266 3678 502 3681
rect 1146 3678 1286 3681
rect 1450 3678 1886 3681
rect 1938 3678 2078 3681
rect 2138 3678 2150 3681
rect 2266 3678 2294 3681
rect 2342 3681 2345 3688
rect 2342 3678 2374 3681
rect 2394 3678 2462 3681
rect 2690 3678 2718 3681
rect 2770 3678 2806 3681
rect 2810 3678 2854 3681
rect 2890 3678 2894 3681
rect 2898 3678 2966 3681
rect 3066 3678 3102 3681
rect 3166 3681 3169 3688
rect 3166 3678 3206 3681
rect 3434 3678 3734 3681
rect 4002 3678 4113 3681
rect 4122 3678 4134 3681
rect 4138 3678 4166 3681
rect -26 3671 -22 3672
rect -26 3668 6 3671
rect 114 3668 134 3671
rect 226 3668 286 3671
rect 290 3668 345 3671
rect 326 3662 329 3668
rect 342 3662 345 3668
rect 630 3668 662 3671
rect 870 3671 873 3678
rect 2150 3672 2153 3678
rect 870 3668 910 3671
rect 930 3668 1046 3671
rect 1050 3668 1206 3671
rect 1246 3668 1350 3671
rect 1442 3668 1470 3671
rect 1746 3668 1798 3671
rect 2202 3668 2310 3671
rect 2314 3668 2425 3671
rect 2434 3668 2494 3671
rect 2590 3671 2593 3678
rect 2546 3668 2593 3671
rect 2630 3668 2654 3671
rect 2682 3668 2734 3671
rect 2762 3668 2774 3671
rect 2834 3668 2846 3671
rect 2914 3668 2934 3671
rect 2994 3668 3102 3671
rect 3114 3668 3118 3671
rect 3186 3668 3190 3671
rect 3210 3668 3214 3671
rect 3226 3668 3230 3671
rect 3450 3668 3630 3671
rect 3666 3668 3814 3671
rect 3930 3668 4030 3671
rect 4034 3668 4102 3671
rect 4110 3671 4113 3678
rect 4142 3672 4145 3678
rect 4110 3668 4126 3671
rect 4146 3668 4174 3671
rect 4178 3668 4222 3671
rect 4262 3671 4265 3678
rect 4226 3668 4265 3671
rect 4466 3668 4510 3671
rect 4514 3668 4566 3671
rect 382 3662 385 3668
rect 542 3662 545 3668
rect 630 3662 633 3668
rect 1246 3662 1249 3668
rect 58 3658 94 3661
rect 98 3658 126 3661
rect 730 3658 910 3661
rect 914 3658 918 3661
rect 986 3658 1030 3661
rect 1726 3661 1729 3668
rect 2134 3662 2137 3668
rect 1726 3658 1846 3661
rect 1890 3658 1918 3661
rect 1922 3658 1958 3661
rect 1970 3658 1982 3661
rect 2146 3658 2198 3661
rect 2226 3658 2270 3661
rect 2274 3658 2390 3661
rect 2394 3658 2406 3661
rect 2422 3661 2425 3668
rect 2422 3658 2438 3661
rect 2442 3658 2454 3661
rect 2582 3658 2590 3661
rect 2630 3661 2633 3668
rect 2750 3662 2753 3668
rect 2950 3662 2953 3668
rect 2594 3658 2633 3661
rect 2642 3658 2662 3661
rect 2706 3658 2710 3661
rect 2730 3658 2742 3661
rect 2802 3658 2846 3661
rect 3082 3658 3118 3661
rect 3134 3661 3137 3668
rect 3134 3658 3150 3661
rect 3170 3658 3222 3661
rect 3314 3658 3342 3661
rect 3346 3658 3414 3661
rect 3546 3658 3550 3661
rect 3730 3658 3742 3661
rect 3914 3658 4022 3661
rect 4026 3658 4030 3661
rect 4042 3658 4094 3661
rect 4122 3658 4150 3661
rect 4154 3658 4182 3661
rect 4186 3658 4214 3661
rect 4266 3658 4278 3661
rect 4282 3658 4406 3661
rect 1054 3652 1057 3658
rect 1590 3652 1593 3658
rect -26 3651 -22 3652
rect -26 3648 70 3651
rect 114 3648 190 3651
rect 626 3648 798 3651
rect 802 3648 838 3651
rect 1130 3648 1150 3651
rect 1826 3648 1942 3651
rect 1986 3648 1990 3651
rect 2026 3648 2270 3651
rect 2278 3648 2286 3651
rect 2290 3648 2302 3651
rect 2330 3648 2350 3651
rect 2470 3651 2473 3658
rect 2870 3652 2873 3658
rect 2354 3648 2473 3651
rect 2482 3648 2518 3651
rect 2554 3648 2558 3651
rect 2602 3648 2630 3651
rect 2634 3648 2774 3651
rect 2814 3648 2862 3651
rect 2946 3648 3014 3651
rect 3042 3648 3086 3651
rect 3106 3648 3150 3651
rect 3182 3648 3294 3651
rect 3410 3648 3438 3651
rect 4026 3648 4033 3651
rect 4058 3648 4070 3651
rect 4082 3648 4150 3651
rect 4186 3648 4190 3651
rect 4314 3648 4526 3651
rect 4530 3648 4542 3651
rect 778 3638 782 3641
rect 1378 3638 1790 3641
rect 1794 3638 1862 3641
rect 2006 3641 2009 3648
rect 2574 3642 2577 3648
rect 2814 3642 2817 3648
rect 3182 3642 3185 3648
rect 4030 3642 4033 3648
rect 1954 3638 2014 3641
rect 2170 3638 2206 3641
rect 2234 3638 2262 3641
rect 2266 3638 2334 3641
rect 2338 3638 2382 3641
rect 2386 3638 2406 3641
rect 2482 3638 2526 3641
rect 2650 3638 2702 3641
rect 2706 3638 2737 3641
rect 2746 3638 2790 3641
rect 2834 3638 2838 3641
rect 2970 3638 3054 3641
rect 3074 3638 3118 3641
rect 3218 3638 3366 3641
rect 4322 3638 4326 3641
rect 4338 3638 4374 3641
rect 4378 3638 4478 3641
rect 4502 3638 4518 3641
rect 2734 3632 2737 3638
rect 4502 3632 4505 3638
rect 618 3628 774 3631
rect 778 3628 862 3631
rect 1890 3628 2102 3631
rect 2130 3628 2286 3631
rect 2370 3628 2430 3631
rect 2474 3628 2518 3631
rect 2522 3628 2590 3631
rect 2610 3628 2686 3631
rect 2738 3628 2822 3631
rect 3082 3628 3174 3631
rect 3258 3628 3281 3631
rect 3890 3628 3990 3631
rect 3994 3628 4214 3631
rect 1442 3618 1654 3621
rect 2138 3618 2142 3621
rect 2190 3618 2198 3621
rect 2202 3618 2262 3621
rect 2278 3618 2726 3621
rect 2830 3618 2838 3621
rect 2842 3618 2990 3621
rect 3014 3621 3017 3628
rect 3278 3622 3281 3628
rect 3014 3618 3214 3621
rect 3226 3618 3270 3621
rect 3274 3618 3278 3621
rect 3694 3618 4022 3621
rect 4234 3618 4366 3621
rect 4370 3618 4374 3621
rect 4378 3618 4446 3621
rect 4450 3618 4574 3621
rect 2278 3611 2281 3618
rect 2114 3608 2281 3611
rect 2290 3608 2470 3611
rect 2726 3611 2729 3618
rect 3694 3612 3697 3618
rect 2726 3608 3022 3611
rect 3250 3608 3438 3611
rect 3594 3608 3694 3611
rect 496 3603 498 3607
rect 502 3603 505 3607
rect 510 3603 512 3607
rect 1520 3603 1522 3607
rect 1526 3603 1529 3607
rect 1534 3603 1536 3607
rect 2494 3602 2497 3608
rect 2544 3603 2546 3607
rect 2550 3603 2553 3607
rect 2558 3603 2560 3607
rect 3568 3603 3570 3607
rect 3574 3603 3577 3607
rect 3582 3603 3584 3607
rect 1802 3598 2089 3601
rect 2098 3598 2438 3601
rect 2506 3598 2518 3601
rect 2594 3598 2694 3601
rect 2994 3598 3238 3601
rect 3410 3598 3462 3601
rect 3594 3598 3774 3601
rect 3778 3598 4270 3601
rect 1250 3588 1414 3591
rect 2018 3588 2070 3591
rect 2086 3591 2089 3598
rect 2086 3588 2190 3591
rect 2218 3588 2310 3591
rect 2434 3588 2465 3591
rect 2490 3588 2662 3591
rect 2770 3588 3030 3591
rect 3106 3588 3326 3591
rect 3406 3588 3510 3591
rect 3546 3588 3726 3591
rect 3730 3588 3902 3591
rect 4226 3588 4462 3591
rect 410 3578 494 3581
rect 1918 3581 1921 3588
rect 2462 3582 2465 3588
rect 3406 3582 3409 3588
rect 1918 3578 2446 3581
rect 2490 3578 2537 3581
rect 2842 3578 2862 3581
rect 2866 3578 2950 3581
rect 2954 3578 2974 3581
rect 2986 3578 2998 3581
rect 3114 3578 3190 3581
rect 3338 3578 3358 3581
rect 3474 3578 3614 3581
rect 3618 3578 4014 3581
rect 4330 3578 4534 3581
rect 4538 3578 4566 3581
rect 2534 3572 2537 3578
rect 202 3568 374 3571
rect 378 3568 486 3571
rect 490 3568 558 3571
rect 746 3568 766 3571
rect 1650 3568 1742 3571
rect 2458 3568 2462 3571
rect 2490 3568 2494 3571
rect 2506 3568 2510 3571
rect 2634 3568 2646 3571
rect 2662 3568 2710 3571
rect 2778 3568 2782 3571
rect 2858 3568 2886 3571
rect 2890 3568 2990 3571
rect 2994 3568 3006 3571
rect 3098 3568 3150 3571
rect 3154 3568 3230 3571
rect 3234 3568 3286 3571
rect 3290 3568 3310 3571
rect 3330 3568 3334 3571
rect 3394 3568 3726 3571
rect 3738 3568 3798 3571
rect 3818 3568 3878 3571
rect 3890 3568 4422 3571
rect 4426 3568 4430 3571
rect 290 3558 318 3561
rect 322 3558 446 3561
rect 466 3558 526 3561
rect 746 3558 798 3561
rect 1146 3558 1174 3561
rect 1394 3558 1918 3561
rect 1966 3558 2022 3561
rect 2142 3561 2145 3568
rect 2138 3558 2145 3561
rect 2162 3558 2166 3561
rect 2178 3558 2390 3561
rect 2662 3561 2665 3568
rect 2450 3558 2665 3561
rect 2722 3558 2806 3561
rect 2810 3558 3006 3561
rect 3082 3558 3374 3561
rect 3386 3558 3398 3561
rect 3426 3558 3430 3561
rect 3746 3558 3886 3561
rect 3906 3558 3982 3561
rect 3986 3558 4342 3561
rect 4346 3558 4518 3561
rect 4522 3558 4590 3561
rect -26 3551 -22 3552
rect -26 3548 6 3551
rect 126 3551 129 3558
rect 790 3552 793 3558
rect 66 3548 129 3551
rect 402 3548 414 3551
rect 418 3548 454 3551
rect 762 3548 782 3551
rect 890 3548 1078 3551
rect 1082 3548 1086 3551
rect 566 3542 569 3548
rect 26 3538 70 3541
rect 418 3538 438 3541
rect 630 3541 633 3548
rect 646 3541 649 3548
rect 1258 3548 1390 3551
rect 1394 3548 1398 3551
rect 1446 3548 1494 3551
rect 1446 3542 1449 3548
rect 1514 3548 1518 3551
rect 1538 3548 1574 3551
rect 1578 3548 1622 3551
rect 1626 3548 1785 3551
rect 1686 3542 1689 3548
rect 1782 3542 1785 3548
rect 1966 3551 1969 3558
rect 2670 3552 2673 3558
rect 1866 3548 1969 3551
rect 1978 3548 1982 3551
rect 2066 3548 2102 3551
rect 1814 3542 1817 3548
rect 2378 3548 2638 3551
rect 2770 3548 2782 3551
rect 2842 3548 2846 3551
rect 2850 3548 2886 3551
rect 2890 3548 2982 3551
rect 3018 3548 3110 3551
rect 3542 3551 3545 3558
rect 3490 3548 3545 3551
rect 3742 3552 3745 3558
rect 3754 3548 3926 3551
rect 2654 3542 2657 3548
rect 578 3538 649 3541
rect 978 3538 990 3541
rect 1034 3538 1161 3541
rect 1354 3538 1382 3541
rect 1890 3538 1918 3541
rect 1922 3538 1982 3541
rect 1986 3538 2038 3541
rect 2042 3538 2054 3541
rect 2058 3538 2094 3541
rect 2146 3538 2166 3541
rect 2306 3538 2310 3541
rect 2322 3538 2326 3541
rect 2418 3538 2422 3541
rect 2434 3538 2446 3541
rect 2530 3538 2542 3541
rect 2562 3538 2606 3541
rect 2682 3538 2894 3541
rect 2922 3538 2966 3541
rect 3126 3541 3129 3548
rect 4242 3548 4318 3551
rect 3126 3538 3150 3541
rect 3186 3538 3278 3541
rect 3298 3538 3342 3541
rect 3402 3538 3414 3541
rect 3418 3538 3494 3541
rect 3578 3538 3686 3541
rect 3690 3538 3806 3541
rect 3998 3541 4001 3548
rect 4110 3541 4113 3548
rect 3954 3538 4206 3541
rect 4218 3538 4222 3541
rect 4350 3541 4353 3548
rect 4226 3538 4353 3541
rect 4498 3538 4510 3541
rect 1062 3532 1065 3538
rect 1158 3532 1161 3538
rect 2478 3532 2481 3538
rect -26 3531 -22 3532
rect -26 3528 30 3531
rect 130 3528 230 3531
rect 322 3528 670 3531
rect 1274 3528 1422 3531
rect 1426 3528 1446 3531
rect 1722 3528 1862 3531
rect 1978 3528 1998 3531
rect 2010 3528 2038 3531
rect 2170 3528 2238 3531
rect 2282 3528 2382 3531
rect 2418 3528 2422 3531
rect 2490 3528 2686 3531
rect 2690 3528 3046 3531
rect 3058 3528 3086 3531
rect 3090 3528 3358 3531
rect 3510 3531 3513 3538
rect 3510 3528 3654 3531
rect 4334 3528 4494 3531
rect 90 3518 190 3521
rect 1210 3518 1846 3521
rect 1954 3518 2014 3521
rect 2018 3518 2190 3521
rect 2194 3518 2270 3521
rect 2394 3518 2478 3521
rect 2522 3518 2710 3521
rect 2714 3518 2806 3521
rect 2810 3518 2870 3521
rect 2874 3518 2942 3521
rect 2946 3518 2966 3521
rect 3066 3518 3094 3521
rect 3226 3518 3254 3521
rect 3314 3518 3318 3521
rect 3338 3518 3342 3521
rect 3862 3521 3865 3528
rect 4334 3522 4337 3528
rect 3862 3518 3886 3521
rect 726 3512 729 3518
rect 3462 3512 3465 3518
rect 1626 3508 1654 3511
rect 1946 3508 1982 3511
rect 2250 3508 2350 3511
rect 2826 3508 2862 3511
rect 4186 3508 4230 3511
rect 4234 3508 4254 3511
rect 4258 3508 4406 3511
rect 1000 3503 1002 3507
rect 1006 3503 1009 3507
rect 1014 3503 1016 3507
rect 2024 3503 2026 3507
rect 2030 3503 2033 3507
rect 2038 3503 2040 3507
rect 2414 3502 2417 3508
rect 2654 3502 2657 3508
rect 2918 3502 2921 3508
rect 3048 3503 3050 3507
rect 3054 3503 3057 3507
rect 3062 3503 3064 3507
rect 4080 3503 4082 3507
rect 4086 3503 4089 3507
rect 4094 3503 4096 3507
rect 1954 3498 2006 3501
rect 2250 3498 2366 3501
rect 2678 3498 2782 3501
rect 2930 3498 3014 3501
rect 3154 3498 3294 3501
rect 3522 3498 4070 3501
rect 4106 3498 4246 3501
rect 4250 3498 4294 3501
rect 378 3488 529 3491
rect 538 3488 606 3491
rect 754 3488 806 3491
rect 1026 3488 1030 3491
rect 1146 3488 1246 3491
rect 1418 3488 1502 3491
rect 1786 3488 1790 3491
rect 1922 3488 1942 3491
rect 1970 3488 2134 3491
rect 2234 3488 2262 3491
rect 2266 3488 2422 3491
rect 2678 3491 2681 3498
rect 2582 3488 2681 3491
rect 2690 3488 2694 3491
rect 2914 3488 3222 3491
rect 3506 3488 3726 3491
rect 3730 3488 4126 3491
rect 82 3478 142 3481
rect 230 3481 233 3488
rect 146 3478 310 3481
rect 314 3478 374 3481
rect 426 3478 446 3481
rect 474 3478 478 3481
rect 526 3481 529 3488
rect 526 3478 558 3481
rect 750 3481 753 3488
rect 666 3478 753 3481
rect 830 3482 833 3488
rect 2582 3482 2585 3488
rect 1346 3478 1438 3481
rect 1770 3478 1902 3481
rect 1938 3478 1998 3481
rect 2002 3478 2094 3481
rect 2098 3478 2142 3481
rect 2194 3478 2198 3481
rect 2218 3478 2350 3481
rect 2370 3478 2438 3481
rect 2506 3478 2566 3481
rect 2666 3478 2830 3481
rect 2834 3478 2894 3481
rect 2914 3478 3518 3481
rect 3626 3478 3742 3481
rect 3794 3478 3862 3481
rect 3866 3478 4110 3481
rect 4322 3478 4366 3481
rect 4370 3478 4382 3481
rect 34 3468 54 3471
rect 82 3468 94 3471
rect 98 3468 118 3471
rect 122 3468 286 3471
rect 394 3468 438 3471
rect 738 3468 750 3471
rect 942 3471 945 3478
rect 898 3468 945 3471
rect 1482 3468 1638 3471
rect 1906 3468 1942 3471
rect 1962 3468 1990 3471
rect 2026 3468 2030 3471
rect 2050 3468 2142 3471
rect 2146 3468 2174 3471
rect 2266 3468 2302 3471
rect 2434 3468 2454 3471
rect 2490 3468 2526 3471
rect 2530 3468 2622 3471
rect 2690 3468 2726 3471
rect 2874 3468 2878 3471
rect 2938 3468 2942 3471
rect 3010 3468 3022 3471
rect 3042 3468 3102 3471
rect 3218 3468 3254 3471
rect 3290 3468 3318 3471
rect 3362 3468 3390 3471
rect 3394 3468 3414 3471
rect 3434 3468 3470 3471
rect 3498 3468 3510 3471
rect 3514 3468 3574 3471
rect 3834 3468 4006 3471
rect 4010 3468 4222 3471
rect 4282 3468 4350 3471
rect 4362 3468 4430 3471
rect 4434 3468 4454 3471
rect 50 3458 126 3461
rect 226 3458 230 3461
rect 290 3458 302 3461
rect 306 3458 366 3461
rect 510 3461 513 3468
rect 510 3458 662 3461
rect 1310 3461 1313 3468
rect 1202 3458 1313 3461
rect 1362 3458 1398 3461
rect 1402 3458 1494 3461
rect 1574 3458 1974 3461
rect 2010 3458 2070 3461
rect 2074 3458 2094 3461
rect 2146 3458 2294 3461
rect 2374 3461 2377 3468
rect 2346 3458 2377 3461
rect 2530 3458 2598 3461
rect 2646 3461 2649 3468
rect 2634 3458 2649 3461
rect 2666 3458 2694 3461
rect 2822 3461 2825 3468
rect 2838 3461 2841 3468
rect 2822 3458 2841 3461
rect 2902 3461 2905 3468
rect 3142 3462 3145 3468
rect 2874 3458 2905 3461
rect 2914 3458 2926 3461
rect 2970 3458 2990 3461
rect 2994 3458 3030 3461
rect 3082 3458 3086 3461
rect 3106 3458 3126 3461
rect 3162 3458 3166 3461
rect 3218 3458 3278 3461
rect 3346 3458 3350 3461
rect 3370 3458 3374 3461
rect 3466 3458 3478 3461
rect 3654 3461 3657 3468
rect 3610 3458 3657 3461
rect 3746 3458 3766 3461
rect 3786 3458 3846 3461
rect 3866 3458 3886 3461
rect 3946 3459 3950 3461
rect 3946 3458 3953 3459
rect 4034 3458 4254 3461
rect 4258 3458 4294 3461
rect 4330 3458 4390 3461
rect 4518 3461 4521 3468
rect 4506 3458 4521 3461
rect 254 3452 257 3458
rect 1574 3452 1577 3458
rect -26 3451 -22 3452
rect -26 3448 6 3451
rect 178 3448 254 3451
rect 450 3448 462 3451
rect 466 3448 470 3451
rect 498 3448 518 3451
rect 930 3448 958 3451
rect 1258 3448 1382 3451
rect 1442 3448 1454 3451
rect 1674 3448 2086 3451
rect 2094 3448 2102 3451
rect 2106 3448 2158 3451
rect 2190 3448 2206 3451
rect 2234 3448 2254 3451
rect 2286 3448 2294 3451
rect 2298 3448 2318 3451
rect 2446 3451 2449 3458
rect 2798 3452 2801 3458
rect 2446 3448 2478 3451
rect 2626 3448 2670 3451
rect 2674 3448 2734 3451
rect 2738 3448 2782 3451
rect 2818 3448 2846 3451
rect 2858 3448 2886 3451
rect 2898 3448 2918 3451
rect 2938 3448 2942 3451
rect 3094 3451 3097 3458
rect 3018 3448 3118 3451
rect 3122 3448 3150 3451
rect 3178 3448 3198 3451
rect 3226 3448 3278 3451
rect 3282 3448 3326 3451
rect 3466 3448 3609 3451
rect 3618 3448 3726 3451
rect 3754 3448 3782 3451
rect 3886 3448 4038 3451
rect 4106 3448 4310 3451
rect 4362 3448 4374 3451
rect 4542 3451 4545 3458
rect 4434 3448 4545 3451
rect 2190 3442 2193 3448
rect 458 3438 502 3441
rect 730 3438 1590 3441
rect 1930 3438 1950 3441
rect 1954 3438 1958 3441
rect 2242 3438 2334 3441
rect 2382 3441 2385 3448
rect 2382 3438 2390 3441
rect 2474 3438 2486 3441
rect 2522 3438 2574 3441
rect 2578 3438 2614 3441
rect 2626 3438 2654 3441
rect 2690 3438 2694 3441
rect 2730 3438 2806 3441
rect 2810 3438 2838 3441
rect 2882 3438 2958 3441
rect 2998 3441 3001 3448
rect 3606 3442 3609 3448
rect 3886 3442 3889 3448
rect 2978 3438 3022 3441
rect 3154 3438 3198 3441
rect 3314 3438 3350 3441
rect 3530 3438 3598 3441
rect 4194 3438 4382 3441
rect 4394 3438 4502 3441
rect 4506 3438 4510 3441
rect 4550 3441 4553 3448
rect 4526 3438 4553 3441
rect 4526 3432 4529 3438
rect 826 3428 870 3431
rect 874 3428 1230 3431
rect 1938 3428 2198 3431
rect 2242 3428 2366 3431
rect 2418 3428 2430 3431
rect 2434 3428 2670 3431
rect 2938 3428 2966 3431
rect 3002 3428 3014 3431
rect 3234 3428 3430 3431
rect 3602 3428 3990 3431
rect 3994 3428 4222 3431
rect 786 3418 822 3421
rect 1154 3418 1198 3421
rect 1562 3418 1598 3421
rect 2206 3421 2209 3428
rect 2206 3418 2494 3421
rect 2506 3418 2862 3421
rect 2886 3421 2889 3428
rect 2886 3418 2990 3421
rect 1610 3408 1702 3411
rect 1810 3408 1910 3411
rect 2682 3408 2686 3411
rect 2762 3408 2974 3411
rect 3042 3408 3310 3411
rect 3322 3408 3534 3411
rect 496 3403 498 3407
rect 502 3403 505 3407
rect 510 3403 512 3407
rect 1520 3403 1522 3407
rect 1526 3403 1529 3407
rect 1534 3403 1536 3407
rect 2544 3403 2546 3407
rect 2550 3403 2553 3407
rect 2558 3403 2560 3407
rect 3568 3403 3570 3407
rect 3574 3403 3577 3407
rect 3582 3403 3584 3407
rect 1866 3398 2214 3401
rect 2306 3398 2510 3401
rect 2738 3398 2822 3401
rect 2834 3398 2886 3401
rect 3138 3398 3398 3401
rect 1042 3388 1070 3391
rect 1106 3388 1246 3391
rect 1450 3388 1550 3391
rect 2122 3388 2254 3391
rect 2282 3388 2334 3391
rect 2402 3388 2430 3391
rect 2530 3388 2550 3391
rect 2610 3388 2646 3391
rect 2674 3388 2678 3391
rect 2786 3388 2822 3391
rect 2842 3388 2846 3391
rect 3098 3388 3190 3391
rect 3410 3388 3462 3391
rect 4106 3388 4110 3391
rect 4178 3388 4566 3391
rect 434 3378 558 3381
rect 586 3378 694 3381
rect 1210 3378 1270 3381
rect 2118 3378 2150 3381
rect 2450 3378 2630 3381
rect 2658 3378 2734 3381
rect 2754 3378 2846 3381
rect 2898 3378 2926 3381
rect 2962 3378 2998 3381
rect 3114 3378 3118 3381
rect 3154 3378 3166 3381
rect 3194 3378 3470 3381
rect 3482 3378 3502 3381
rect 3618 3378 3638 3381
rect 3734 3381 3737 3388
rect 3734 3378 3886 3381
rect 4322 3378 4486 3381
rect 4490 3378 4494 3381
rect 34 3368 206 3371
rect 546 3368 654 3371
rect 1910 3371 1913 3378
rect 2118 3372 2121 3378
rect 1698 3368 1913 3371
rect 1922 3368 1961 3371
rect 2250 3368 2254 3371
rect 2322 3368 2366 3371
rect 2418 3368 2438 3371
rect 2522 3368 2526 3371
rect 2570 3368 2606 3371
rect 2618 3368 2742 3371
rect 2778 3368 2782 3371
rect 2818 3368 2830 3371
rect 2914 3368 3361 3371
rect 3370 3368 3745 3371
rect 3850 3368 4126 3371
rect 34 3358 110 3361
rect 142 3358 366 3361
rect 570 3358 726 3361
rect 1222 3361 1225 3368
rect 1958 3362 1961 3368
rect 1222 3358 1326 3361
rect 1546 3358 1630 3361
rect 1666 3358 1798 3361
rect 1994 3358 2102 3361
rect 2114 3358 2134 3361
rect 2142 3361 2145 3368
rect 2262 3362 2265 3368
rect 3358 3362 3361 3368
rect 3742 3362 3745 3368
rect 2142 3358 2166 3361
rect 2178 3358 2230 3361
rect 2314 3358 2438 3361
rect 2442 3358 2486 3361
rect 2490 3358 2582 3361
rect 2786 3358 2934 3361
rect 2962 3358 2966 3361
rect 3002 3358 3006 3361
rect 3074 3358 3134 3361
rect 3154 3358 3158 3361
rect 3170 3358 3174 3361
rect 3202 3358 3241 3361
rect 3282 3358 3294 3361
rect 3378 3358 3462 3361
rect 3482 3358 3670 3361
rect 4334 3361 4337 3368
rect 4314 3358 4337 3361
rect 4514 3358 4542 3361
rect 142 3352 145 3358
rect -26 3351 -22 3352
rect -26 3348 6 3351
rect 58 3348 142 3351
rect 162 3348 302 3351
rect 306 3348 470 3351
rect 642 3348 678 3351
rect 794 3348 1134 3351
rect 1138 3348 1142 3351
rect 1194 3348 1270 3351
rect 1414 3351 1417 3358
rect 3238 3352 3241 3358
rect 1298 3348 1417 3351
rect 1582 3348 1590 3351
rect 1594 3348 1670 3351
rect 1478 3342 1481 3348
rect 1762 3348 1766 3351
rect 1786 3348 1849 3351
rect 1954 3348 2094 3351
rect 2098 3348 2110 3351
rect 2202 3348 2238 3351
rect 2242 3348 2286 3351
rect 2298 3348 2302 3351
rect 2306 3348 2334 3351
rect 2338 3348 2374 3351
rect 2482 3348 2598 3351
rect 2610 3348 2734 3351
rect 2826 3348 2846 3351
rect 2906 3348 2918 3351
rect 2994 3348 2998 3351
rect 3090 3348 3110 3351
rect 3282 3348 3366 3351
rect 3378 3348 3398 3351
rect 3402 3348 3430 3351
rect 3450 3348 3526 3351
rect 3538 3348 3550 3351
rect 3650 3348 3686 3351
rect 3690 3348 3726 3351
rect 3786 3348 3830 3351
rect 3890 3348 3921 3351
rect 4282 3348 4326 3351
rect 4330 3348 4358 3351
rect 4454 3351 4457 3358
rect 4454 3348 4518 3351
rect 4522 3348 4558 3351
rect 1846 3342 1849 3348
rect 34 3338 54 3341
rect 346 3338 366 3341
rect 530 3338 590 3341
rect 594 3338 630 3341
rect 890 3338 926 3341
rect 930 3338 934 3341
rect 946 3338 1017 3341
rect 1066 3338 1113 3341
rect 1562 3338 1598 3341
rect 1666 3338 1686 3341
rect 1962 3338 2094 3341
rect 2098 3338 2102 3341
rect 2106 3338 2118 3341
rect 2182 3341 2185 3348
rect 2122 3338 2185 3341
rect 2194 3338 2342 3341
rect 2390 3341 2393 3348
rect 2346 3338 2393 3341
rect 2410 3338 2446 3341
rect 2690 3338 2790 3341
rect 2806 3341 2809 3348
rect 2806 3338 2854 3341
rect 2882 3338 2913 3341
rect 2922 3338 2961 3341
rect 2970 3338 2974 3341
rect 3262 3341 3265 3348
rect 3918 3342 3921 3348
rect 3258 3338 3265 3341
rect 3290 3338 3310 3341
rect 3322 3338 3342 3341
rect 3370 3338 3406 3341
rect 3490 3338 3510 3341
rect 3514 3338 3534 3341
rect 3538 3338 3558 3341
rect 3562 3338 3582 3341
rect 3586 3338 3622 3341
rect 3626 3338 3646 3341
rect 3686 3338 3694 3341
rect 3698 3338 3774 3341
rect 4210 3338 4294 3341
rect 4314 3338 4318 3341
rect 4322 3338 4398 3341
rect 646 3332 649 3338
rect 1014 3332 1017 3338
rect 1110 3332 1113 3338
rect 2910 3332 2913 3338
rect 2958 3332 2961 3338
rect 114 3328 190 3331
rect 378 3328 470 3331
rect 682 3328 710 3331
rect 1234 3328 1358 3331
rect 1362 3328 1422 3331
rect 1426 3328 1526 3331
rect 1530 3328 1566 3331
rect 1898 3328 1990 3331
rect 2026 3328 2054 3331
rect 2114 3328 2358 3331
rect 2370 3328 2374 3331
rect 2402 3328 2526 3331
rect 2530 3328 2558 3331
rect 2802 3328 2870 3331
rect 2966 3328 3022 3331
rect 3246 3328 3262 3331
rect 3322 3328 3326 3331
rect 3354 3328 3382 3331
rect 3458 3328 3510 3331
rect 3514 3328 3670 3331
rect 3674 3328 3702 3331
rect 3938 3328 4030 3331
rect 4034 3328 4129 3331
rect 4274 3328 4478 3331
rect 4482 3328 4534 3331
rect 186 3318 230 3321
rect 270 3321 273 3328
rect 726 3322 729 3328
rect 2694 3322 2697 3328
rect 270 3318 318 3321
rect 322 3318 358 3321
rect 362 3318 398 3321
rect 410 3318 438 3321
rect 602 3318 614 3321
rect 994 3318 1030 3321
rect 1210 3318 1222 3321
rect 1322 3318 1502 3321
rect 1682 3318 2049 3321
rect 2130 3318 2254 3321
rect 2282 3318 2286 3321
rect 2370 3318 2374 3321
rect 2382 3318 2486 3321
rect 2786 3318 2790 3321
rect 2834 3318 2838 3321
rect 2966 3321 2969 3328
rect 3126 3322 3129 3328
rect 3206 3322 3209 3328
rect 3246 3322 3249 3328
rect 3310 3322 3313 3328
rect 4126 3322 4129 3328
rect 2882 3318 2969 3321
rect 2978 3318 2998 3321
rect 3034 3318 3054 3321
rect 3066 3318 3070 3321
rect 3330 3318 3750 3321
rect 438 3312 441 3318
rect 798 3312 801 3318
rect 298 3308 422 3311
rect 538 3308 774 3311
rect 1130 3308 1574 3311
rect 1690 3308 1702 3311
rect 2046 3311 2049 3318
rect 2046 3308 2214 3311
rect 2382 3311 2385 3318
rect 2550 3312 2553 3318
rect 2630 3312 2633 3318
rect 3166 3312 3169 3318
rect 2282 3308 2385 3311
rect 2394 3308 2398 3311
rect 2706 3308 2710 3311
rect 2850 3308 2878 3311
rect 2898 3308 2910 3311
rect 3130 3308 3142 3311
rect 3186 3308 3230 3311
rect 3522 3308 3702 3311
rect 4322 3308 4366 3311
rect 4482 3308 4494 3311
rect 4506 3308 4510 3311
rect 1000 3303 1002 3307
rect 1006 3303 1009 3307
rect 1014 3303 1016 3307
rect 2024 3303 2026 3307
rect 2030 3303 2033 3307
rect 2038 3303 2040 3307
rect 2886 3302 2889 3308
rect 2934 3302 2937 3308
rect 3048 3303 3050 3307
rect 3054 3303 3057 3307
rect 3062 3303 3064 3307
rect 4080 3303 4082 3307
rect 4086 3303 4089 3307
rect 4094 3303 4096 3307
rect 74 3298 174 3301
rect 610 3298 654 3301
rect 698 3298 742 3301
rect 1450 3298 1822 3301
rect 1826 3298 1926 3301
rect 2058 3298 2126 3301
rect 2170 3298 2342 3301
rect 2362 3298 2462 3301
rect 2514 3298 2566 3301
rect 2906 3298 2926 3301
rect 3106 3298 3222 3301
rect 3306 3298 3646 3301
rect 3954 3298 3982 3301
rect 3986 3298 4025 3301
rect 4498 3298 4558 3301
rect 234 3288 262 3291
rect 266 3288 302 3291
rect 306 3288 382 3291
rect 626 3288 718 3291
rect 722 3288 750 3291
rect 1234 3288 1398 3291
rect 1442 3288 1494 3291
rect 1498 3288 1662 3291
rect 1810 3288 1830 3291
rect 1834 3288 1902 3291
rect 1906 3288 1934 3291
rect 2018 3288 2022 3291
rect 2098 3288 2190 3291
rect 2290 3288 2294 3291
rect 2386 3288 2470 3291
rect 2538 3288 2633 3291
rect 2642 3288 2974 3291
rect 3026 3288 3102 3291
rect 3114 3288 3390 3291
rect 4022 3291 4025 3298
rect 4022 3288 4342 3291
rect 4394 3288 4566 3291
rect 2630 3282 2633 3288
rect 242 3278 393 3281
rect 402 3278 454 3281
rect 498 3278 510 3281
rect 1290 3278 1430 3281
rect 1482 3278 1518 3281
rect 1922 3278 2174 3281
rect 2186 3278 2406 3281
rect 2938 3278 2942 3281
rect 2986 3278 3094 3281
rect 3250 3278 3342 3281
rect 3354 3278 3406 3281
rect 3426 3278 3430 3281
rect 3530 3278 3662 3281
rect 3702 3281 3705 3288
rect 3674 3278 3705 3281
rect 3862 3281 3865 3288
rect 4014 3281 4017 3288
rect 3862 3278 4017 3281
rect 4370 3278 4526 3281
rect 66 3268 110 3271
rect 242 3268 294 3271
rect 322 3268 326 3271
rect 390 3271 393 3278
rect 390 3268 446 3271
rect 450 3268 470 3271
rect 490 3268 545 3271
rect 818 3268 854 3271
rect 1266 3268 1486 3271
rect 1514 3268 1926 3271
rect 1938 3268 2062 3271
rect 2218 3268 2225 3271
rect 2250 3268 2254 3271
rect 2346 3268 2422 3271
rect 2466 3268 2470 3271
rect 2570 3268 2614 3271
rect 2618 3268 2638 3271
rect 2666 3268 2670 3271
rect 2674 3268 2718 3271
rect 2870 3268 2910 3271
rect 2946 3268 2982 3271
rect 3066 3268 3102 3271
rect 3150 3271 3153 3278
rect 4214 3272 4217 3278
rect 3150 3268 3182 3271
rect 3186 3268 3262 3271
rect 3298 3268 3302 3271
rect 3314 3268 3398 3271
rect 3402 3268 3894 3271
rect 3994 3268 4118 3271
rect 4122 3268 4214 3271
rect 4250 3268 4262 3271
rect 90 3258 129 3261
rect 210 3258 270 3261
rect 310 3261 313 3268
rect 542 3262 545 3268
rect 290 3258 313 3261
rect 370 3258 374 3261
rect 786 3258 814 3261
rect 1190 3261 1193 3268
rect 2222 3262 2225 3268
rect 2870 3262 2873 3268
rect 2910 3262 2913 3268
rect 2942 3262 2945 3268
rect 3278 3262 3281 3268
rect 1190 3258 1238 3261
rect 1242 3258 1334 3261
rect 1378 3258 1422 3261
rect 1442 3258 1470 3261
rect 1554 3258 1654 3261
rect 1658 3258 1734 3261
rect 1738 3258 1774 3261
rect 1790 3258 1862 3261
rect 1866 3258 1950 3261
rect 2258 3258 2262 3261
rect 2306 3258 2574 3261
rect 2602 3258 2606 3261
rect 2618 3258 2670 3261
rect 2714 3258 2750 3261
rect 2962 3258 2966 3261
rect 2994 3258 3078 3261
rect 3138 3258 3214 3261
rect 3218 3258 3230 3261
rect 3234 3258 3254 3261
rect 3406 3258 3414 3261
rect 3418 3258 3505 3261
rect 3698 3258 3702 3261
rect 4026 3258 4214 3261
rect 4258 3258 4278 3261
rect 4366 3261 4369 3268
rect 4526 3262 4529 3268
rect 4366 3258 4414 3261
rect 126 3252 129 3258
rect 1790 3252 1793 3258
rect 2094 3252 2097 3258
rect 3502 3252 3505 3258
rect 218 3248 230 3251
rect 298 3248 558 3251
rect 626 3248 790 3251
rect 794 3248 838 3251
rect 842 3248 1350 3251
rect 1378 3248 1382 3251
rect 1434 3248 1774 3251
rect 2226 3248 2350 3251
rect 2394 3248 2414 3251
rect 2418 3248 2470 3251
rect 2514 3248 2542 3251
rect 2546 3248 2646 3251
rect 2650 3248 2678 3251
rect 2682 3248 2766 3251
rect 2858 3248 2918 3251
rect 2922 3248 2942 3251
rect 3010 3248 3022 3251
rect 3026 3248 3118 3251
rect 3218 3248 3286 3251
rect 3290 3248 3310 3251
rect 3610 3248 3798 3251
rect 4250 3248 4257 3251
rect 4546 3248 4566 3251
rect 4254 3242 4257 3248
rect 346 3238 382 3241
rect 714 3238 958 3241
rect 1442 3238 1710 3241
rect 1890 3238 2390 3241
rect 2418 3238 2454 3241
rect 2594 3238 2614 3241
rect 2634 3238 2638 3241
rect 2714 3238 2822 3241
rect 2826 3238 2846 3241
rect 2850 3238 2894 3241
rect 2970 3238 3014 3241
rect 3090 3238 3174 3241
rect 3178 3238 3198 3241
rect 3562 3238 3670 3241
rect 4266 3238 4430 3241
rect 762 3228 790 3231
rect 962 3228 1342 3231
rect 1410 3228 1630 3231
rect 1882 3228 2206 3231
rect 2218 3228 2798 3231
rect 3198 3231 3201 3238
rect 3198 3228 3366 3231
rect 3442 3228 3446 3231
rect 3458 3228 4390 3231
rect 106 3218 214 3221
rect 666 3218 790 3221
rect 810 3218 2742 3221
rect 2754 3218 2806 3221
rect 2826 3218 2862 3221
rect 2882 3218 3222 3221
rect 3522 3218 3566 3221
rect 3570 3218 3662 3221
rect 3666 3218 3718 3221
rect 3722 3218 3766 3221
rect 4106 3218 4326 3221
rect 730 3208 766 3211
rect 770 3208 1038 3211
rect 1042 3208 1102 3211
rect 1122 3208 1158 3211
rect 1410 3208 1414 3211
rect 1578 3208 1606 3211
rect 1986 3208 2142 3211
rect 2162 3208 2246 3211
rect 2330 3208 2398 3211
rect 2402 3208 2494 3211
rect 2578 3208 2622 3211
rect 2682 3208 2694 3211
rect 2698 3208 2734 3211
rect 2738 3208 2822 3211
rect 2826 3208 2854 3211
rect 2906 3208 2966 3211
rect 2970 3208 3038 3211
rect 3042 3208 3110 3211
rect 3114 3208 3134 3211
rect 3162 3208 3270 3211
rect 4226 3208 4326 3211
rect 496 3203 498 3207
rect 502 3203 505 3207
rect 510 3203 512 3207
rect 1478 3202 1481 3208
rect 1520 3203 1522 3207
rect 1526 3203 1529 3207
rect 1534 3203 1536 3207
rect 2544 3203 2546 3207
rect 2550 3203 2553 3207
rect 2558 3203 2560 3207
rect 3568 3203 3570 3207
rect 3574 3203 3577 3207
rect 3582 3203 3584 3207
rect 922 3198 1414 3201
rect 1954 3198 1974 3201
rect 2210 3198 2286 3201
rect 2314 3198 2342 3201
rect 2354 3198 2358 3201
rect 2370 3198 2502 3201
rect 2578 3198 2726 3201
rect 2730 3198 2798 3201
rect 2802 3198 2990 3201
rect 2994 3198 3230 3201
rect 3234 3198 3294 3201
rect 4074 3198 4406 3201
rect 986 3188 1017 3191
rect 1014 3182 1017 3188
rect 1102 3188 1550 3191
rect 1586 3188 2158 3191
rect 2194 3188 2814 3191
rect 2858 3188 2878 3191
rect 3226 3188 3710 3191
rect 3778 3188 3958 3191
rect 3962 3188 4142 3191
rect 4194 3188 4206 3191
rect 1102 3182 1105 3188
rect 238 3178 246 3181
rect 250 3178 694 3181
rect 1466 3178 1553 3181
rect 1550 3172 1553 3178
rect 2146 3178 2230 3181
rect 2274 3178 2598 3181
rect 2602 3178 2806 3181
rect 3034 3178 3158 3181
rect 3178 3178 3182 3181
rect 3226 3178 3286 3181
rect 4406 3181 4409 3188
rect 4010 3178 4073 3181
rect 4406 3178 4430 3181
rect -26 3168 -22 3172
rect 34 3168 38 3171
rect 42 3168 86 3171
rect 90 3168 238 3171
rect 242 3168 294 3171
rect 298 3168 302 3171
rect 338 3168 350 3171
rect 770 3168 814 3171
rect 1630 3171 1633 3178
rect 2838 3172 2841 3178
rect 2918 3172 2921 3178
rect 4070 3172 4073 3178
rect 1630 3168 1694 3171
rect 1722 3168 1838 3171
rect 2074 3168 2166 3171
rect 2178 3168 2206 3171
rect 2314 3168 2438 3171
rect 2458 3168 2462 3171
rect 2482 3168 2486 3171
rect 2498 3168 2510 3171
rect 2534 3168 2662 3171
rect 2738 3168 2774 3171
rect 3018 3168 3022 3171
rect 3106 3168 3110 3171
rect 3154 3168 3158 3171
rect 3170 3168 3254 3171
rect 4266 3168 4534 3171
rect -26 3161 -23 3168
rect -26 3158 102 3161
rect 202 3158 238 3161
rect 258 3158 270 3161
rect 282 3158 342 3161
rect 386 3158 406 3161
rect 1334 3161 1337 3168
rect 1414 3161 1417 3168
rect 1334 3158 1417 3161
rect 1602 3158 1654 3161
rect 2222 3161 2225 3168
rect 2090 3158 2225 3161
rect 2230 3161 2233 3168
rect 2254 3161 2257 3168
rect 2230 3158 2257 3161
rect 2534 3161 2537 3168
rect 2402 3158 2537 3161
rect 2546 3158 2630 3161
rect 2650 3158 2654 3161
rect 2666 3158 2670 3161
rect 2782 3161 2785 3168
rect 2762 3158 2785 3161
rect 2834 3158 3278 3161
rect 3686 3161 3689 3168
rect 3686 3158 3822 3161
rect 3882 3158 3950 3161
rect 3954 3158 4198 3161
rect 4262 3161 4265 3168
rect 4262 3158 4286 3161
rect 4414 3158 4446 3161
rect 4554 3158 4566 3161
rect 4570 3158 4590 3161
rect -26 3148 -22 3152
rect 18 3148 30 3151
rect 66 3148 78 3151
rect 146 3148 150 3151
rect 194 3148 254 3151
rect 258 3148 294 3151
rect 298 3148 326 3151
rect 346 3148 374 3151
rect 402 3148 446 3151
rect 450 3148 470 3151
rect 490 3148 502 3151
rect 566 3151 569 3158
rect 538 3148 569 3151
rect 730 3148 798 3151
rect 1150 3151 1153 3158
rect 1806 3152 1809 3158
rect 1018 3148 1153 3151
rect 1258 3148 1510 3151
rect 1530 3148 1590 3151
rect 1594 3148 1625 3151
rect 1658 3148 1686 3151
rect 1698 3148 1726 3151
rect 1918 3151 1921 3158
rect 2382 3152 2385 3158
rect 1918 3148 1990 3151
rect -26 3141 -23 3148
rect 1622 3142 1625 3148
rect 2010 3148 2062 3151
rect 2066 3148 2185 3151
rect 2266 3148 2294 3151
rect 2298 3148 2318 3151
rect 2338 3148 2358 3151
rect 2410 3148 2414 3151
rect 2482 3148 2622 3151
rect 2650 3148 2854 3151
rect 2866 3148 2870 3151
rect 2882 3148 3238 3151
rect 3258 3148 3286 3151
rect 3290 3148 3302 3151
rect 3306 3148 3350 3151
rect 3354 3148 3374 3151
rect 3574 3151 3577 3158
rect 4414 3152 4417 3158
rect 3562 3148 3577 3151
rect 3666 3148 3678 3151
rect 3682 3148 3734 3151
rect 3754 3148 3894 3151
rect -26 3138 6 3141
rect 130 3138 150 3141
rect 186 3138 190 3141
rect 262 3138 278 3141
rect 354 3138 366 3141
rect 386 3138 422 3141
rect 426 3138 454 3141
rect 530 3138 681 3141
rect 962 3138 1022 3141
rect 1546 3138 1606 3141
rect 2082 3138 2086 3141
rect 2106 3138 2166 3141
rect 2170 3138 2174 3141
rect 2182 3141 2185 3148
rect 3918 3148 3966 3151
rect 4082 3148 4278 3151
rect 4330 3148 4334 3151
rect 4482 3148 4502 3151
rect 4506 3148 4510 3151
rect 3918 3142 3921 3148
rect 4046 3142 4049 3148
rect 4438 3142 4441 3148
rect 2182 3138 2302 3141
rect 2466 3138 2494 3141
rect 2514 3138 2598 3141
rect 2618 3138 2622 3141
rect 2666 3138 2742 3141
rect 2746 3138 2806 3141
rect 2810 3138 2886 3141
rect 2946 3138 2974 3141
rect 3018 3138 3054 3141
rect 3250 3138 3313 3141
rect 3362 3138 3430 3141
rect 3498 3138 3670 3141
rect 4298 3138 4350 3141
rect 4354 3138 4374 3141
rect 4410 3138 4422 3141
rect 4466 3138 4486 3141
rect 4490 3138 4510 3141
rect 4562 3138 4566 3141
rect 262 3132 265 3138
rect 582 3132 585 3138
rect 678 3132 681 3138
rect 1406 3132 1409 3138
rect 3310 3132 3313 3138
rect 4118 3132 4121 3138
rect -26 3128 -22 3132
rect 50 3128 94 3131
rect 98 3128 246 3131
rect 314 3128 334 3131
rect 338 3128 430 3131
rect 458 3128 550 3131
rect 954 3128 1334 3131
rect 1554 3128 1566 3131
rect 1578 3128 1614 3131
rect 1994 3128 2094 3131
rect 2098 3128 2150 3131
rect 2162 3128 2182 3131
rect 2346 3128 2350 3131
rect 2434 3128 2494 3131
rect 2530 3128 2678 3131
rect 2802 3128 2838 3131
rect 2874 3128 2878 3131
rect 2938 3128 2942 3131
rect 2986 3128 2990 3131
rect 2994 3128 3134 3131
rect 3186 3128 3246 3131
rect 3642 3128 3750 3131
rect 4122 3128 4350 3131
rect -26 3121 -23 3128
rect 2846 3122 2849 3128
rect -26 3118 54 3121
rect 258 3118 262 3121
rect 370 3118 406 3121
rect 514 3118 542 3121
rect 666 3118 670 3121
rect 770 3118 886 3121
rect 890 3118 1302 3121
rect 1322 3118 1390 3121
rect 1554 3118 1566 3121
rect 1570 3118 1606 3121
rect 1610 3118 1646 3121
rect 1682 3118 2190 3121
rect 2402 3118 2417 3121
rect 2466 3118 2470 3121
rect 2482 3118 2486 3121
rect 2498 3118 2542 3121
rect 2626 3118 2742 3121
rect 2770 3118 2774 3121
rect 2890 3118 2942 3121
rect 3034 3118 3086 3121
rect 3170 3118 3254 3121
rect 3298 3118 3502 3121
rect 3506 3118 3982 3121
rect 4082 3118 4177 3121
rect 2414 3112 2417 3118
rect 4174 3112 4177 3118
rect 178 3108 262 3111
rect 266 3108 318 3111
rect 322 3108 430 3111
rect 442 3108 598 3111
rect 786 3108 814 3111
rect 858 3108 934 3111
rect 1490 3108 1590 3111
rect 1594 3108 1686 3111
rect 1690 3108 1718 3111
rect 2146 3108 2174 3111
rect 2282 3108 2310 3111
rect 2346 3108 2358 3111
rect 2442 3108 2510 3111
rect 2698 3108 2734 3111
rect 2754 3108 2774 3111
rect 3098 3108 3254 3111
rect 3298 3108 3470 3111
rect 3642 3108 3646 3111
rect 4178 3108 4270 3111
rect 4274 3108 4294 3111
rect 4442 3108 4446 3111
rect 1000 3103 1002 3107
rect 1006 3103 1009 3107
rect 1014 3103 1016 3107
rect 2024 3103 2026 3107
rect 2030 3103 2033 3107
rect 2038 3103 2040 3107
rect 2646 3102 2649 3108
rect 3048 3103 3050 3107
rect 3054 3103 3057 3107
rect 3062 3103 3064 3107
rect 4080 3103 4082 3107
rect 4086 3103 4089 3107
rect 4094 3103 4096 3107
rect 402 3098 702 3101
rect 834 3098 958 3101
rect 1562 3098 1694 3101
rect 2130 3098 2150 3101
rect 2266 3098 2294 3101
rect 2298 3098 2318 3101
rect 2322 3098 2382 3101
rect 2386 3098 2582 3101
rect 2698 3098 2702 3101
rect 2738 3098 2830 3101
rect 2866 3098 2894 3101
rect 3034 3098 3041 3101
rect 3258 3098 3606 3101
rect 4282 3098 4302 3101
rect 4394 3098 4486 3101
rect 1294 3092 1297 3098
rect 1790 3092 1793 3098
rect 154 3088 182 3091
rect 250 3088 326 3091
rect 778 3088 854 3091
rect 858 3088 998 3091
rect 1442 3088 1486 3091
rect 1522 3088 1606 3091
rect 1882 3088 1886 3091
rect 1994 3088 1998 3091
rect 2074 3088 2238 3091
rect 2258 3088 2294 3091
rect 2322 3088 2374 3091
rect 2394 3088 2438 3091
rect 2442 3088 2846 3091
rect 3038 3091 3041 3098
rect 3038 3088 3054 3091
rect 3130 3088 3230 3091
rect 3274 3088 3350 3091
rect 4154 3088 4438 3091
rect 226 3078 246 3081
rect 326 3081 329 3088
rect 326 3078 398 3081
rect 690 3078 694 3081
rect 754 3078 766 3081
rect 1106 3078 1326 3081
rect 1458 3078 1670 3081
rect 2154 3078 2182 3081
rect 2186 3078 2214 3081
rect 2274 3078 2526 3081
rect 2538 3078 2678 3081
rect 2682 3078 2822 3081
rect 2854 3081 2857 3088
rect 3030 3082 3033 3088
rect 2854 3078 2910 3081
rect 3074 3078 3094 3081
rect 3154 3078 3158 3081
rect 3178 3078 3214 3081
rect 3330 3078 3510 3081
rect 3514 3078 3686 3081
rect 4114 3078 4270 3081
rect 4410 3078 4566 3081
rect 6 3072 9 3078
rect 42 3068 78 3071
rect 338 3068 390 3071
rect 570 3068 574 3071
rect 578 3068 830 3071
rect 1386 3068 1390 3071
rect 1402 3068 1542 3071
rect 1678 3071 1681 3078
rect 2254 3072 2257 3078
rect 1678 3068 1726 3071
rect 1762 3068 2078 3071
rect 2162 3068 2254 3071
rect 2258 3068 2310 3071
rect 2322 3068 2414 3071
rect 2426 3068 2438 3071
rect 2482 3068 2486 3071
rect 2522 3068 2558 3071
rect 2602 3068 2606 3071
rect 2610 3068 2646 3071
rect 2878 3068 2894 3071
rect 2898 3068 2902 3071
rect 2994 3068 3078 3071
rect 3114 3068 3198 3071
rect 3282 3068 3294 3071
rect 3362 3068 3382 3071
rect 3466 3068 3486 3071
rect 3546 3068 3702 3071
rect 3998 3071 4001 3078
rect 3998 3068 4150 3071
rect 4390 3071 4393 3078
rect 4282 3068 4393 3071
rect 4458 3068 4478 3071
rect 4482 3068 4510 3071
rect 4538 3068 4542 3071
rect 18 3058 30 3061
rect 174 3061 177 3068
rect 162 3058 177 3061
rect 262 3058 286 3061
rect 546 3058 590 3061
rect 594 3058 750 3061
rect 762 3058 774 3061
rect 862 3061 865 3068
rect 794 3058 910 3061
rect 914 3058 1022 3061
rect 1374 3061 1377 3068
rect 1354 3058 1518 3061
rect 1562 3058 1582 3061
rect 1850 3059 1854 3061
rect 1846 3058 1854 3059
rect 2878 3062 2881 3068
rect 2042 3059 2046 3061
rect 2038 3058 2046 3059
rect 2114 3058 2174 3061
rect 2178 3058 2198 3061
rect 2298 3058 2358 3061
rect 2426 3058 2454 3061
rect 2554 3058 2566 3061
rect 2650 3058 2654 3061
rect 2914 3058 2918 3061
rect 3002 3058 3006 3061
rect 3010 3058 3022 3061
rect 3066 3058 3110 3061
rect 3114 3058 3118 3061
rect 3178 3058 3182 3061
rect 3210 3058 3214 3061
rect 3242 3058 3486 3061
rect 3506 3058 3518 3061
rect 3538 3058 3617 3061
rect 3634 3058 3726 3061
rect 3802 3058 3878 3061
rect 4098 3058 4118 3061
rect 4170 3058 4302 3061
rect 4490 3058 4534 3061
rect 4538 3058 4582 3061
rect 262 3052 265 3058
rect 3142 3052 3145 3058
rect 3614 3052 3617 3058
rect -26 3051 -22 3052
rect -26 3048 6 3051
rect 114 3048 190 3051
rect 274 3048 278 3051
rect 330 3048 342 3051
rect 402 3048 486 3051
rect 522 3048 598 3051
rect 602 3048 630 3051
rect 658 3048 662 3051
rect 706 3048 710 3051
rect 754 3048 766 3051
rect 1326 3048 1454 3051
rect 1546 3048 1558 3051
rect 1642 3048 1846 3051
rect 1954 3048 2198 3051
rect 2206 3048 2214 3051
rect 2290 3048 2297 3051
rect 2362 3048 2366 3051
rect 2438 3048 2470 3051
rect 2522 3048 2606 3051
rect 2610 3048 2630 3051
rect 2634 3048 2662 3051
rect 2682 3048 2710 3051
rect 2714 3048 2742 3051
rect 2914 3048 2918 3051
rect 2978 3048 3006 3051
rect 3034 3048 3110 3051
rect 3170 3048 3182 3051
rect 3194 3048 3222 3051
rect 3226 3048 3238 3051
rect 3274 3048 3310 3051
rect 3322 3048 3510 3051
rect 4066 3048 4158 3051
rect 4290 3048 4350 3051
rect 4370 3048 4374 3051
rect 4470 3048 4518 3051
rect 34 3038 38 3041
rect 306 3038 310 3041
rect 626 3038 678 3041
rect 990 3041 993 3048
rect 1326 3042 1329 3048
rect 2294 3042 2297 3048
rect 2438 3042 2441 3048
rect 4470 3042 4473 3048
rect 990 3038 1046 3041
rect 1382 3038 1414 3041
rect 2122 3038 2166 3041
rect 2534 3038 2590 3041
rect 2706 3038 2726 3041
rect 2730 3038 2790 3041
rect 2842 3038 2862 3041
rect 2866 3038 2974 3041
rect 3018 3038 3030 3041
rect 3034 3038 3046 3041
rect 3122 3038 3126 3041
rect 3370 3038 3454 3041
rect 3458 3038 4030 3041
rect 4322 3038 4462 3041
rect 4530 3038 4534 3041
rect 150 3032 153 3038
rect 1382 3032 1385 3038
rect 2534 3032 2537 3038
rect 274 3028 430 3031
rect 786 3028 838 3031
rect 842 3028 1014 3031
rect 1762 3028 2062 3031
rect 2162 3028 2238 3031
rect 2290 3028 2318 3031
rect 2730 3028 2766 3031
rect 2770 3028 2822 3031
rect 2842 3028 2846 3031
rect 2906 3028 2934 3031
rect 3042 3028 3182 3031
rect 3394 3028 4254 3031
rect 4282 3028 4446 3031
rect 4562 3028 4574 3031
rect 754 3018 758 3021
rect 1586 3018 2118 3021
rect 2122 3018 2214 3021
rect 2250 3018 2486 3021
rect 2762 3018 3406 3021
rect 3490 3018 3673 3021
rect 3682 3018 3686 3021
rect 3690 3018 4206 3021
rect 1666 3008 1873 3011
rect 2210 3008 2406 3011
rect 2410 3008 2534 3011
rect 2778 3008 3470 3011
rect 3670 3011 3673 3018
rect 3670 3008 3710 3011
rect 496 3003 498 3007
rect 502 3003 505 3007
rect 510 3003 512 3007
rect 1520 3003 1522 3007
rect 1526 3003 1529 3007
rect 1534 3003 1536 3007
rect 378 2998 398 3001
rect 522 2998 630 3001
rect 634 2998 646 3001
rect 650 2998 782 3001
rect 1186 2998 1230 3001
rect 1282 2998 1286 3001
rect 1450 2998 1494 3001
rect 1858 2998 1862 3001
rect 1870 3001 1873 3008
rect 2544 3003 2546 3007
rect 2550 3003 2553 3007
rect 2558 3003 2560 3007
rect 3568 3003 3570 3007
rect 3574 3003 3577 3007
rect 3582 3003 3584 3007
rect 1870 2998 2134 3001
rect 2138 2998 2166 3001
rect 2178 2998 2190 3001
rect 2314 2998 2390 3001
rect 2890 2998 2934 3001
rect 3146 2998 3286 3001
rect 122 2988 158 2991
rect 162 2988 702 2991
rect 746 2988 790 2991
rect 1170 2988 2758 2991
rect 3106 2988 3270 2991
rect 3290 2988 3462 2991
rect 3466 2988 3934 2991
rect 402 2978 494 2981
rect 642 2978 654 2981
rect 658 2978 678 2981
rect 682 2978 726 2981
rect 730 2978 782 2981
rect 786 2978 798 2981
rect 802 2978 822 2981
rect 1370 2978 1649 2981
rect 1666 2978 2206 2981
rect 2238 2978 2262 2981
rect 2310 2978 2334 2981
rect 2346 2978 2590 2981
rect 2594 2978 3478 2981
rect 3666 2978 3742 2981
rect 4122 2978 4558 2981
rect 346 2968 438 2971
rect 442 2968 526 2971
rect 610 2968 926 2971
rect 1418 2968 1462 2971
rect 1646 2971 1649 2978
rect 1646 2968 1814 2971
rect 2238 2971 2241 2978
rect 2310 2972 2313 2978
rect 1906 2968 2241 2971
rect 2250 2968 2262 2971
rect 2378 2968 2414 2971
rect 3026 2968 3030 2971
rect 3338 2968 3646 2971
rect 3698 2968 3854 2971
rect 3858 2968 3998 2971
rect 4514 2968 4566 2971
rect 4570 2968 4574 2971
rect 314 2958 406 2961
rect 534 2961 537 2968
rect 534 2958 542 2961
rect 746 2958 750 2961
rect 986 2958 1070 2961
rect 1090 2958 2566 2961
rect 2754 2958 2769 2961
rect 2786 2958 2798 2961
rect 2914 2958 2918 2961
rect 2922 2958 2926 2961
rect 2930 2958 3230 2961
rect 3250 2958 3854 2961
rect 4322 2958 4326 2961
rect 4410 2958 4422 2961
rect -26 2951 -22 2952
rect -26 2948 6 2951
rect 250 2948 566 2951
rect 650 2948 662 2951
rect 670 2951 673 2958
rect 710 2951 713 2958
rect 2766 2952 2769 2958
rect 4550 2952 4553 2958
rect 670 2948 734 2951
rect 738 2948 798 2951
rect 994 2948 1222 2951
rect 1226 2948 1230 2951
rect 1398 2948 1422 2951
rect 14 2941 17 2948
rect 14 2938 150 2941
rect 650 2938 678 2941
rect 754 2938 790 2941
rect 894 2941 897 2948
rect 910 2941 913 2948
rect 1398 2942 1401 2948
rect 1530 2948 1534 2951
rect 2034 2948 2134 2951
rect 894 2938 913 2941
rect 994 2938 1062 2941
rect 1550 2941 1553 2948
rect 2014 2942 2017 2948
rect 2226 2948 2230 2951
rect 2402 2948 2430 2951
rect 2466 2948 2502 2951
rect 2510 2948 2518 2951
rect 2522 2948 2534 2951
rect 2538 2948 2614 2951
rect 2690 2948 2758 2951
rect 3362 2948 3393 2951
rect 3418 2948 3510 2951
rect 3514 2948 3630 2951
rect 3674 2948 3702 2951
rect 3706 2948 3718 2951
rect 4298 2948 4326 2951
rect 4354 2948 4406 2951
rect 3390 2942 3393 2948
rect 1550 2938 1678 2941
rect 1682 2938 1734 2941
rect 2030 2938 2062 2941
rect 2114 2938 2118 2941
rect 2154 2938 2158 2941
rect 2202 2938 2270 2941
rect 2282 2938 2286 2941
rect 2386 2938 2454 2941
rect 2490 2938 2566 2941
rect 2610 2938 2630 2941
rect 2634 2938 2670 2941
rect 2674 2938 2710 2941
rect 2842 2938 2982 2941
rect 2998 2938 3038 2941
rect 3098 2938 3134 2941
rect 3138 2938 3174 2941
rect 3298 2938 3318 2941
rect 3322 2938 3342 2941
rect 3538 2938 3566 2941
rect 3714 2938 3782 2941
rect 4166 2941 4169 2948
rect 4182 2941 4185 2948
rect 4166 2938 4254 2941
rect 4274 2938 4286 2941
rect 4322 2938 4334 2941
rect 4546 2938 4566 2941
rect 2030 2932 2033 2938
rect 2998 2932 3001 2938
rect 178 2928 318 2931
rect 570 2928 598 2931
rect 666 2928 718 2931
rect 1074 2928 1078 2931
rect 1410 2928 1662 2931
rect 2122 2928 2350 2931
rect 2386 2928 2398 2931
rect 2446 2928 2478 2931
rect 2498 2928 2510 2931
rect 2522 2928 2806 2931
rect 2810 2928 2854 2931
rect 3010 2928 3030 2931
rect 3074 2928 3078 2931
rect 3082 2928 3110 2931
rect 3162 2928 3190 2931
rect 3242 2928 3326 2931
rect 4034 2928 4398 2931
rect 4462 2931 4465 2938
rect 4518 2931 4521 2938
rect 4462 2928 4521 2931
rect 158 2918 166 2921
rect 170 2918 310 2921
rect 614 2921 617 2928
rect 2446 2922 2449 2928
rect 614 2918 702 2921
rect 938 2918 1606 2921
rect 1890 2918 1910 2921
rect 1914 2918 2438 2921
rect 2458 2918 2750 2921
rect 2754 2918 2758 2921
rect 2914 2918 2958 2921
rect 2962 2918 3246 2921
rect 3274 2918 3510 2921
rect 3538 2918 3558 2921
rect 3562 2918 4198 2921
rect 4258 2918 4382 2921
rect 4386 2918 4454 2921
rect 466 2908 566 2911
rect 586 2908 654 2911
rect 658 2908 670 2911
rect 690 2908 774 2911
rect 778 2908 814 2911
rect 1082 2908 1166 2911
rect 1282 2908 1382 2911
rect 1674 2908 1694 2911
rect 2050 2908 2302 2911
rect 2402 2908 2414 2911
rect 2434 2908 2670 2911
rect 2690 2908 2886 2911
rect 2890 2908 2894 2911
rect 2962 2908 2966 2911
rect 3194 2908 3222 2911
rect 3226 2908 3246 2911
rect 3314 2908 3678 2911
rect 4242 2908 4310 2911
rect 4314 2908 4382 2911
rect 1000 2903 1002 2907
rect 1006 2903 1009 2907
rect 1014 2903 1016 2907
rect 2024 2903 2026 2907
rect 2030 2903 2033 2907
rect 2038 2903 2040 2907
rect 3048 2903 3050 2907
rect 3054 2903 3057 2907
rect 3062 2903 3064 2907
rect 3278 2902 3281 2908
rect 4080 2903 4082 2907
rect 4086 2903 4089 2907
rect 4094 2903 4096 2907
rect 306 2898 366 2901
rect 370 2898 478 2901
rect 482 2898 534 2901
rect 554 2898 614 2901
rect 618 2898 630 2901
rect 1066 2898 1086 2901
rect 1354 2898 1382 2901
rect 1450 2898 1574 2901
rect 1578 2898 1590 2901
rect 1634 2898 1846 2901
rect 1906 2898 1942 2901
rect 2050 2898 2054 2901
rect 2234 2898 2366 2901
rect 2650 2898 2670 2901
rect 2818 2898 3006 2901
rect 3082 2898 3198 2901
rect 3218 2898 3238 2901
rect 3346 2898 3454 2901
rect 3458 2898 3502 2901
rect 3506 2898 3526 2901
rect 3810 2898 3814 2901
rect 4362 2898 4558 2901
rect 694 2892 697 2898
rect 266 2888 334 2891
rect 442 2888 582 2891
rect 594 2888 638 2891
rect 658 2888 686 2891
rect 874 2888 886 2891
rect 1106 2888 1142 2891
rect 1370 2888 1382 2891
rect 1466 2888 1486 2891
rect 1666 2888 1790 2891
rect 1794 2888 1830 2891
rect 1842 2888 1910 2891
rect 1930 2888 2238 2891
rect 2354 2888 2430 2891
rect 2522 2888 2526 2891
rect 2850 2888 3254 2891
rect 3338 2888 3342 2891
rect 3498 2888 3862 2891
rect 4266 2888 4486 2891
rect 34 2878 62 2881
rect 74 2878 158 2881
rect 538 2878 590 2881
rect 602 2878 646 2881
rect 666 2878 870 2881
rect 874 2878 878 2881
rect 882 2878 918 2881
rect 1346 2878 1462 2881
rect 1594 2878 1774 2881
rect 1778 2878 1806 2881
rect 1826 2878 2150 2881
rect 2162 2878 2630 2881
rect 2866 2878 2966 2881
rect 3082 2878 3086 2881
rect 3302 2881 3305 2888
rect 3302 2878 3318 2881
rect 3690 2878 3918 2881
rect 4142 2881 4145 2888
rect 4142 2878 4342 2881
rect 4402 2878 4470 2881
rect -26 2871 -22 2872
rect -26 2868 86 2871
rect 114 2868 126 2871
rect 546 2868 710 2871
rect 810 2868 854 2871
rect 862 2868 910 2871
rect 958 2871 961 2878
rect 914 2868 961 2871
rect 1294 2871 1297 2878
rect 1226 2868 1297 2871
rect 1462 2871 1465 2878
rect 1462 2868 1550 2871
rect 1650 2868 1654 2871
rect 1770 2868 1830 2871
rect 1850 2868 1950 2871
rect 2218 2868 2350 2871
rect 2442 2868 2462 2871
rect 2634 2868 2726 2871
rect 2882 2868 2982 2871
rect 3266 2868 3350 2871
rect 3650 2868 3774 2871
rect 3850 2868 3966 2871
rect 4322 2868 4358 2871
rect 4362 2868 4422 2871
rect 4426 2868 4542 2871
rect 4582 2871 4585 2878
rect 4562 2868 4585 2871
rect 66 2858 142 2861
rect 146 2858 270 2861
rect 274 2858 286 2861
rect 482 2858 526 2861
rect 530 2858 550 2861
rect 594 2858 662 2861
rect 666 2858 686 2861
rect 706 2858 710 2861
rect 810 2858 814 2861
rect 862 2861 865 2868
rect 842 2858 865 2861
rect 890 2858 950 2861
rect 1034 2858 1038 2861
rect 1158 2858 1230 2861
rect 1558 2858 1582 2861
rect 1598 2861 1601 2868
rect 1598 2858 1622 2861
rect 1650 2858 1726 2861
rect 1730 2858 1798 2861
rect 2086 2861 2089 2868
rect 2026 2858 2134 2861
rect 2182 2861 2185 2868
rect 2138 2858 2185 2861
rect 2374 2861 2377 2868
rect 2502 2862 2505 2868
rect 2614 2862 2617 2868
rect 2758 2862 2761 2868
rect 2330 2858 2377 2861
rect 2426 2858 2470 2861
rect 2538 2858 2566 2861
rect 2594 2858 2606 2861
rect 2626 2858 2646 2861
rect 2650 2858 2678 2861
rect 2862 2861 2865 2868
rect 2842 2858 2865 2861
rect 2954 2858 3054 2861
rect 3058 2858 3070 2861
rect 3190 2861 3193 2868
rect 3146 2858 3193 2861
rect 3338 2858 3390 2861
rect 3518 2861 3521 2868
rect 3606 2861 3609 2868
rect 3518 2858 3609 2861
rect 3666 2858 3670 2861
rect 3706 2858 3726 2861
rect 3730 2858 3870 2861
rect 3874 2858 3910 2861
rect 4110 2861 4113 2868
rect 4598 2862 4601 2868
rect 4110 2858 4158 2861
rect 4330 2858 4398 2861
rect 4402 2858 4446 2861
rect 4450 2858 4550 2861
rect 4554 2858 4582 2861
rect 1158 2852 1161 2858
rect 1558 2852 1561 2858
rect 2310 2852 2313 2858
rect 2406 2852 2409 2858
rect -26 2851 -22 2852
rect -26 2848 6 2851
rect 114 2848 190 2851
rect 274 2848 366 2851
rect 434 2848 878 2851
rect 942 2848 966 2851
rect 1626 2848 1654 2851
rect 1738 2848 1758 2851
rect 1914 2848 2118 2851
rect 2618 2848 2673 2851
rect 2738 2848 2766 2851
rect 2770 2848 2774 2851
rect 2842 2848 2886 2851
rect 2930 2848 2953 2851
rect 2978 2848 3006 2851
rect 3010 2848 3094 2851
rect 3234 2848 3262 2851
rect 3266 2848 3294 2851
rect 3438 2851 3441 2858
rect 3306 2848 3441 2851
rect 3506 2848 3926 2851
rect 4378 2848 4414 2851
rect 4474 2848 4598 2851
rect 942 2842 945 2848
rect 2670 2842 2673 2848
rect 2950 2842 2953 2848
rect 402 2838 438 2841
rect 446 2838 494 2841
rect 498 2838 558 2841
rect 698 2838 742 2841
rect 950 2838 1046 2841
rect 1050 2838 2454 2841
rect 2570 2838 2598 2841
rect 2602 2838 2649 2841
rect 2738 2838 2790 2841
rect 2986 2838 3662 2841
rect 3730 2838 3758 2841
rect 3762 2838 3854 2841
rect 3858 2838 3950 2841
rect 4562 2838 4566 2841
rect 446 2832 449 2838
rect 542 2828 574 2831
rect 578 2828 598 2831
rect 818 2828 846 2831
rect 950 2831 953 2838
rect 850 2828 953 2831
rect 2010 2828 2086 2831
rect 2090 2828 2158 2831
rect 2354 2828 2422 2831
rect 2482 2828 2638 2831
rect 2646 2831 2649 2838
rect 2646 2828 2702 2831
rect 2706 2828 2806 2831
rect 2810 2828 2942 2831
rect 3210 2828 3398 2831
rect 3674 2828 3742 2831
rect 3746 2828 4270 2831
rect 542 2822 545 2828
rect 642 2818 686 2821
rect 1266 2818 1446 2821
rect 1450 2818 3246 2821
rect 3394 2818 4438 2821
rect 814 2812 817 2818
rect 2010 2808 2478 2811
rect 2578 2808 2710 2811
rect 3250 2808 3358 2811
rect 3986 2808 4078 2811
rect 496 2803 498 2807
rect 502 2803 505 2807
rect 510 2803 512 2807
rect 1520 2803 1522 2807
rect 1526 2803 1529 2807
rect 1534 2803 1536 2807
rect 2544 2803 2546 2807
rect 2550 2803 2553 2807
rect 2558 2803 2560 2807
rect 3568 2803 3570 2807
rect 3574 2803 3577 2807
rect 3582 2803 3584 2807
rect 954 2798 1486 2801
rect 2178 2798 2294 2801
rect 2578 2798 3334 2801
rect 3810 2798 3838 2801
rect 3842 2798 4238 2801
rect 474 2788 862 2791
rect 866 2788 894 2791
rect 1130 2788 1190 2791
rect 1194 2788 1406 2791
rect 2574 2791 2577 2798
rect 1410 2788 2577 2791
rect 3154 2788 4102 2791
rect 4106 2788 4174 2791
rect 1802 2778 1902 2781
rect 1978 2778 2046 2781
rect 2090 2778 2094 2781
rect 2202 2778 2254 2781
rect 2298 2778 2494 2781
rect 2522 2778 2545 2781
rect 2570 2778 2886 2781
rect 2938 2778 3006 2781
rect 3362 2778 3750 2781
rect 3754 2778 4462 2781
rect 2542 2772 2545 2778
rect 4598 2772 4601 2778
rect 1274 2768 1310 2771
rect 1482 2768 1518 2771
rect 1682 2768 1686 2771
rect 1762 2768 1902 2771
rect 1914 2768 2126 2771
rect 2850 2768 2870 2771
rect 2938 2768 2958 2771
rect 2962 2768 2966 2771
rect 2970 2768 3006 2771
rect 3010 2768 3030 2771
rect 3034 2768 3078 2771
rect 3162 2768 3246 2771
rect 3258 2768 3294 2771
rect 4002 2768 4030 2771
rect 350 2761 353 2768
rect 350 2758 462 2761
rect 614 2761 617 2768
rect 694 2762 697 2768
rect 2614 2762 2617 2768
rect 614 2758 622 2761
rect 770 2758 814 2761
rect 834 2758 1022 2761
rect 1282 2758 1310 2761
rect 1618 2758 1694 2761
rect 1698 2758 1750 2761
rect 1754 2758 1790 2761
rect 1810 2758 1862 2761
rect 1930 2758 2006 2761
rect 2114 2758 2486 2761
rect 2490 2758 2526 2761
rect 2698 2758 2702 2761
rect 2770 2758 2814 2761
rect 2818 2758 2974 2761
rect 2978 2758 3142 2761
rect 3226 2758 3366 2761
rect 3370 2758 3414 2761
rect 3646 2761 3649 2768
rect 3514 2758 3942 2761
rect 3946 2758 3998 2761
rect 4242 2758 4262 2761
rect 4266 2758 4310 2761
rect 4314 2758 4454 2761
rect 710 2752 713 2758
rect -26 2751 -22 2752
rect -26 2748 14 2751
rect 50 2748 142 2751
rect 258 2748 614 2751
rect 634 2748 638 2751
rect 658 2748 710 2751
rect 714 2748 734 2751
rect 738 2748 846 2751
rect 850 2748 862 2751
rect 898 2748 1126 2751
rect 1418 2748 1422 2751
rect 1602 2748 1662 2751
rect 1666 2748 1726 2751
rect 1730 2748 1774 2751
rect 1778 2748 1814 2751
rect 1822 2748 1886 2751
rect 614 2742 617 2748
rect 1822 2742 1825 2748
rect 26 2738 70 2741
rect 626 2738 670 2741
rect 874 2738 910 2741
rect 938 2738 1030 2741
rect 1034 2738 1105 2741
rect 1586 2738 1734 2741
rect 1990 2741 1993 2748
rect 2154 2748 2286 2751
rect 2330 2748 2334 2751
rect 2450 2748 2622 2751
rect 2906 2748 2934 2751
rect 3018 2748 3062 2751
rect 3138 2748 3190 2751
rect 3194 2748 3222 2751
rect 3242 2748 3281 2751
rect 3470 2751 3473 2758
rect 3458 2748 3473 2751
rect 3690 2748 3878 2751
rect 2310 2742 2313 2748
rect 3278 2742 3281 2748
rect 1990 2738 2022 2741
rect 2338 2738 2350 2741
rect 2354 2738 2366 2741
rect 2370 2738 2382 2741
rect 2386 2738 2406 2741
rect 2410 2738 2462 2741
rect 2602 2738 2646 2741
rect 2650 2738 2694 2741
rect 2698 2738 2726 2741
rect 2730 2738 2734 2741
rect 2810 2738 2830 2741
rect 2834 2738 2862 2741
rect 2866 2738 2886 2741
rect 3402 2738 3582 2741
rect 3662 2741 3665 2748
rect 3922 2748 4038 2751
rect 4082 2748 4142 2751
rect 4386 2748 4390 2751
rect 3602 2738 3665 2741
rect 3778 2738 3814 2741
rect 4130 2738 4206 2741
rect 4234 2738 4238 2741
rect 4242 2738 4278 2741
rect 4306 2738 4342 2741
rect 1102 2732 1105 2738
rect -26 2731 -22 2732
rect -26 2728 6 2731
rect 98 2728 158 2731
rect 658 2728 702 2731
rect 706 2728 718 2731
rect 1378 2728 1590 2731
rect 1746 2728 2014 2731
rect 2018 2728 2086 2731
rect 2090 2728 2110 2731
rect 2258 2728 2494 2731
rect 2738 2728 2990 2731
rect 3314 2728 3422 2731
rect 3426 2728 3502 2731
rect 3506 2728 3518 2731
rect 3522 2728 3566 2731
rect 3778 2728 3782 2731
rect 3786 2728 4038 2731
rect 4058 2728 4158 2731
rect 4290 2728 4302 2731
rect 74 2718 318 2721
rect 826 2718 1238 2721
rect 1682 2718 1742 2721
rect 1794 2718 1830 2721
rect 1866 2718 1894 2721
rect 2162 2718 2406 2721
rect 2594 2718 2814 2721
rect 2914 2718 3102 2721
rect 3434 2718 3798 2721
rect 3842 2718 3926 2721
rect 3930 2718 4318 2721
rect 694 2712 697 2718
rect 82 2708 190 2711
rect 722 2708 742 2711
rect 746 2708 846 2711
rect 850 2708 854 2711
rect 858 2708 878 2711
rect 1090 2708 1118 2711
rect 1466 2708 1758 2711
rect 2322 2708 2446 2711
rect 2466 2708 2614 2711
rect 2682 2708 2726 2711
rect 2994 2708 2998 2711
rect 3178 2708 3262 2711
rect 3362 2708 3742 2711
rect 4210 2708 4358 2711
rect 1000 2703 1002 2707
rect 1006 2703 1009 2707
rect 1014 2703 1016 2707
rect 2024 2703 2026 2707
rect 2030 2703 2033 2707
rect 2038 2703 2040 2707
rect 3048 2703 3050 2707
rect 3054 2703 3057 2707
rect 3062 2703 3064 2707
rect 4080 2703 4082 2707
rect 4086 2703 4089 2707
rect 4094 2703 4096 2707
rect 654 2698 702 2701
rect 1642 2698 1670 2701
rect 2058 2698 2374 2701
rect 2410 2698 2478 2701
rect 2634 2698 2662 2701
rect 2674 2698 2830 2701
rect 3098 2698 3126 2701
rect 3674 2698 3710 2701
rect 3714 2698 3830 2701
rect 3938 2698 3966 2701
rect 4130 2698 4142 2701
rect 4182 2698 4230 2701
rect 654 2692 657 2698
rect 1558 2692 1561 2698
rect 3198 2692 3201 2698
rect 146 2688 414 2691
rect 602 2688 654 2691
rect 882 2688 886 2691
rect 1186 2688 1214 2691
rect 1594 2688 1897 2691
rect 1978 2688 2030 2691
rect 2034 2688 2070 2691
rect 2114 2688 2118 2691
rect 2386 2688 2390 2691
rect 2482 2688 2486 2691
rect 2498 2688 2982 2691
rect 2986 2688 3038 2691
rect 3090 2688 3094 2691
rect 3346 2688 3390 2691
rect 3730 2688 3790 2691
rect 3810 2688 3982 2691
rect 4182 2691 4185 2698
rect 4042 2688 4185 2691
rect 14 2681 17 2688
rect 14 2678 142 2681
rect 582 2681 585 2688
rect 1894 2682 1897 2688
rect 582 2678 622 2681
rect 642 2678 646 2681
rect 682 2678 686 2681
rect 730 2678 814 2681
rect 842 2678 886 2681
rect 1658 2678 1702 2681
rect 1730 2678 1798 2681
rect 1994 2678 2102 2681
rect 2182 2681 2185 2688
rect 2454 2682 2457 2688
rect 2106 2678 2222 2681
rect 2250 2678 2286 2681
rect 2618 2678 2846 2681
rect 2882 2678 3030 2681
rect 3034 2678 3142 2681
rect 3186 2678 3278 2681
rect 3662 2681 3665 2688
rect 3662 2678 3678 2681
rect 3698 2678 3742 2681
rect 3798 2681 3801 2688
rect 3770 2678 3801 2681
rect 4002 2678 4022 2681
rect 4122 2678 4206 2681
rect 4274 2678 4286 2681
rect 4314 2678 4358 2681
rect -26 2671 -22 2672
rect -26 2668 22 2671
rect 50 2668 70 2671
rect 122 2668 222 2671
rect 562 2668 734 2671
rect 746 2668 766 2671
rect 794 2668 902 2671
rect 1338 2668 1481 2671
rect 1614 2671 1617 2678
rect 1578 2668 1617 2671
rect 1770 2668 1774 2671
rect 2242 2668 2286 2671
rect 2290 2668 2334 2671
rect 2606 2671 2609 2678
rect 2546 2668 2609 2671
rect 2890 2668 2902 2671
rect 3122 2668 3198 2671
rect 3402 2668 3406 2671
rect 3442 2668 3446 2671
rect 3474 2668 3534 2671
rect 3650 2668 3686 2671
rect 3738 2668 3785 2671
rect 3794 2668 3806 2671
rect 3898 2668 3902 2671
rect 3942 2671 3945 2678
rect 3906 2668 3945 2671
rect 3986 2668 4014 2671
rect 4042 2668 4046 2671
rect 4050 2668 4086 2671
rect 4090 2668 4246 2671
rect 4258 2668 4270 2671
rect 4338 2668 4374 2671
rect 4406 2671 4409 2678
rect 4378 2668 4409 2671
rect 82 2658 102 2661
rect 106 2658 134 2661
rect 186 2658 246 2661
rect 254 2661 257 2668
rect 254 2658 302 2661
rect 350 2661 353 2668
rect 350 2658 398 2661
rect 594 2658 702 2661
rect 730 2658 734 2661
rect 754 2658 758 2661
rect 834 2658 1022 2661
rect 1142 2661 1145 2668
rect 1382 2662 1385 2668
rect 1478 2662 1481 2668
rect 1142 2658 1222 2661
rect 1322 2658 1326 2661
rect 1622 2661 1625 2668
rect 1622 2658 1646 2661
rect 1694 2658 1702 2661
rect 1706 2658 1726 2661
rect 1830 2661 1833 2668
rect 1738 2658 1833 2661
rect 2182 2658 2190 2661
rect 2306 2658 2350 2661
rect 2550 2658 2566 2661
rect 2726 2661 2729 2668
rect 2706 2658 2729 2661
rect 2914 2658 2950 2661
rect 3098 2658 3150 2661
rect 3154 2658 3174 2661
rect 3266 2658 3273 2661
rect 3394 2658 3750 2661
rect 3782 2661 3785 2668
rect 3782 2658 3841 2661
rect 3930 2658 3958 2661
rect 4090 2658 4126 2661
rect 4210 2658 4214 2661
rect 4330 2658 4350 2661
rect 318 2652 321 2658
rect -26 2651 -22 2652
rect -26 2648 6 2651
rect 370 2648 542 2651
rect 602 2648 606 2651
rect 626 2648 646 2651
rect 650 2648 670 2651
rect 714 2648 718 2651
rect 734 2651 737 2658
rect 734 2648 766 2651
rect 1318 2651 1321 2658
rect 2182 2652 2185 2658
rect 2550 2652 2553 2658
rect 3270 2652 3273 2658
rect 3838 2652 3841 2658
rect 970 2648 1321 2651
rect 1370 2648 1398 2651
rect 1642 2648 1646 2651
rect 2258 2648 2262 2651
rect 2362 2648 2430 2651
rect 2586 2648 2670 2651
rect 2674 2648 2718 2651
rect 2722 2648 2822 2651
rect 2826 2648 2838 2651
rect 2850 2648 2918 2651
rect 2962 2648 3006 2651
rect 3210 2648 3214 2651
rect 3370 2648 3382 2651
rect 3386 2648 3398 2651
rect 3402 2648 3422 2651
rect 3426 2648 3446 2651
rect 3466 2648 3710 2651
rect 3746 2648 3774 2651
rect 3946 2648 3958 2651
rect 3962 2648 3966 2651
rect 4058 2648 4062 2651
rect 4170 2648 4206 2651
rect 4210 2648 4214 2651
rect 4306 2648 4318 2651
rect 4354 2648 4374 2651
rect 4378 2648 4398 2651
rect 4402 2648 4454 2651
rect 490 2638 566 2641
rect 570 2638 614 2641
rect 698 2638 750 2641
rect 1218 2638 1350 2641
rect 1354 2638 2934 2641
rect 2938 2638 3374 2641
rect 3402 2638 3622 2641
rect 4066 2638 4158 2641
rect 4174 2638 4182 2641
rect 4174 2632 4177 2638
rect 2050 2628 2230 2631
rect 2234 2628 2241 2631
rect 2306 2628 2310 2631
rect 2322 2628 2382 2631
rect 2386 2628 2766 2631
rect 2954 2628 2974 2631
rect 2994 2628 3150 2631
rect 3282 2628 3670 2631
rect 298 2618 366 2621
rect 490 2618 2078 2621
rect 2090 2618 2910 2621
rect 3226 2618 3638 2621
rect 3918 2621 3921 2628
rect 3890 2618 3958 2621
rect 546 2608 886 2611
rect 2114 2608 2350 2611
rect 2362 2608 2422 2611
rect 2426 2608 2518 2611
rect 2786 2608 3534 2611
rect 3634 2608 3646 2611
rect 496 2603 498 2607
rect 502 2603 505 2607
rect 510 2603 512 2607
rect 1022 2602 1025 2608
rect 1520 2603 1522 2607
rect 1526 2603 1529 2607
rect 1534 2603 1536 2607
rect 2544 2603 2546 2607
rect 2550 2603 2553 2607
rect 2558 2603 2560 2607
rect 3568 2603 3570 2607
rect 3574 2603 3577 2607
rect 3582 2603 3584 2607
rect 658 2598 798 2601
rect 1450 2598 1494 2601
rect 1786 2598 1846 2601
rect 2242 2598 2430 2601
rect 2570 2598 2958 2601
rect 3354 2598 3366 2601
rect 3698 2598 3902 2601
rect 3906 2598 4150 2601
rect 762 2588 1030 2591
rect 1466 2588 1502 2591
rect 1562 2588 1566 2591
rect 1802 2588 1806 2591
rect 2138 2588 2142 2591
rect 2146 2588 2318 2591
rect 2394 2588 2462 2591
rect 2546 2588 2614 2591
rect 2754 2588 3014 2591
rect 3322 2588 3350 2591
rect 1662 2582 1665 2588
rect 706 2578 790 2581
rect 794 2578 862 2581
rect 2194 2578 2750 2581
rect 2986 2578 3158 2581
rect 3162 2578 3310 2581
rect 3378 2578 3494 2581
rect 3602 2578 3622 2581
rect 3626 2578 3742 2581
rect 4042 2578 4286 2581
rect 386 2568 686 2571
rect 690 2568 710 2571
rect 1146 2568 1262 2571
rect 1546 2568 1598 2571
rect 1602 2568 1734 2571
rect 2218 2568 2238 2571
rect 2242 2568 2318 2571
rect 2458 2568 2678 2571
rect 2690 2568 2710 2571
rect 2758 2571 2761 2578
rect 2758 2568 2814 2571
rect 2826 2568 2854 2571
rect 2930 2568 2934 2571
rect 3010 2568 3022 2571
rect 3026 2568 3150 2571
rect 3154 2568 3206 2571
rect 3210 2568 3214 2571
rect 3338 2568 3382 2571
rect 3490 2568 3574 2571
rect 3834 2568 3910 2571
rect 3914 2568 3926 2571
rect 4050 2568 4102 2571
rect 4138 2568 4158 2571
rect 4234 2568 4302 2571
rect 4330 2568 4342 2571
rect 4434 2568 4438 2571
rect 2862 2562 2865 2568
rect -26 2561 -22 2562
rect -26 2558 6 2561
rect 50 2558 190 2561
rect 634 2558 638 2561
rect 690 2558 758 2561
rect 850 2558 926 2561
rect 1082 2558 1086 2561
rect 1970 2558 2054 2561
rect 2090 2558 2358 2561
rect 2434 2558 2462 2561
rect 2610 2558 2662 2561
rect 2666 2558 2801 2561
rect 2906 2558 3078 2561
rect 3290 2558 3302 2561
rect 3306 2558 3326 2561
rect 3462 2561 3465 2568
rect 3426 2558 3465 2561
rect 3474 2558 3534 2561
rect 3638 2561 3641 2568
rect 4230 2562 4233 2568
rect 3570 2558 3641 2561
rect 3650 2558 3654 2561
rect 3738 2558 3742 2561
rect 3754 2558 3758 2561
rect 3762 2558 3798 2561
rect 3826 2558 3942 2561
rect 3978 2558 4006 2561
rect 4082 2558 4134 2561
rect 4258 2558 4278 2561
rect 4306 2558 4310 2561
rect 4314 2558 4334 2561
rect 4346 2558 4406 2561
rect 4474 2558 4518 2561
rect 4522 2558 4534 2561
rect 2798 2552 2801 2558
rect 3198 2552 3201 2558
rect 58 2548 70 2551
rect 226 2548 462 2551
rect 514 2548 630 2551
rect 658 2548 718 2551
rect 722 2548 726 2551
rect 770 2548 838 2551
rect 874 2548 902 2551
rect 922 2548 1078 2551
rect 1102 2548 1150 2551
rect 1730 2548 1734 2551
rect 1890 2548 1910 2551
rect 1914 2548 1950 2551
rect 1954 2548 1982 2551
rect 1994 2548 2126 2551
rect 2130 2548 2310 2551
rect 2466 2548 2726 2551
rect 2746 2548 2793 2551
rect 2802 2548 2870 2551
rect 2874 2548 2910 2551
rect 3322 2548 3398 2551
rect 3418 2548 3550 2551
rect 3554 2548 4214 2551
rect 4218 2548 4238 2551
rect 4242 2548 4470 2551
rect 4546 2548 4550 2551
rect 286 2542 289 2548
rect 1102 2542 1105 2548
rect -26 2538 -22 2542
rect 26 2538 70 2541
rect 378 2538 401 2541
rect 426 2538 526 2541
rect 598 2538 694 2541
rect 794 2538 822 2541
rect 858 2538 918 2541
rect 922 2538 942 2541
rect 994 2538 1030 2541
rect 1210 2538 1270 2541
rect 1730 2538 1830 2541
rect 1946 2538 1966 2541
rect 1994 2538 1998 2541
rect 2002 2538 2126 2541
rect 2130 2538 2142 2541
rect 2318 2541 2321 2548
rect 2790 2542 2793 2548
rect 2318 2538 2438 2541
rect 2530 2538 2678 2541
rect 2682 2538 2782 2541
rect 2794 2538 2902 2541
rect 2910 2541 2913 2548
rect 2910 2538 2926 2541
rect 2966 2541 2969 2548
rect 2966 2538 2990 2541
rect 3250 2538 3262 2541
rect 3338 2538 3422 2541
rect 3434 2538 3438 2541
rect 3486 2538 3518 2541
rect 3522 2538 3558 2541
rect 3634 2538 3670 2541
rect 3730 2538 3846 2541
rect 3850 2538 3894 2541
rect 3914 2538 3926 2541
rect 3962 2538 3974 2541
rect 4066 2538 4142 2541
rect 4186 2538 4190 2541
rect 4274 2538 4318 2541
rect 4330 2538 4350 2541
rect 4354 2538 4438 2541
rect 4486 2541 4489 2548
rect 4486 2538 4518 2541
rect -26 2531 -23 2538
rect 398 2532 401 2538
rect 598 2532 601 2538
rect -26 2528 30 2531
rect 50 2528 142 2531
rect 474 2528 494 2531
rect 650 2528 686 2531
rect 822 2531 825 2538
rect 3486 2532 3489 2538
rect 822 2528 870 2531
rect 874 2528 894 2531
rect 898 2528 910 2531
rect 1634 2528 1838 2531
rect 1858 2528 1990 2531
rect 2562 2528 2654 2531
rect 2658 2528 2742 2531
rect 2754 2528 2830 2531
rect 2842 2528 2974 2531
rect 2978 2528 3318 2531
rect 3538 2528 3542 2531
rect 3546 2528 3558 2531
rect 3646 2528 3822 2531
rect 3922 2528 4086 2531
rect 4254 2531 4257 2538
rect 4202 2528 4257 2531
rect 4338 2528 4342 2531
rect 4386 2528 4398 2531
rect 4418 2528 4438 2531
rect 4442 2528 4446 2531
rect 266 2518 294 2521
rect 298 2518 470 2521
rect 482 2518 486 2521
rect 562 2518 742 2521
rect 842 2518 958 2521
rect 1122 2518 1294 2521
rect 1298 2518 2246 2521
rect 2362 2518 2366 2521
rect 2370 2518 2886 2521
rect 2962 2518 2966 2521
rect 3202 2518 3206 2521
rect 3430 2521 3433 2528
rect 3646 2522 3649 2528
rect 3430 2518 3622 2521
rect 3698 2518 3702 2521
rect 3722 2518 3902 2521
rect 3906 2518 3966 2521
rect 4182 2521 4185 2528
rect 4066 2518 4185 2521
rect 4194 2518 4558 2521
rect 450 2508 486 2511
rect 642 2508 742 2511
rect 1522 2508 1742 2511
rect 2130 2508 2294 2511
rect 2842 2508 2854 2511
rect 2938 2508 2958 2511
rect 3266 2508 3526 2511
rect 3530 2508 3734 2511
rect 3754 2508 3990 2511
rect 4194 2508 4254 2511
rect 4258 2508 4462 2511
rect 4466 2508 4494 2511
rect 4498 2508 4518 2511
rect 1000 2503 1002 2507
rect 1006 2503 1009 2507
rect 1014 2503 1016 2507
rect 2024 2503 2026 2507
rect 2030 2503 2033 2507
rect 2038 2503 2040 2507
rect 3048 2503 3050 2507
rect 3054 2503 3057 2507
rect 3062 2503 3064 2507
rect 4080 2503 4082 2507
rect 4086 2503 4089 2507
rect 4094 2503 4096 2507
rect 250 2498 358 2501
rect 586 2498 638 2501
rect 762 2498 993 2501
rect 1362 2498 1518 2501
rect 1666 2498 1670 2501
rect 2098 2498 2174 2501
rect 2178 2498 2206 2501
rect 2218 2498 2281 2501
rect 2290 2498 2390 2501
rect 2610 2498 2926 2501
rect 3074 2498 3078 2501
rect 3082 2498 3238 2501
rect 3258 2498 3350 2501
rect 3602 2498 3702 2501
rect 3706 2498 3782 2501
rect 4138 2498 4174 2501
rect 4186 2498 4278 2501
rect 4322 2498 4326 2501
rect 4330 2498 4390 2501
rect 758 2488 774 2491
rect 842 2488 862 2491
rect 890 2488 982 2491
rect 990 2491 993 2498
rect 1646 2492 1649 2498
rect 990 2488 1046 2491
rect 1458 2488 1462 2491
rect 1466 2488 1486 2491
rect 1986 2488 2022 2491
rect 2042 2488 2046 2491
rect 2250 2488 2270 2491
rect 2278 2491 2281 2498
rect 2278 2488 2350 2491
rect 2482 2488 2510 2491
rect 2514 2488 2918 2491
rect 3226 2488 3238 2491
rect 3274 2488 3294 2491
rect 3434 2488 3481 2491
rect 758 2482 761 2488
rect 74 2478 158 2481
rect 162 2478 270 2481
rect 274 2478 334 2481
rect 554 2478 566 2481
rect 802 2478 846 2481
rect 850 2478 878 2481
rect 882 2478 886 2481
rect 978 2478 1030 2481
rect 1034 2478 1038 2481
rect 1102 2481 1105 2488
rect 1102 2478 1142 2481
rect 1762 2478 1806 2481
rect 2522 2478 2526 2481
rect 2578 2478 2582 2481
rect 2594 2478 2598 2481
rect 2810 2478 2862 2481
rect 2926 2481 2929 2488
rect 3478 2482 3481 2488
rect 3690 2488 3694 2491
rect 3818 2488 3966 2491
rect 4038 2488 4086 2491
rect 4114 2488 4334 2491
rect 3486 2482 3489 2488
rect 2882 2478 2929 2481
rect 3102 2478 3110 2481
rect 3114 2478 3166 2481
rect 3186 2478 3342 2481
rect 3466 2478 3470 2481
rect 3558 2481 3561 2488
rect 4038 2482 4041 2488
rect 3514 2478 3561 2481
rect 3578 2478 3638 2481
rect 3642 2478 3782 2481
rect 3786 2478 3830 2481
rect 3834 2478 3838 2481
rect 3886 2478 3894 2481
rect 3898 2478 3934 2481
rect 3978 2478 4030 2481
rect 4170 2478 4198 2481
rect 4290 2478 4342 2481
rect 4370 2478 4430 2481
rect 4450 2478 4486 2481
rect 4582 2481 4585 2488
rect 4562 2478 4585 2481
rect 4590 2482 4593 2488
rect 918 2472 921 2478
rect 34 2468 54 2471
rect 482 2468 574 2471
rect 1010 2468 1014 2471
rect 1086 2471 1089 2478
rect 1086 2468 1110 2471
rect 1130 2468 1182 2471
rect 1202 2468 1294 2471
rect 1374 2471 1377 2478
rect 1470 2471 1473 2478
rect 1306 2468 1473 2471
rect 1874 2468 2078 2471
rect 2142 2471 2145 2478
rect 2758 2472 2761 2478
rect 2774 2472 2777 2478
rect 2142 2468 2174 2471
rect 2266 2468 2318 2471
rect 2338 2468 2454 2471
rect 2514 2468 2574 2471
rect 2578 2468 2630 2471
rect 2978 2468 2982 2471
rect 2990 2468 3062 2471
rect 3066 2468 3310 2471
rect 3438 2471 3441 2478
rect 3438 2468 3478 2471
rect 3482 2468 3526 2471
rect 3530 2468 3542 2471
rect 3586 2468 3590 2471
rect 3642 2468 3646 2471
rect 3650 2468 3686 2471
rect 3690 2468 3750 2471
rect 3758 2468 3790 2471
rect 3818 2468 3830 2471
rect 3986 2468 4046 2471
rect 4050 2468 4078 2471
rect 4082 2468 4118 2471
rect 4138 2468 4142 2471
rect 4146 2468 4174 2471
rect 4214 2468 4254 2471
rect 4362 2468 4382 2471
rect 4434 2468 4449 2471
rect 58 2458 62 2461
rect 206 2461 209 2468
rect 146 2458 209 2461
rect 330 2458 417 2461
rect 698 2458 702 2461
rect 726 2461 729 2468
rect 726 2458 774 2461
rect 878 2461 881 2468
rect 842 2458 881 2461
rect 926 2462 929 2468
rect 1074 2458 1118 2461
rect 1154 2458 1494 2461
rect 1514 2458 1534 2461
rect 1538 2458 1630 2461
rect 1678 2461 1681 2468
rect 1774 2461 1777 2468
rect 1634 2458 1777 2461
rect 1802 2459 1806 2461
rect 1798 2458 1806 2459
rect 2110 2461 2113 2468
rect 2502 2462 2505 2468
rect 2110 2458 2230 2461
rect 2234 2458 2254 2461
rect 2586 2458 2758 2461
rect 2790 2461 2793 2468
rect 2990 2462 2993 2468
rect 2790 2458 2857 2461
rect 2874 2458 2974 2461
rect 3122 2458 3126 2461
rect 3138 2458 3230 2461
rect 3338 2458 3358 2461
rect 3418 2458 3518 2461
rect 3522 2458 3606 2461
rect 3666 2458 3689 2461
rect 3758 2461 3761 2468
rect 4214 2462 4217 2468
rect 4446 2462 4449 2468
rect 3698 2458 3761 2461
rect 3770 2458 3806 2461
rect 3818 2458 3942 2461
rect 3958 2458 4070 2461
rect 4162 2458 4190 2461
rect 4234 2458 4246 2461
rect 4338 2458 4406 2461
rect 414 2452 417 2458
rect 1902 2452 1905 2458
rect 2390 2452 2393 2458
rect 2854 2452 2857 2458
rect -26 2451 -22 2452
rect -26 2448 6 2451
rect 34 2448 118 2451
rect 482 2448 518 2451
rect 522 2448 606 2451
rect 610 2448 614 2451
rect 658 2448 894 2451
rect 986 2448 1390 2451
rect 1546 2448 1686 2451
rect 2210 2448 2222 2451
rect 2226 2448 2249 2451
rect 2482 2448 2526 2451
rect 2530 2448 2598 2451
rect 2602 2448 2734 2451
rect 3178 2448 3206 2451
rect 3290 2448 3302 2451
rect 3306 2448 3326 2451
rect 3354 2448 3438 2451
rect 3650 2448 3654 2451
rect 3658 2448 3670 2451
rect 3686 2451 3689 2458
rect 3958 2452 3961 2458
rect 3686 2448 3710 2451
rect 3754 2448 3774 2451
rect 3798 2448 3846 2451
rect 3930 2448 3934 2451
rect 4346 2448 4366 2451
rect 4414 2451 4417 2458
rect 4414 2448 4454 2451
rect 4490 2448 4526 2451
rect 346 2438 510 2441
rect 514 2438 614 2441
rect 618 2438 630 2441
rect 894 2441 897 2448
rect 2246 2442 2249 2448
rect 3798 2442 3801 2448
rect 894 2438 1094 2441
rect 1154 2438 1254 2441
rect 1258 2438 1606 2441
rect 2278 2438 2422 2441
rect 2642 2438 3214 2441
rect 3330 2438 3414 2441
rect 3530 2438 3798 2441
rect 3858 2438 3974 2441
rect 3994 2438 4006 2441
rect 4290 2438 4374 2441
rect 282 2428 862 2431
rect 866 2428 1078 2431
rect 1130 2428 1406 2431
rect 1410 2428 1494 2431
rect 2278 2431 2281 2438
rect 1498 2428 2281 2431
rect 2286 2428 3182 2431
rect 3302 2431 3305 2438
rect 3302 2428 3494 2431
rect 3562 2428 3814 2431
rect 3842 2428 4494 2431
rect 862 2418 870 2421
rect 874 2418 974 2421
rect 1426 2418 1662 2421
rect 2286 2421 2289 2428
rect 1802 2418 2289 2421
rect 2322 2418 2566 2421
rect 2682 2418 2902 2421
rect 2922 2418 4358 2421
rect 4566 2421 4569 2428
rect 4370 2418 4569 2421
rect 1554 2408 1558 2411
rect 2098 2408 2342 2411
rect 2570 2408 2934 2411
rect 2946 2408 3230 2411
rect 3242 2408 3398 2411
rect 3594 2408 4006 2411
rect 4018 2408 4046 2411
rect 4074 2408 4318 2411
rect 4442 2408 4590 2411
rect 496 2403 498 2407
rect 502 2403 505 2407
rect 510 2403 512 2407
rect 1520 2403 1522 2407
rect 1526 2403 1529 2407
rect 1534 2403 1536 2407
rect 1662 2402 1665 2408
rect 2544 2403 2546 2407
rect 2550 2403 2553 2407
rect 2558 2403 2560 2407
rect 3568 2403 3570 2407
rect 3574 2403 3577 2407
rect 3582 2403 3584 2407
rect 986 2398 998 2401
rect 2202 2398 2302 2401
rect 2882 2398 2918 2401
rect 2954 2398 3246 2401
rect 3266 2398 3358 2401
rect 3826 2398 3910 2401
rect 4050 2398 4478 2401
rect 874 2388 1206 2391
rect 1234 2388 1358 2391
rect 1362 2388 2318 2391
rect 2346 2388 2414 2391
rect 2778 2388 2798 2391
rect 2810 2388 3190 2391
rect 3218 2388 3302 2391
rect 3306 2388 3350 2391
rect 3474 2388 3742 2391
rect 3754 2388 3918 2391
rect 4210 2388 4214 2391
rect 4482 2388 4526 2391
rect 46 2381 49 2388
rect 46 2378 94 2381
rect 98 2378 110 2381
rect 114 2378 190 2381
rect 194 2378 230 2381
rect 234 2378 262 2381
rect 266 2378 390 2381
rect 394 2378 406 2381
rect 970 2378 998 2381
rect 1618 2378 2454 2381
rect 2458 2378 2998 2381
rect 3178 2378 3366 2381
rect 3514 2378 3550 2381
rect 3630 2378 3638 2381
rect 3642 2378 3670 2381
rect 3882 2378 3926 2381
rect 4034 2378 4062 2381
rect 4066 2378 4430 2381
rect 178 2368 582 2371
rect 722 2368 934 2371
rect 990 2368 1158 2371
rect 1330 2368 1374 2371
rect 1378 2368 1798 2371
rect 1898 2368 1950 2371
rect 2762 2368 2870 2371
rect 2874 2368 3262 2371
rect 3266 2368 3366 2371
rect 3378 2368 4118 2371
rect 4210 2368 4214 2371
rect 4242 2368 4278 2371
rect 4346 2368 4350 2371
rect 4410 2368 4502 2371
rect 4518 2371 4521 2378
rect 4514 2368 4521 2371
rect 4542 2371 4545 2378
rect 4538 2368 4545 2371
rect 990 2362 993 2368
rect -26 2361 -22 2362
rect -26 2358 22 2361
rect 146 2358 190 2361
rect 194 2358 206 2361
rect 210 2358 342 2361
rect 730 2358 918 2361
rect 1002 2358 1014 2361
rect 1018 2358 1062 2361
rect 1226 2358 1254 2361
rect 1410 2358 1414 2361
rect 1658 2358 1702 2361
rect 1978 2358 2174 2361
rect 2246 2361 2249 2368
rect 2246 2358 2278 2361
rect 2314 2358 2334 2361
rect 2374 2361 2377 2368
rect 4406 2362 4409 2368
rect 2338 2358 2406 2361
rect 2410 2358 2478 2361
rect 2706 2358 2806 2361
rect 2854 2358 2862 2361
rect 2866 2358 2902 2361
rect 2922 2358 2961 2361
rect 162 2348 273 2351
rect 330 2348 574 2351
rect 578 2348 646 2351
rect 690 2348 710 2351
rect 746 2348 894 2351
rect 954 2348 1262 2351
rect 1382 2348 1446 2351
rect 1918 2351 1921 2358
rect 1918 2348 1998 2351
rect -26 2341 -22 2342
rect -26 2338 6 2341
rect 30 2341 33 2348
rect 270 2342 273 2348
rect 926 2342 929 2348
rect 1382 2342 1385 2348
rect 2074 2348 2118 2351
rect 2174 2351 2177 2358
rect 2582 2352 2585 2358
rect 2814 2352 2817 2358
rect 2958 2352 2961 2358
rect 3018 2358 3054 2361
rect 3198 2358 3206 2361
rect 3210 2358 3230 2361
rect 3234 2358 3310 2361
rect 3354 2358 3542 2361
rect 3602 2358 3630 2361
rect 3690 2358 3710 2361
rect 3714 2358 3750 2361
rect 3810 2358 3833 2361
rect 3850 2358 3870 2361
rect 3922 2358 3950 2361
rect 3970 2358 3998 2361
rect 4146 2358 4150 2361
rect 4194 2358 4273 2361
rect 4338 2358 4366 2361
rect 4474 2358 4542 2361
rect 2974 2352 2977 2358
rect 3830 2352 3833 2358
rect 3998 2352 4001 2358
rect 4270 2352 4273 2358
rect 2138 2348 2222 2351
rect 2234 2348 2254 2351
rect 2266 2348 2278 2351
rect 2282 2348 2446 2351
rect 2602 2348 2654 2351
rect 2714 2348 2758 2351
rect 2762 2348 2782 2351
rect 2834 2348 2838 2351
rect 2906 2348 2926 2351
rect 2986 2348 3094 2351
rect 3098 2348 3134 2351
rect 3138 2348 3262 2351
rect 3266 2348 3350 2351
rect 3402 2348 3406 2351
rect 3458 2348 3486 2351
rect 3490 2348 3518 2351
rect 3554 2348 3590 2351
rect 3626 2348 3646 2351
rect 3706 2348 3814 2351
rect 3858 2348 3862 2351
rect 3946 2348 3974 2351
rect 4018 2348 4022 2351
rect 4218 2348 4222 2351
rect 4274 2348 4278 2351
rect 4330 2348 4366 2351
rect 4370 2348 4422 2351
rect 4498 2348 4510 2351
rect 4582 2351 4585 2358
rect 4578 2348 4585 2351
rect 30 2338 206 2341
rect 586 2338 678 2341
rect 746 2338 798 2341
rect 1018 2338 1062 2341
rect 1098 2338 1142 2341
rect 1194 2338 1262 2341
rect 1282 2338 1358 2341
rect 1650 2338 1694 2341
rect 1698 2338 1790 2341
rect 2130 2338 2150 2341
rect 2202 2338 2206 2341
rect 2394 2338 2422 2341
rect 2458 2338 2486 2341
rect 2530 2338 2718 2341
rect 2738 2338 2742 2341
rect 2762 2338 3006 2341
rect 3042 2338 3070 2341
rect 3114 2338 3158 2341
rect 3242 2338 3270 2341
rect 3306 2338 3321 2341
rect 14 2331 17 2338
rect 14 2328 150 2331
rect 178 2328 206 2331
rect 678 2331 681 2338
rect 2918 2332 2921 2338
rect 3318 2332 3321 2338
rect 3402 2338 3414 2341
rect 3434 2338 3438 2341
rect 3602 2338 3606 2341
rect 3658 2338 3726 2341
rect 3770 2338 3782 2341
rect 3786 2338 3862 2341
rect 3970 2338 3974 2341
rect 3978 2338 4006 2341
rect 4150 2341 4153 2348
rect 4018 2338 4153 2341
rect 4178 2338 4406 2341
rect 4410 2338 4574 2341
rect 3366 2332 3369 2338
rect 4158 2332 4161 2338
rect 678 2328 814 2331
rect 818 2328 862 2331
rect 878 2328 894 2331
rect 954 2328 958 2331
rect 1730 2328 1950 2331
rect 1954 2328 2174 2331
rect 2298 2328 2302 2331
rect 2362 2328 2366 2331
rect 2466 2328 2470 2331
rect 2646 2328 2654 2331
rect 2658 2328 2902 2331
rect 3010 2328 3094 2331
rect 3098 2328 3118 2331
rect 3122 2328 3206 2331
rect 3210 2328 3270 2331
rect 3378 2328 3430 2331
rect 3458 2328 3502 2331
rect 3562 2328 3590 2331
rect 3594 2328 3686 2331
rect 3746 2328 3790 2331
rect 3866 2328 3918 2331
rect 4130 2328 4158 2331
rect 4170 2328 4246 2331
rect 4250 2328 4262 2331
rect 4314 2328 4318 2331
rect 4346 2328 4430 2331
rect 4466 2328 4478 2331
rect 4482 2328 4534 2331
rect 4562 2328 4566 2331
rect 214 2318 222 2321
rect 226 2318 398 2321
rect 454 2321 457 2328
rect 878 2322 881 2328
rect 454 2318 510 2321
rect 942 2321 945 2328
rect 942 2318 974 2321
rect 986 2318 1078 2321
rect 1754 2318 1758 2321
rect 1922 2318 2182 2321
rect 2618 2318 2718 2321
rect 2842 2318 2950 2321
rect 2954 2318 2982 2321
rect 3002 2318 3254 2321
rect 3258 2318 3406 2321
rect 3626 2318 3694 2321
rect 3786 2318 4086 2321
rect 4194 2318 4254 2321
rect 4258 2318 4382 2321
rect 4402 2318 4470 2321
rect 4546 2318 4558 2321
rect 122 2308 214 2311
rect 218 2308 318 2311
rect 322 2308 454 2311
rect 458 2308 830 2311
rect 834 2308 902 2311
rect 1210 2308 1438 2311
rect 2170 2308 2246 2311
rect 2410 2308 2742 2311
rect 2770 2308 2814 2311
rect 3082 2308 3150 2311
rect 3154 2308 3214 2311
rect 3306 2308 3534 2311
rect 3690 2308 3774 2311
rect 3778 2308 3870 2311
rect 4210 2308 4246 2311
rect 4250 2308 4302 2311
rect 4314 2308 4326 2311
rect 4378 2308 4382 2311
rect 1000 2303 1002 2307
rect 1006 2303 1009 2307
rect 1014 2303 1016 2307
rect 2024 2303 2026 2307
rect 2030 2303 2033 2307
rect 2038 2303 2040 2307
rect 3048 2303 3050 2307
rect 3054 2303 3057 2307
rect 3062 2303 3064 2307
rect 4080 2303 4082 2307
rect 4086 2303 4089 2307
rect 4094 2303 4096 2307
rect 514 2298 886 2301
rect 1370 2298 1374 2301
rect 1442 2298 1486 2301
rect 1490 2298 1574 2301
rect 1578 2298 1590 2301
rect 1826 2298 1846 2301
rect 2050 2298 2158 2301
rect 2202 2298 2350 2301
rect 2538 2298 2630 2301
rect 2682 2298 2686 2301
rect 2690 2298 2734 2301
rect 2778 2298 2854 2301
rect 2866 2298 2990 2301
rect 3122 2298 3174 2301
rect 3250 2298 3382 2301
rect 3410 2298 3601 2301
rect 3642 2298 3702 2301
rect 3706 2298 3798 2301
rect 3842 2298 3910 2301
rect 4258 2298 4494 2301
rect 4522 2298 4574 2301
rect 302 2291 305 2298
rect 302 2288 310 2291
rect 338 2288 358 2291
rect 958 2288 966 2291
rect 970 2288 1078 2291
rect 1354 2288 1470 2291
rect 1650 2288 1886 2291
rect 1890 2288 2238 2291
rect 2266 2288 2270 2291
rect 2330 2288 2398 2291
rect 2522 2288 2566 2291
rect 2634 2288 2678 2291
rect 2690 2288 2726 2291
rect 2730 2288 3510 2291
rect 3514 2288 3550 2291
rect 3554 2288 3590 2291
rect 3598 2291 3601 2298
rect 3598 2288 3822 2291
rect 4130 2288 4294 2291
rect 4298 2288 4390 2291
rect 4474 2288 4486 2291
rect 1086 2282 1089 2288
rect 1102 2282 1105 2288
rect 234 2278 238 2281
rect 306 2278 350 2281
rect 650 2278 798 2281
rect 894 2278 958 2281
rect 978 2278 990 2281
rect 1034 2278 1038 2281
rect 1322 2278 1382 2281
rect 1554 2278 1670 2281
rect 1674 2278 1886 2281
rect 1890 2278 1982 2281
rect 2218 2278 2574 2281
rect 2754 2278 2758 2281
rect 2778 2278 2782 2281
rect 2786 2278 2814 2281
rect 2886 2278 2894 2281
rect 2898 2278 2926 2281
rect 3002 2278 3030 2281
rect 3154 2278 3206 2281
rect 3226 2278 3238 2281
rect 3274 2278 3310 2281
rect 3434 2278 3438 2281
rect 3586 2278 3646 2281
rect 3650 2278 3670 2281
rect 3674 2278 3678 2281
rect 3730 2278 3753 2281
rect -26 2271 -22 2272
rect -26 2268 126 2271
rect 154 2268 174 2271
rect 330 2268 342 2271
rect 350 2271 353 2278
rect 470 2272 473 2278
rect 894 2272 897 2278
rect 350 2268 470 2271
rect 714 2268 734 2271
rect 778 2268 878 2271
rect 930 2268 1022 2271
rect 1082 2268 1398 2271
rect 1578 2268 1582 2271
rect 1922 2268 1926 2271
rect 2158 2271 2161 2278
rect 2158 2268 2182 2271
rect 2206 2271 2209 2278
rect 3494 2272 3497 2278
rect 3750 2272 3753 2278
rect 3810 2278 3825 2281
rect 3866 2278 3870 2281
rect 3874 2278 3894 2281
rect 3914 2278 3966 2281
rect 3986 2278 3998 2281
rect 4070 2278 4166 2281
rect 4262 2278 4302 2281
rect 4470 2281 4473 2288
rect 4386 2278 4473 2281
rect 3758 2272 3761 2278
rect 2206 2268 2262 2271
rect 2282 2268 2334 2271
rect 2338 2268 2358 2271
rect 2386 2268 2390 2271
rect 2666 2268 2670 2271
rect 2698 2268 2710 2271
rect 2714 2268 3006 2271
rect 3010 2268 3062 2271
rect 3066 2268 3094 2271
rect 3170 2268 3174 2271
rect 3178 2268 3190 2271
rect 3290 2268 3334 2271
rect 3370 2268 3494 2271
rect 3538 2268 3598 2271
rect 3794 2268 3814 2271
rect 3822 2271 3825 2278
rect 3822 2268 3910 2271
rect 3946 2268 3974 2271
rect 4070 2271 4073 2278
rect 4262 2272 4265 2278
rect 4010 2268 4073 2271
rect 4090 2268 4094 2271
rect 4118 2268 4134 2271
rect 4346 2268 4409 2271
rect 4450 2268 4454 2271
rect 170 2258 233 2261
rect 386 2258 545 2261
rect 730 2258 793 2261
rect 1074 2258 1137 2261
rect 1242 2258 1598 2261
rect 1610 2258 2326 2261
rect 2502 2261 2505 2268
rect 2502 2258 2566 2261
rect 2602 2258 2630 2261
rect 2642 2258 2734 2261
rect 2738 2258 2838 2261
rect 2882 2258 2889 2261
rect 2898 2258 2918 2261
rect 2938 2258 2942 2261
rect 2962 2258 2974 2261
rect 3106 2258 3118 2261
rect 3142 2261 3145 2268
rect 4118 2262 4121 2268
rect 4326 2262 4329 2268
rect 4406 2262 4409 2268
rect 3142 2258 3182 2261
rect 3226 2258 3326 2261
rect 3426 2258 3446 2261
rect 3474 2258 3478 2261
rect 3554 2258 3662 2261
rect 3666 2258 3686 2261
rect 3746 2258 3798 2261
rect 3826 2258 3846 2261
rect 4050 2258 4086 2261
rect 4138 2258 4174 2261
rect 4178 2258 4190 2261
rect 4202 2258 4270 2261
rect 4306 2258 4310 2261
rect 4378 2258 4393 2261
rect 4450 2258 4494 2261
rect 230 2252 233 2258
rect 542 2252 545 2258
rect 790 2252 793 2258
rect 1134 2252 1137 2258
rect 2894 2252 2897 2258
rect 4390 2252 4393 2258
rect 4526 2252 4529 2258
rect -26 2251 -22 2252
rect -26 2248 6 2251
rect 690 2248 774 2251
rect 2018 2248 2022 2251
rect 2186 2248 2230 2251
rect 2250 2248 2313 2251
rect 2402 2248 2566 2251
rect 2578 2248 2606 2251
rect 2610 2248 2614 2251
rect 2690 2248 2710 2251
rect 2714 2248 2774 2251
rect 2794 2248 2878 2251
rect 2906 2248 3022 2251
rect 3026 2248 3046 2251
rect 3050 2248 3110 2251
rect 3114 2248 3118 2251
rect 3138 2248 3158 2251
rect 3178 2248 3262 2251
rect 3346 2248 3374 2251
rect 3402 2248 3430 2251
rect 3538 2248 3558 2251
rect 3610 2248 3622 2251
rect 3626 2248 3654 2251
rect 3898 2248 3942 2251
rect 4050 2248 4070 2251
rect 4098 2248 4118 2251
rect 4178 2248 4254 2251
rect 4258 2248 4334 2251
rect 4346 2248 4350 2251
rect 2310 2242 2313 2248
rect 546 2238 734 2241
rect 738 2238 910 2241
rect 914 2238 950 2241
rect 954 2238 998 2241
rect 1002 2238 1038 2241
rect 1210 2238 2262 2241
rect 2330 2238 2758 2241
rect 2810 2238 2862 2241
rect 2890 2238 2942 2241
rect 2958 2238 2966 2241
rect 2970 2238 3222 2241
rect 3234 2238 3294 2241
rect 3362 2238 3422 2241
rect 3434 2238 3446 2241
rect 3482 2238 3750 2241
rect 4014 2241 4017 2248
rect 3954 2238 4062 2241
rect 4066 2238 4126 2241
rect 4154 2238 4198 2241
rect 4218 2238 4225 2241
rect 4330 2238 4486 2241
rect 4506 2238 4526 2241
rect 4566 2241 4569 2248
rect 4546 2238 4569 2241
rect 4222 2232 4225 2238
rect 4494 2232 4497 2238
rect -26 2231 -22 2232
rect -26 2228 78 2231
rect 306 2228 470 2231
rect 474 2228 534 2231
rect 538 2228 966 2231
rect 1282 2228 1478 2231
rect 1866 2228 2158 2231
rect 2162 2228 2414 2231
rect 2434 2228 2478 2231
rect 2482 2228 2606 2231
rect 2658 2228 2750 2231
rect 2762 2228 2806 2231
rect 2842 2228 3286 2231
rect 3386 2228 3822 2231
rect 3842 2228 4022 2231
rect 4034 2228 4190 2231
rect 4290 2228 4345 2231
rect 4342 2222 4345 2228
rect 938 2218 1422 2221
rect 1474 2218 2350 2221
rect 2514 2218 2910 2221
rect 3186 2218 3302 2221
rect 3394 2218 3638 2221
rect 3994 2218 4030 2221
rect 4130 2218 4158 2221
rect 4442 2218 4574 2221
rect -26 2211 -22 2212
rect -26 2208 54 2211
rect 762 2208 1302 2211
rect 1610 2208 2534 2211
rect 2610 2208 2630 2211
rect 2634 2208 2654 2211
rect 2762 2208 3390 2211
rect 3874 2208 4078 2211
rect 4090 2208 4134 2211
rect 4298 2208 4350 2211
rect 4434 2208 4478 2211
rect 496 2203 498 2207
rect 502 2203 505 2207
rect 510 2203 512 2207
rect 1520 2203 1522 2207
rect 1526 2203 1529 2207
rect 1534 2203 1536 2207
rect 2544 2203 2546 2207
rect 2550 2203 2553 2207
rect 2558 2203 2560 2207
rect 3568 2203 3570 2207
rect 3574 2203 3577 2207
rect 3582 2203 3584 2207
rect 590 2198 1062 2201
rect 1706 2198 1998 2201
rect 2002 2198 2310 2201
rect 2570 2198 3038 2201
rect 3234 2198 3462 2201
rect 3714 2198 4014 2201
rect 4026 2198 4094 2201
rect 4458 2198 4478 2201
rect -26 2191 -22 2192
rect -26 2188 38 2191
rect 98 2188 334 2191
rect 590 2191 593 2198
rect 1078 2192 1081 2198
rect 338 2188 593 2191
rect 602 2188 678 2191
rect 1138 2188 1622 2191
rect 1626 2188 2214 2191
rect 2434 2188 2438 2191
rect 2442 2188 2542 2191
rect 2682 2188 2910 2191
rect 3266 2188 3270 2191
rect 3398 2188 3593 2191
rect 3986 2188 4134 2191
rect 4330 2188 4334 2191
rect 26 2178 318 2181
rect 522 2178 606 2181
rect 826 2178 854 2181
rect 970 2178 1286 2181
rect 1290 2178 1310 2181
rect 1330 2178 1777 2181
rect 1858 2178 2102 2181
rect 2106 2178 2190 2181
rect 2226 2178 2230 2181
rect 2234 2178 2246 2181
rect 2250 2178 2254 2181
rect 2258 2178 2366 2181
rect 2918 2181 2921 2188
rect 2402 2178 2921 2181
rect 3010 2178 3062 2181
rect 3066 2178 3113 2181
rect 3134 2181 3137 2188
rect 3122 2178 3137 2181
rect 3146 2178 3302 2181
rect 3306 2178 3350 2181
rect 3398 2181 3401 2188
rect 3590 2182 3593 2188
rect 3354 2178 3401 2181
rect 3458 2178 3486 2181
rect 3498 2178 3518 2181
rect 3594 2178 3782 2181
rect 4058 2178 4134 2181
rect 4146 2178 4182 2181
rect 4290 2178 4374 2181
rect -26 2171 -22 2172
rect 6 2171 9 2178
rect 1774 2172 1777 2178
rect -26 2168 9 2171
rect 74 2168 110 2171
rect 202 2168 366 2171
rect 370 2168 430 2171
rect 434 2168 478 2171
rect 578 2168 1246 2171
rect 1322 2168 1422 2171
rect 1434 2168 1686 2171
rect 2114 2168 3078 2171
rect 3110 2171 3113 2178
rect 3110 2168 3150 2171
rect 3250 2168 3270 2171
rect 3274 2168 3382 2171
rect 3442 2168 3502 2171
rect 3666 2168 3750 2171
rect 4254 2171 4257 2178
rect 3978 2168 4257 2171
rect 4346 2168 4358 2171
rect 4362 2168 4430 2171
rect 3438 2162 3441 2168
rect 122 2158 238 2161
rect 242 2158 310 2161
rect 386 2158 566 2161
rect 794 2158 870 2161
rect 882 2158 1134 2161
rect 1154 2158 1158 2161
rect 1186 2158 1214 2161
rect 1218 2158 1345 2161
rect 1410 2158 1414 2161
rect 1434 2158 1438 2161
rect 1474 2158 1502 2161
rect 1506 2158 1726 2161
rect 2274 2158 2310 2161
rect 2314 2158 2321 2161
rect 2378 2158 2422 2161
rect 2426 2158 2441 2161
rect 2458 2158 2582 2161
rect 2658 2158 2662 2161
rect 2674 2158 2686 2161
rect 2738 2158 2782 2161
rect 2786 2158 2806 2161
rect 2810 2158 2838 2161
rect 2930 2158 3038 2161
rect 3042 2158 3358 2161
rect 3490 2158 3510 2161
rect 3598 2161 3601 2168
rect 3766 2162 3769 2168
rect 3522 2158 3601 2161
rect 3626 2158 3686 2161
rect 3706 2158 3710 2161
rect 3790 2161 3793 2168
rect 3786 2158 3793 2161
rect 3818 2158 3830 2161
rect 4050 2158 4206 2161
rect 4210 2158 4510 2161
rect -26 2151 -22 2152
rect -26 2148 110 2151
rect 182 2148 294 2151
rect 450 2148 454 2151
rect 466 2148 790 2151
rect 810 2148 841 2151
rect 182 2142 185 2148
rect 318 2141 321 2148
rect 422 2141 425 2148
rect 838 2142 841 2148
rect 882 2148 902 2151
rect 1114 2148 1142 2151
rect 1146 2148 1326 2151
rect 1342 2151 1345 2158
rect 1342 2148 1689 2151
rect 1698 2148 1742 2151
rect 1746 2148 1774 2151
rect 1854 2151 1857 2158
rect 1854 2148 1934 2151
rect 2214 2151 2217 2158
rect 2438 2152 2441 2158
rect 2210 2148 2217 2151
rect 2234 2148 2286 2151
rect 2314 2148 2326 2151
rect 2346 2148 2350 2151
rect 2354 2148 2398 2151
rect 2598 2151 2601 2158
rect 4046 2152 4049 2158
rect 2598 2148 2606 2151
rect 2682 2148 2686 2151
rect 2798 2148 2838 2151
rect 2946 2148 3006 2151
rect 3026 2148 3030 2151
rect 3042 2148 3134 2151
rect 3226 2148 3230 2151
rect 3362 2148 3382 2151
rect 3402 2148 3406 2151
rect 3422 2148 3454 2151
rect 3562 2148 3606 2151
rect 3730 2148 3758 2151
rect 3794 2148 3798 2151
rect 3802 2148 3822 2151
rect 3834 2148 3862 2151
rect 3866 2148 3894 2151
rect 3930 2148 3998 2151
rect 4066 2148 4078 2151
rect 4122 2148 4126 2151
rect 4162 2148 4182 2151
rect 4210 2148 4230 2151
rect 4266 2148 4294 2151
rect 4306 2148 4310 2151
rect 4434 2148 4438 2151
rect 4454 2148 4470 2151
rect 4506 2148 4590 2151
rect 846 2142 849 2148
rect 318 2138 425 2141
rect 514 2138 726 2141
rect 1086 2141 1089 2148
rect 1334 2142 1337 2148
rect 1686 2142 1689 2148
rect 2454 2142 2457 2148
rect 2462 2142 2465 2148
rect 2798 2142 2801 2148
rect 3182 2142 3185 2148
rect 3422 2142 3425 2148
rect 1086 2138 1134 2141
rect 1202 2138 1222 2141
rect 1450 2138 1454 2141
rect 1514 2138 1670 2141
rect 1698 2138 1702 2141
rect 1730 2138 1734 2141
rect 1778 2138 1782 2141
rect 2202 2138 2206 2141
rect 2250 2138 2270 2141
rect 2290 2138 2318 2141
rect 2322 2138 2406 2141
rect 2642 2138 2654 2141
rect 2658 2138 2678 2141
rect 2682 2138 2710 2141
rect 2914 2138 2998 2141
rect 3002 2138 3030 2141
rect 3034 2138 3078 2141
rect 3082 2138 3166 2141
rect 3218 2138 3222 2141
rect 3250 2138 3257 2141
rect 3274 2138 3278 2141
rect 3322 2138 3406 2141
rect 3494 2141 3497 2148
rect 3542 2141 3545 2148
rect 3494 2138 3545 2141
rect 3554 2138 3646 2141
rect 3674 2138 3750 2141
rect 3754 2138 3782 2141
rect 3786 2138 3814 2141
rect 3858 2138 3934 2141
rect 4034 2138 4054 2141
rect 4074 2138 4110 2141
rect 4130 2138 4166 2141
rect 4186 2138 4214 2141
rect 4230 2141 4233 2148
rect 4230 2138 4270 2141
rect 4278 2138 4286 2141
rect 4318 2141 4321 2148
rect 4454 2142 4457 2148
rect 4290 2138 4350 2141
rect 4386 2138 4430 2141
rect 4498 2138 4502 2141
rect 102 2131 105 2138
rect 102 2128 534 2131
rect 682 2128 686 2131
rect 754 2128 830 2131
rect 834 2128 910 2131
rect 914 2128 974 2131
rect 978 2128 990 2131
rect 1098 2128 1110 2131
rect 1162 2128 1206 2131
rect 1466 2128 1494 2131
rect 1682 2128 1718 2131
rect 1722 2128 1758 2131
rect 1998 2131 2001 2138
rect 3254 2132 3257 2138
rect 3782 2132 3785 2138
rect 1986 2128 2238 2131
rect 2282 2128 2366 2131
rect 2370 2128 2478 2131
rect 2546 2128 2782 2131
rect 2786 2128 2798 2131
rect 2802 2128 2822 2131
rect 2826 2128 2838 2131
rect 2946 2128 2974 2131
rect 2982 2128 3094 2131
rect 3106 2128 3110 2131
rect 3122 2128 3158 2131
rect 3170 2128 3174 2131
rect 3274 2128 3334 2131
rect 3514 2128 3550 2131
rect 3554 2128 3558 2131
rect 3674 2128 3678 2131
rect 3682 2128 3734 2131
rect 3850 2128 3862 2131
rect 3906 2128 3910 2131
rect 4170 2128 4182 2131
rect 4186 2128 4198 2131
rect 4214 2131 4217 2138
rect 4214 2128 4326 2131
rect 4434 2128 4478 2131
rect 4482 2128 4486 2131
rect 314 2118 326 2121
rect 1398 2121 1401 2128
rect 2982 2122 2985 2128
rect 3646 2122 3649 2128
rect 330 2118 1225 2121
rect 1398 2118 1689 2121
rect 1698 2118 1710 2121
rect 2018 2118 2046 2121
rect 2234 2118 2302 2121
rect 2330 2118 2382 2121
rect 2450 2118 2758 2121
rect 2770 2118 2782 2121
rect 3042 2118 3086 2121
rect 3106 2118 3118 2121
rect 3322 2118 3366 2121
rect 3434 2118 3502 2121
rect 3522 2118 3550 2121
rect 3658 2118 3702 2121
rect 3770 2118 3838 2121
rect 3966 2121 3969 2128
rect 4398 2122 4401 2128
rect 3858 2118 3969 2121
rect 4066 2118 4134 2121
rect 4258 2118 4262 2121
rect 4298 2118 4350 2121
rect 4410 2118 4438 2121
rect 4450 2118 4454 2121
rect 4458 2118 4462 2121
rect 4466 2118 4550 2121
rect 690 2108 974 2111
rect 1222 2111 1225 2118
rect 1222 2108 1438 2111
rect 1686 2111 1689 2118
rect 1686 2108 1750 2111
rect 1754 2108 2014 2111
rect 2538 2108 2878 2111
rect 2882 2108 2894 2111
rect 3138 2108 3254 2111
rect 3330 2108 3374 2111
rect 3378 2108 3494 2111
rect 3634 2108 3694 2111
rect 3874 2108 3878 2111
rect 4258 2108 4310 2111
rect 1000 2103 1002 2107
rect 1006 2103 1009 2107
rect 1014 2103 1016 2107
rect 2024 2103 2026 2107
rect 2030 2103 2033 2107
rect 2038 2103 2040 2107
rect 3048 2103 3050 2107
rect 3054 2103 3057 2107
rect 3062 2103 3064 2107
rect 4080 2103 4082 2107
rect 4086 2103 4089 2107
rect 4094 2103 4096 2107
rect 394 2098 454 2101
rect 458 2098 542 2101
rect 562 2098 662 2101
rect 666 2098 750 2101
rect 778 2098 990 2101
rect 1386 2098 1406 2101
rect 1522 2098 1542 2101
rect 1714 2098 1742 2101
rect 2234 2098 2406 2101
rect 2586 2098 2742 2101
rect 2762 2098 2934 2101
rect 2938 2098 2958 2101
rect 3098 2098 3153 2101
rect 3162 2098 3206 2101
rect 3218 2098 3238 2101
rect 3402 2098 3814 2101
rect 3866 2098 3974 2101
rect 3978 2098 3990 2101
rect 4010 2098 4070 2101
rect 4194 2098 4222 2101
rect 4226 2098 4486 2101
rect -26 2091 -22 2092
rect -26 2088 265 2091
rect 314 2088 334 2091
rect 338 2088 342 2091
rect 346 2088 470 2091
rect 802 2088 846 2091
rect 922 2088 966 2091
rect 986 2088 1070 2091
rect 1362 2088 1406 2091
rect 1466 2088 1510 2091
rect 1514 2088 1625 2091
rect 1658 2088 1766 2091
rect 1846 2088 1854 2091
rect 1858 2088 2270 2091
rect 2298 2088 2350 2091
rect 2354 2088 2390 2091
rect 2394 2088 2462 2091
rect 2486 2088 2494 2091
rect 2498 2088 2662 2091
rect 2682 2088 2737 2091
rect 2866 2088 2950 2091
rect 2958 2091 2961 2098
rect 2958 2088 3046 2091
rect 3106 2088 3134 2091
rect 3150 2091 3153 2098
rect 3150 2088 3214 2091
rect 3274 2088 3278 2091
rect 3386 2088 3438 2091
rect 3498 2088 3622 2091
rect 3714 2088 3782 2091
rect 3818 2088 4158 2091
rect 4162 2088 4262 2091
rect 4538 2088 4598 2091
rect 262 2082 265 2088
rect 782 2082 785 2088
rect 1078 2082 1081 2088
rect 1622 2082 1625 2088
rect 2734 2082 2737 2088
rect 266 2078 286 2081
rect 314 2078 438 2081
rect 594 2078 694 2081
rect 970 2078 1006 2081
rect 1018 2078 1054 2081
rect 1058 2078 1070 2081
rect 1098 2078 1102 2081
rect 1226 2078 1230 2081
rect 1234 2078 1294 2081
rect 1298 2078 1422 2081
rect 1578 2078 1598 2081
rect 1602 2078 1606 2081
rect 1674 2078 1734 2081
rect 1794 2078 1886 2081
rect 1922 2078 1966 2081
rect 1982 2078 1990 2081
rect 1994 2078 2166 2081
rect 2226 2078 2246 2081
rect 2346 2078 2606 2081
rect 2706 2078 2710 2081
rect 2874 2078 2934 2081
rect 2938 2078 2942 2081
rect 2954 2078 3366 2081
rect 3370 2078 3542 2081
rect 3642 2078 3678 2081
rect 3682 2078 3686 2081
rect 3690 2078 3822 2081
rect 3850 2078 3870 2081
rect 3898 2078 3958 2081
rect 4002 2078 4014 2081
rect 4042 2078 4190 2081
rect 4258 2078 4262 2081
rect 4314 2078 4350 2081
rect 4354 2078 4374 2081
rect 4430 2081 4433 2088
rect 4386 2078 4433 2081
rect 4490 2078 4510 2081
rect -26 2071 -22 2072
rect 30 2071 33 2078
rect -26 2068 33 2071
rect 282 2068 286 2071
rect 330 2068 398 2071
rect 406 2068 670 2071
rect 818 2068 838 2071
rect 866 2068 886 2071
rect 890 2068 894 2071
rect 910 2071 913 2078
rect 4270 2072 4273 2078
rect 910 2068 1038 2071
rect 1042 2068 1174 2071
rect 1210 2068 1246 2071
rect 1354 2068 1366 2071
rect 1386 2068 1406 2071
rect 1570 2068 1689 2071
rect 1706 2068 1710 2071
rect 1930 2068 2094 2071
rect 2098 2068 2294 2071
rect 2330 2068 2406 2071
rect 2426 2068 2470 2071
rect 2474 2068 2478 2071
rect 2482 2068 2526 2071
rect 2586 2068 2590 2071
rect 2602 2068 2622 2071
rect 2690 2068 2710 2071
rect 2722 2068 2726 2071
rect 2730 2068 2758 2071
rect 2858 2068 2878 2071
rect 2954 2068 2982 2071
rect 3010 2068 3182 2071
rect 3378 2068 3518 2071
rect 3618 2068 3630 2071
rect 3706 2068 3718 2071
rect 3746 2068 3750 2071
rect 3818 2068 4046 2071
rect 4154 2068 4246 2071
rect 4346 2068 4358 2071
rect 4394 2068 4438 2071
rect 4474 2068 4510 2071
rect 4570 2068 4574 2071
rect 214 2061 217 2068
rect 270 2061 273 2068
rect 214 2058 273 2061
rect 298 2058 310 2061
rect 318 2061 321 2068
rect 318 2058 342 2061
rect 406 2061 409 2068
rect 1246 2062 1249 2068
rect 386 2058 409 2061
rect 482 2058 526 2061
rect 530 2058 638 2061
rect 770 2058 806 2061
rect 810 2058 862 2061
rect 874 2058 878 2061
rect 994 2058 1030 2061
rect 1034 2058 1046 2061
rect 1058 2058 1094 2061
rect 1266 2058 1326 2061
rect 1470 2061 1473 2068
rect 1470 2058 1534 2061
rect 1550 2061 1553 2068
rect 1686 2062 1689 2068
rect 1550 2058 1566 2061
rect 1594 2058 1638 2061
rect 1666 2058 1673 2061
rect 1786 2059 1790 2061
rect 1786 2058 1793 2059
rect 1886 2061 1889 2068
rect 1834 2058 1990 2061
rect 1994 2058 2102 2061
rect 2122 2059 2126 2061
rect 2118 2058 2126 2059
rect 2138 2058 2278 2061
rect 2298 2058 2318 2061
rect 2410 2058 2414 2061
rect 2442 2058 2446 2061
rect 2450 2058 2478 2061
rect 2482 2058 2518 2061
rect 2634 2058 2646 2061
rect 2682 2058 2758 2061
rect 2762 2058 2934 2061
rect 2938 2058 3014 2061
rect 3074 2058 3078 2061
rect 3082 2058 3094 2061
rect 3114 2058 3190 2061
rect 3226 2058 3254 2061
rect 3258 2058 3286 2061
rect 3290 2058 3334 2061
rect 3394 2058 3406 2061
rect 3410 2058 3470 2061
rect 3474 2058 3590 2061
rect 3658 2058 3686 2061
rect 3706 2058 3726 2061
rect 3730 2058 3766 2061
rect 3778 2058 4014 2061
rect 4170 2058 4302 2061
rect 4306 2058 4318 2061
rect 4322 2058 4374 2061
rect 4434 2058 4478 2061
rect 4482 2058 4494 2061
rect 4554 2058 4558 2061
rect 4562 2058 4598 2061
rect 1670 2052 1673 2058
rect -26 2051 -22 2052
rect -26 2048 6 2051
rect 254 2048 358 2051
rect 458 2048 462 2051
rect 498 2048 521 2051
rect 530 2048 622 2051
rect 626 2048 646 2051
rect 658 2048 806 2051
rect 882 2048 894 2051
rect 978 2048 982 2051
rect 986 2048 1134 2051
rect 1282 2048 1302 2051
rect 1306 2048 1342 2051
rect 1378 2048 1390 2051
rect 1394 2048 1566 2051
rect 1742 2051 1745 2058
rect 1742 2048 2158 2051
rect 2170 2048 2190 2051
rect 2202 2048 2302 2051
rect 2410 2048 2494 2051
rect 2530 2048 2574 2051
rect 2778 2048 2862 2051
rect 2898 2048 2918 2051
rect 2930 2048 2950 2051
rect 3094 2051 3097 2058
rect 3094 2048 3150 2051
rect 3178 2048 3230 2051
rect 3370 2048 3374 2051
rect 3382 2051 3385 2058
rect 3774 2052 3777 2058
rect 4454 2052 4457 2058
rect 3382 2048 3438 2051
rect 3578 2048 3582 2051
rect 3626 2048 3630 2051
rect 3762 2048 3766 2051
rect 3802 2048 3806 2051
rect 3882 2048 3886 2051
rect 3930 2048 3950 2051
rect 4006 2048 4182 2051
rect 4194 2048 4238 2051
rect 4290 2048 4350 2051
rect 254 2042 257 2048
rect 470 2042 473 2048
rect 26 2038 142 2041
rect 146 2038 246 2041
rect 322 2038 350 2041
rect 354 2038 470 2041
rect 474 2038 502 2041
rect 518 2041 521 2048
rect 1326 2042 1329 2048
rect 3782 2042 3785 2048
rect 518 2038 710 2041
rect 794 2038 798 2041
rect 842 2038 886 2041
rect 1162 2038 1310 2041
rect 1402 2038 1694 2041
rect 1714 2038 1758 2041
rect 2050 2038 3494 2041
rect 3498 2038 3774 2041
rect 3794 2038 3814 2041
rect 4006 2041 4009 2048
rect 3842 2038 4009 2041
rect 4014 2038 4022 2041
rect 4026 2038 4030 2041
rect 4098 2038 4542 2041
rect 4546 2038 4550 2041
rect 170 2028 494 2031
rect 682 2028 1430 2031
rect 1578 2028 1630 2031
rect 1634 2028 1721 2031
rect 1866 2028 2006 2031
rect 2250 2028 2254 2031
rect 2270 2028 2278 2031
rect 2282 2028 2326 2031
rect 2354 2028 2438 2031
rect 2714 2028 2750 2031
rect 2754 2028 2766 2031
rect 2806 2028 2814 2031
rect 2818 2028 2870 2031
rect 2874 2028 2974 2031
rect 3186 2028 3246 2031
rect 3266 2028 3782 2031
rect 3786 2028 4126 2031
rect 4210 2028 4406 2031
rect 4410 2028 4462 2031
rect 490 2018 766 2021
rect 1338 2018 1366 2021
rect 1502 2021 1505 2028
rect 1718 2022 1721 2028
rect 1502 2018 1646 2021
rect 1666 2018 1702 2021
rect 1730 2018 1806 2021
rect 1810 2018 2598 2021
rect 2602 2018 2662 2021
rect 2890 2018 3022 2021
rect 3090 2018 3302 2021
rect 3306 2018 3326 2021
rect 3330 2018 3350 2021
rect 3362 2018 3614 2021
rect 3618 2018 3625 2021
rect 3802 2018 3966 2021
rect 3970 2018 4046 2021
rect 4114 2018 4182 2021
rect 4186 2018 4278 2021
rect 4282 2018 4302 2021
rect 4330 2018 4342 2021
rect 122 2008 478 2011
rect 826 2008 1510 2011
rect 1898 2008 1902 2011
rect 1922 2008 2054 2011
rect 2058 2008 2494 2011
rect 2610 2008 2646 2011
rect 2650 2008 2726 2011
rect 2882 2008 3150 2011
rect 3194 2008 3398 2011
rect 3754 2008 3974 2011
rect 3978 2008 3998 2011
rect 4426 2008 4534 2011
rect 4538 2008 4582 2011
rect 496 2003 498 2007
rect 502 2003 505 2007
rect 510 2003 512 2007
rect 1520 2003 1522 2007
rect 1526 2003 1529 2007
rect 1534 2003 1536 2007
rect 2544 2003 2546 2007
rect 2550 2003 2553 2007
rect 2558 2003 2560 2007
rect 3568 2003 3570 2007
rect 3574 2003 3577 2007
rect 3582 2003 3584 2007
rect 50 1998 150 2001
rect 1194 1998 1222 2001
rect 1434 1998 1438 2001
rect 1546 1998 1822 2001
rect 2106 1998 2214 2001
rect 2258 1998 2286 2001
rect 2570 1998 2894 2001
rect 2898 1998 3142 2001
rect 3778 1998 3854 2001
rect 3866 1998 3934 2001
rect 4058 1998 4102 2001
rect 4106 1998 4398 2001
rect 98 1988 342 1991
rect 414 1991 417 1998
rect 3686 1992 3689 1998
rect 346 1988 558 1991
rect 642 1988 694 1991
rect 894 1988 902 1991
rect 906 1988 1718 1991
rect 1730 1988 2478 1991
rect 2482 1988 2534 1991
rect 3006 1988 3014 1991
rect 3018 1988 3174 1991
rect 3178 1988 3182 1991
rect 3522 1988 3678 1991
rect 3810 1988 3838 1991
rect 3842 1988 4054 1991
rect 4194 1988 4246 1991
rect 258 1978 294 1981
rect 298 1978 366 1981
rect 482 1978 606 1981
rect 610 1978 934 1981
rect 1098 1978 1542 1981
rect 1650 1978 1710 1981
rect 1714 1978 1782 1981
rect 1858 1978 1974 1981
rect 2202 1978 2302 1981
rect 2314 1978 2342 1981
rect 2354 1978 2566 1981
rect 2630 1981 2633 1988
rect 2630 1978 2670 1981
rect 2750 1981 2753 1988
rect 2750 1978 2862 1981
rect 2970 1978 3225 1981
rect 3458 1978 3614 1981
rect 3618 1978 3670 1981
rect 3674 1978 4206 1981
rect 4346 1978 4398 1981
rect -26 1971 -22 1972
rect 30 1971 33 1978
rect -26 1968 33 1971
rect 218 1968 374 1971
rect 378 1968 382 1971
rect 398 1971 401 1978
rect 398 1968 526 1971
rect 630 1968 646 1971
rect 706 1968 790 1971
rect 930 1968 990 1971
rect 1122 1968 1174 1971
rect 1602 1968 1678 1971
rect 1762 1968 1854 1971
rect 1898 1968 1934 1971
rect 1938 1968 1958 1971
rect 2010 1968 2062 1971
rect 2086 1971 2089 1978
rect 3222 1972 3225 1978
rect 2086 1968 3022 1971
rect 3162 1968 3166 1971
rect 3226 1968 3358 1971
rect 3514 1968 3518 1971
rect 3534 1968 3542 1971
rect 3546 1968 3550 1971
rect 3562 1968 3678 1971
rect 3706 1968 3710 1971
rect 3722 1968 3726 1971
rect 3818 1968 4150 1971
rect 4194 1968 4246 1971
rect 4250 1968 4294 1971
rect 4306 1968 4390 1971
rect 4406 1971 4409 1978
rect 4494 1971 4497 1978
rect 4394 1968 4401 1971
rect 4406 1968 4497 1971
rect 630 1962 633 1968
rect 26 1958 54 1961
rect 122 1958 270 1961
rect 274 1958 318 1961
rect 330 1958 334 1961
rect 402 1958 422 1961
rect 554 1958 558 1961
rect 802 1958 1334 1961
rect 1522 1958 1614 1961
rect 1618 1958 1638 1961
rect 1722 1958 1774 1961
rect 1802 1958 2430 1961
rect 2446 1958 2454 1961
rect 2458 1958 2470 1961
rect 2474 1958 2518 1961
rect 2674 1958 2678 1961
rect 2710 1958 2838 1961
rect 2842 1958 2910 1961
rect 3034 1958 3038 1961
rect 3042 1958 3046 1961
rect 3074 1958 3254 1961
rect 3258 1958 3374 1961
rect 3490 1958 3654 1961
rect 3658 1958 3814 1961
rect 3826 1958 3830 1961
rect 3842 1958 3934 1961
rect 3962 1958 3966 1961
rect 3986 1958 4078 1961
rect 4162 1958 4166 1961
rect 4170 1958 4318 1961
rect 4402 1958 4406 1961
rect -26 1951 -22 1952
rect -26 1948 6 1951
rect 314 1948 318 1951
rect 478 1948 510 1951
rect 522 1948 534 1951
rect 594 1948 614 1951
rect 662 1951 665 1958
rect 678 1951 681 1958
rect 662 1948 681 1951
rect 1050 1948 1126 1951
rect 1138 1948 1142 1951
rect 1170 1948 1206 1951
rect 1234 1948 1262 1951
rect 1266 1948 1270 1951
rect 1366 1951 1369 1958
rect 2710 1952 2713 1958
rect 1366 1948 1454 1951
rect 1490 1948 1510 1951
rect 1634 1948 1654 1951
rect 1738 1948 1742 1951
rect 1754 1948 2006 1951
rect 2010 1948 2054 1951
rect 2058 1948 2094 1951
rect 2098 1948 2134 1951
rect 2138 1948 2150 1951
rect 2298 1948 2374 1951
rect 2386 1948 2422 1951
rect 2426 1948 2494 1951
rect 2498 1948 2526 1951
rect 2530 1948 2534 1951
rect 2690 1948 2702 1951
rect 2770 1948 2878 1951
rect 2890 1948 2902 1951
rect 2946 1948 3150 1951
rect 3202 1948 3206 1951
rect 3218 1948 3230 1951
rect 3290 1948 3294 1951
rect 3298 1948 3318 1951
rect 3434 1948 3542 1951
rect 3602 1948 3638 1951
rect 3642 1948 3665 1951
rect 3714 1948 3718 1951
rect 3754 1948 3830 1951
rect 3842 1948 3870 1951
rect 3890 1948 3894 1951
rect 3906 1948 3926 1951
rect 3930 1948 3958 1951
rect 3962 1948 4006 1951
rect 4010 1948 4062 1951
rect 4066 1948 4134 1951
rect 4138 1948 4142 1951
rect 4194 1948 4198 1951
rect 4234 1948 4294 1951
rect 4298 1948 4350 1951
rect 4410 1948 4558 1951
rect 478 1942 481 1948
rect 210 1938 249 1941
rect 282 1938 382 1941
rect 538 1938 550 1941
rect 570 1938 582 1941
rect 814 1941 817 1948
rect 762 1938 817 1941
rect 906 1938 910 1941
rect 930 1938 1070 1941
rect 1138 1938 1185 1941
rect 1218 1938 1238 1941
rect 1258 1938 1270 1941
rect 1274 1938 1286 1941
rect 1406 1938 1502 1941
rect 1538 1938 1558 1941
rect 1562 1938 1566 1941
rect 1622 1941 1625 1948
rect 1570 1938 1625 1941
rect 1642 1938 1662 1941
rect 1706 1938 1830 1941
rect 1834 1938 1870 1941
rect 1906 1938 1910 1941
rect 1914 1938 1934 1941
rect 1998 1938 2070 1941
rect 2114 1938 2118 1941
rect 2322 1938 2606 1941
rect 2626 1940 2646 1941
rect 2622 1938 2646 1940
rect 2670 1941 2673 1948
rect 2710 1941 2713 1948
rect 2670 1938 2713 1941
rect 3662 1942 3665 1948
rect 2730 1940 2854 1941
rect 2726 1938 2854 1940
rect 2858 1938 2942 1941
rect 2946 1938 2958 1941
rect 2978 1938 3142 1941
rect 3146 1938 3158 1941
rect 3250 1938 3254 1941
rect 3306 1938 3342 1941
rect 3434 1938 3438 1941
rect 3474 1938 3494 1941
rect 3498 1938 3534 1941
rect 3666 1938 3742 1941
rect 3826 1938 3838 1941
rect 3882 1938 3918 1941
rect 3938 1938 3993 1941
rect 4050 1938 4078 1941
rect 4122 1938 4358 1941
rect 4362 1938 4414 1941
rect 4498 1938 4526 1941
rect 4530 1938 4566 1941
rect 246 1932 249 1938
rect 306 1928 830 1931
rect 978 1928 1057 1931
rect 1082 1928 1126 1931
rect 1138 1928 1142 1931
rect 1182 1931 1185 1938
rect 1294 1932 1297 1938
rect 1406 1932 1409 1938
rect 1182 1928 1262 1931
rect 1554 1928 1590 1931
rect 1594 1928 1614 1931
rect 1618 1928 1798 1931
rect 1826 1928 1830 1931
rect 1842 1928 1870 1931
rect 1998 1931 2001 1938
rect 1938 1928 2001 1931
rect 2010 1928 2014 1931
rect 2182 1931 2185 1938
rect 2182 1928 2190 1931
rect 2278 1931 2281 1938
rect 2258 1928 2398 1931
rect 2402 1928 2422 1931
rect 2538 1928 2558 1931
rect 2562 1928 2686 1931
rect 2730 1928 2734 1931
rect 2754 1928 2798 1931
rect 2842 1928 2889 1931
rect 2938 1928 2942 1931
rect 3002 1928 3038 1931
rect 3114 1928 3166 1931
rect 3414 1931 3417 1938
rect 3378 1928 3417 1931
rect 3538 1928 3718 1931
rect 3758 1931 3761 1938
rect 3846 1932 3849 1938
rect 3990 1932 3993 1938
rect 3758 1928 3782 1931
rect 3938 1928 3958 1931
rect 4026 1928 4030 1931
rect 4042 1928 4049 1931
rect 4058 1928 4070 1931
rect 4154 1928 4166 1931
rect 4178 1928 4406 1931
rect 4458 1928 4470 1931
rect 4490 1928 4550 1931
rect 4554 1928 4566 1931
rect 4570 1928 4582 1931
rect 1054 1922 1057 1928
rect 50 1918 230 1921
rect 234 1918 550 1921
rect 554 1918 734 1921
rect 1150 1921 1153 1928
rect 1150 1918 1198 1921
rect 1286 1921 1289 1928
rect 1226 1918 1334 1921
rect 1474 1918 1494 1921
rect 1498 1918 1566 1921
rect 1634 1918 1934 1921
rect 1946 1918 1998 1921
rect 2006 1918 2110 1921
rect 2154 1918 2422 1921
rect 2462 1921 2465 1928
rect 2886 1922 2889 1928
rect 2462 1918 2654 1921
rect 2658 1918 2702 1921
rect 3042 1918 3302 1921
rect 3314 1918 3334 1921
rect 3438 1921 3441 1928
rect 4046 1922 4049 1928
rect 3338 1918 3758 1921
rect 3762 1918 3998 1921
rect 4066 1918 4142 1921
rect 4258 1918 4262 1921
rect 4298 1918 4302 1921
rect 4386 1918 4446 1921
rect 4522 1918 4566 1921
rect 266 1908 382 1911
rect 482 1908 550 1911
rect 554 1908 670 1911
rect 674 1908 782 1911
rect 1098 1908 1158 1911
rect 1162 1908 1206 1911
rect 1250 1908 1254 1911
rect 1538 1908 1886 1911
rect 1890 1908 1982 1911
rect 2006 1911 2009 1918
rect 4518 1912 4521 1918
rect 1994 1908 2009 1911
rect 2162 1908 2182 1911
rect 2242 1908 2398 1911
rect 2402 1908 2454 1911
rect 2474 1908 2494 1911
rect 2602 1908 2622 1911
rect 2626 1908 2638 1911
rect 2650 1908 2734 1911
rect 3122 1908 3630 1911
rect 3650 1908 3686 1911
rect 3690 1908 3718 1911
rect 3794 1908 3942 1911
rect 3962 1908 3966 1911
rect 3986 1908 4014 1911
rect 4018 1908 4070 1911
rect 4250 1908 4374 1911
rect 4410 1908 4422 1911
rect 4442 1908 4510 1911
rect 1000 1903 1002 1907
rect 1006 1903 1009 1907
rect 1014 1903 1016 1907
rect 2024 1903 2026 1907
rect 2030 1903 2033 1907
rect 2038 1903 2040 1907
rect 3048 1903 3050 1907
rect 3054 1903 3057 1907
rect 3062 1903 3064 1907
rect 4080 1903 4082 1907
rect 4086 1903 4089 1907
rect 4094 1903 4096 1907
rect 326 1898 902 1901
rect 906 1898 934 1901
rect 1114 1898 1742 1901
rect 1802 1898 1950 1901
rect 2146 1898 3038 1901
rect 3354 1898 3766 1901
rect 3778 1898 3798 1901
rect 3802 1898 3830 1901
rect 3834 1898 3854 1901
rect 3858 1898 3870 1901
rect 3922 1898 3974 1901
rect 4042 1898 4054 1901
rect 4210 1898 4294 1901
rect 4298 1898 4342 1901
rect 4354 1898 4366 1901
rect 4370 1898 4430 1901
rect 4434 1898 4510 1901
rect 326 1892 329 1898
rect 26 1888 326 1891
rect 690 1888 726 1891
rect 738 1888 766 1891
rect 1026 1888 1118 1891
rect 1130 1888 1185 1891
rect 1182 1882 1185 1888
rect 1410 1888 1729 1891
rect 1890 1888 2078 1891
rect 2082 1888 2246 1891
rect 2314 1888 2566 1891
rect 2634 1888 2710 1891
rect 2802 1888 2870 1891
rect 3026 1888 3078 1891
rect 3166 1888 3750 1891
rect 3766 1891 3769 1898
rect 3766 1888 4398 1891
rect 4402 1888 4486 1891
rect 4490 1888 4526 1891
rect 1382 1882 1385 1888
rect 1726 1882 1729 1888
rect 410 1878 446 1881
rect 450 1878 614 1881
rect 746 1878 766 1881
rect 770 1878 822 1881
rect 1190 1878 1310 1881
rect 1354 1878 1366 1881
rect 1386 1878 1422 1881
rect 1770 1878 1774 1881
rect 1906 1878 1918 1881
rect 1938 1878 1974 1881
rect 1978 1878 2057 1881
rect 2066 1878 2105 1881
rect 2186 1878 2206 1881
rect 2210 1878 2302 1881
rect 2338 1878 2342 1881
rect 2418 1878 2478 1881
rect 2490 1878 2694 1881
rect 2706 1878 2742 1881
rect 2754 1878 2766 1881
rect 2770 1878 2878 1881
rect 2882 1878 2942 1881
rect 2946 1878 2950 1881
rect 2978 1878 3038 1881
rect 3042 1878 3046 1881
rect 3086 1881 3089 1888
rect 3166 1882 3169 1888
rect 3086 1878 3166 1881
rect 3202 1878 3270 1881
rect 3554 1878 3630 1881
rect 3682 1878 3694 1881
rect 3714 1878 3734 1881
rect 3754 1878 3766 1881
rect 3842 1878 3862 1881
rect 3866 1878 3886 1881
rect 3890 1878 3918 1881
rect 3946 1878 3958 1881
rect 3970 1878 4006 1881
rect 4026 1878 4046 1881
rect 4050 1878 4086 1881
rect 4090 1878 4118 1881
rect 4130 1878 4134 1881
rect 4202 1878 4214 1881
rect 4218 1878 4230 1881
rect 4258 1878 4326 1881
rect 4458 1878 4462 1881
rect 4514 1878 4542 1881
rect 4582 1881 4585 1888
rect 4562 1878 4585 1881
rect -26 1871 -22 1872
rect 6 1871 9 1878
rect 214 1872 217 1878
rect -26 1868 9 1871
rect 134 1868 153 1871
rect 586 1868 598 1871
rect 626 1868 638 1871
rect 642 1868 646 1871
rect 1030 1871 1033 1878
rect 962 1868 1033 1871
rect 1190 1871 1193 1878
rect 1122 1868 1193 1871
rect 1262 1868 1278 1871
rect 1330 1868 1374 1871
rect 1550 1871 1553 1878
rect 1506 1868 1553 1871
rect 1566 1872 1569 1878
rect 1638 1872 1641 1878
rect 1722 1868 1742 1871
rect 1746 1868 1782 1871
rect 1806 1871 1809 1878
rect 1806 1868 1990 1871
rect 2054 1871 2057 1878
rect 2102 1872 2105 1878
rect 2054 1868 2062 1871
rect 2370 1868 2374 1871
rect 2626 1868 2630 1871
rect 2658 1868 2662 1871
rect 2694 1871 2697 1878
rect 4254 1872 4257 1878
rect 2694 1868 3190 1871
rect 3194 1868 3390 1871
rect 3434 1868 3574 1871
rect 3586 1868 3806 1871
rect 3810 1868 4222 1871
rect 4226 1868 4238 1871
rect 4242 1868 4246 1871
rect 4270 1868 4366 1871
rect 4442 1868 4478 1871
rect 4482 1868 4494 1871
rect 4506 1868 4542 1871
rect 4546 1868 4598 1871
rect 134 1862 137 1868
rect 150 1862 153 1868
rect 154 1858 230 1861
rect 250 1859 254 1861
rect 350 1862 353 1868
rect 250 1858 257 1859
rect 370 1858 406 1861
rect 410 1858 526 1861
rect 610 1858 630 1861
rect 710 1861 713 1868
rect 666 1858 713 1861
rect 806 1861 809 1868
rect 838 1861 841 1868
rect 806 1858 841 1861
rect 870 1861 873 1868
rect 1262 1862 1265 1868
rect 870 1858 918 1861
rect 1202 1858 1230 1861
rect 1326 1861 1329 1868
rect 1282 1858 1329 1861
rect 1354 1858 1630 1861
rect 1634 1858 1641 1861
rect 1690 1858 1694 1861
rect 1746 1858 1750 1861
rect 1798 1861 1801 1868
rect 1770 1858 1801 1861
rect 1866 1858 1894 1861
rect 1922 1858 1982 1861
rect 2002 1858 2014 1861
rect 2082 1858 2118 1861
rect 2146 1858 2214 1861
rect 2230 1861 2233 1868
rect 4270 1862 4273 1868
rect 2230 1858 2294 1861
rect 2426 1858 2446 1861
rect 2530 1858 2598 1861
rect 2698 1858 2774 1861
rect 2782 1858 2790 1861
rect 2794 1858 2814 1861
rect 2834 1858 2838 1861
rect 2866 1858 2886 1861
rect 2906 1858 2910 1861
rect 2938 1858 2950 1861
rect 2994 1858 2998 1861
rect 3210 1858 3382 1861
rect 3386 1858 3398 1861
rect 3418 1858 3462 1861
rect 3498 1858 3510 1861
rect 3658 1858 3670 1861
rect 3674 1858 3750 1861
rect 3770 1858 3798 1861
rect 3930 1858 4094 1861
rect 4138 1858 4158 1861
rect 4162 1858 4262 1861
rect 4282 1858 4398 1861
rect 4402 1858 4566 1861
rect -26 1851 -22 1852
rect -26 1848 30 1851
rect 402 1848 430 1851
rect 434 1848 438 1851
rect 442 1848 606 1851
rect 794 1848 838 1851
rect 1178 1848 1246 1851
rect 1298 1848 1414 1851
rect 1458 1848 1662 1851
rect 1690 1848 1734 1851
rect 1738 1848 1774 1851
rect 1778 1848 1814 1851
rect 1834 1848 1894 1851
rect 226 1838 342 1841
rect 622 1841 625 1848
rect 386 1838 625 1841
rect 638 1841 641 1848
rect 638 1838 790 1841
rect 906 1838 910 1841
rect 1186 1838 1342 1841
rect 1662 1841 1665 1848
rect 2174 1842 2177 1851
rect 2186 1848 2190 1851
rect 2230 1848 2254 1851
rect 2306 1848 2422 1851
rect 2426 1848 2430 1851
rect 2434 1848 2486 1851
rect 2514 1848 2558 1851
rect 2562 1848 2598 1851
rect 2722 1848 2793 1851
rect 2810 1848 3070 1851
rect 3162 1848 3166 1851
rect 3202 1848 3238 1851
rect 3242 1848 3566 1851
rect 3570 1848 3638 1851
rect 3898 1848 3942 1851
rect 4002 1848 4014 1851
rect 4018 1848 4038 1851
rect 4282 1848 4286 1851
rect 4322 1848 4414 1851
rect 4474 1848 4486 1851
rect 4490 1848 4561 1851
rect 2230 1842 2233 1848
rect 1662 1838 2166 1841
rect 2262 1841 2265 1848
rect 2790 1842 2793 1848
rect 2262 1838 2286 1841
rect 2490 1838 2614 1841
rect 2650 1838 2670 1841
rect 2922 1838 2942 1841
rect 3034 1838 3222 1841
rect 3290 1838 3350 1841
rect 3418 1838 3473 1841
rect 3522 1838 3838 1841
rect 3866 1838 4030 1841
rect 4110 1841 4113 1848
rect 4558 1842 4561 1848
rect 4110 1838 4158 1841
rect 4290 1838 4462 1841
rect 3470 1832 3473 1838
rect 314 1828 334 1831
rect 354 1828 558 1831
rect 1098 1828 1222 1831
rect 1634 1828 1734 1831
rect 1842 1828 1846 1831
rect 1946 1828 2246 1831
rect 2274 1828 2502 1831
rect 2506 1828 2630 1831
rect 2754 1828 2902 1831
rect 2946 1828 3182 1831
rect 3258 1828 3358 1831
rect 3474 1828 3494 1831
rect 3602 1828 3822 1831
rect 3826 1828 3846 1831
rect 4026 1828 4310 1831
rect 4314 1828 4558 1831
rect 490 1818 678 1821
rect 866 1818 990 1821
rect 994 1818 1046 1821
rect 1698 1818 2206 1821
rect 2254 1821 2257 1828
rect 2254 1818 2566 1821
rect 2942 1821 2945 1828
rect 2850 1818 2945 1821
rect 3234 1818 3270 1821
rect 3274 1818 3310 1821
rect 3578 1818 4110 1821
rect 962 1808 1502 1811
rect 1570 1808 1782 1811
rect 1786 1808 1926 1811
rect 2098 1808 2134 1811
rect 2154 1808 2238 1811
rect 2578 1808 2710 1811
rect 2834 1808 2910 1811
rect 3330 1808 3446 1811
rect 3498 1808 3558 1811
rect 3738 1808 3782 1811
rect 3810 1808 3846 1811
rect 3858 1808 3934 1811
rect 4034 1808 4446 1811
rect 4450 1808 4518 1811
rect 496 1803 498 1807
rect 502 1803 505 1807
rect 510 1803 512 1807
rect 1520 1803 1522 1807
rect 1526 1803 1529 1807
rect 1534 1803 1536 1807
rect 554 1798 582 1801
rect 1162 1798 1190 1801
rect 1194 1798 1198 1801
rect 1762 1798 1902 1801
rect 2134 1801 2137 1808
rect 2544 1803 2546 1807
rect 2550 1803 2553 1807
rect 2558 1803 2560 1807
rect 3568 1803 3570 1807
rect 3574 1803 3577 1807
rect 3582 1803 3584 1807
rect 2134 1798 2198 1801
rect 2406 1798 2534 1801
rect 2650 1798 2694 1801
rect 2770 1798 2854 1801
rect 2858 1798 2878 1801
rect 3154 1798 3158 1801
rect 3162 1798 3366 1801
rect 3386 1798 3390 1801
rect 3402 1798 3486 1801
rect 3530 1798 3550 1801
rect 3770 1798 3862 1801
rect 3882 1798 3974 1801
rect 4002 1798 4366 1801
rect 4434 1798 4438 1801
rect 2406 1792 2409 1798
rect -26 1791 -22 1792
rect -26 1788 38 1791
rect 306 1788 422 1791
rect 1194 1788 1206 1791
rect 1378 1788 1478 1791
rect 1490 1788 1726 1791
rect 1770 1788 1910 1791
rect 1938 1788 1966 1791
rect 1970 1788 2158 1791
rect 2218 1788 2406 1791
rect 2522 1788 3102 1791
rect 3138 1788 3142 1791
rect 3194 1788 3302 1791
rect 3306 1788 3366 1791
rect 3370 1788 3598 1791
rect 3626 1788 3806 1791
rect 3810 1788 3886 1791
rect 3970 1788 3974 1791
rect 3978 1788 4094 1791
rect 4226 1788 4246 1791
rect 4250 1788 4286 1791
rect 394 1778 574 1781
rect 786 1778 1574 1781
rect 1690 1778 2694 1781
rect 2810 1778 2814 1781
rect 2818 1778 3814 1781
rect 3818 1778 3942 1781
rect 3946 1778 4070 1781
rect 4226 1778 4318 1781
rect 4434 1778 4478 1781
rect -26 1771 -22 1772
rect 6 1771 9 1778
rect -26 1768 9 1771
rect 314 1768 318 1771
rect 330 1768 334 1771
rect 554 1768 590 1771
rect 758 1771 761 1778
rect 738 1768 838 1771
rect 1026 1768 1054 1771
rect 1058 1768 1166 1771
rect 1202 1768 1254 1771
rect 1282 1768 1366 1771
rect 1586 1768 1590 1771
rect 1638 1771 1641 1778
rect 1638 1768 1686 1771
rect 1698 1768 1718 1771
rect 1738 1768 1742 1771
rect 1746 1768 1822 1771
rect 1826 1768 1854 1771
rect 1858 1768 1886 1771
rect 1906 1768 2126 1771
rect 2138 1768 2174 1771
rect 2230 1768 2382 1771
rect 2386 1768 2446 1771
rect 2618 1768 2646 1771
rect 2662 1768 2670 1771
rect 2674 1768 3006 1771
rect 3138 1768 3254 1771
rect 3346 1768 3350 1771
rect 3362 1768 3902 1771
rect 4058 1768 4166 1771
rect 4390 1771 4393 1778
rect 4314 1768 4393 1771
rect 2230 1762 2233 1768
rect -26 1758 54 1761
rect 258 1758 366 1761
rect 370 1758 486 1761
rect 490 1758 638 1761
rect 722 1758 894 1761
rect 1050 1758 1094 1761
rect 1130 1758 1134 1761
rect 1186 1758 1270 1761
rect 1514 1758 1606 1761
rect 1610 1758 1950 1761
rect 1954 1758 2070 1761
rect 2074 1758 2182 1761
rect 2186 1758 2214 1761
rect 2218 1758 2222 1761
rect 2250 1758 2318 1761
rect 2322 1758 2342 1761
rect 2474 1758 2510 1761
rect 2594 1758 2662 1761
rect 2690 1758 2694 1761
rect 2698 1758 2814 1761
rect 2862 1758 2934 1761
rect 3162 1758 3166 1761
rect 3170 1758 3270 1761
rect 3290 1758 3310 1761
rect 3354 1758 3414 1761
rect 3450 1758 3462 1761
rect 3514 1758 3598 1761
rect 3682 1758 3686 1761
rect 3762 1758 3766 1761
rect 3778 1758 4206 1761
rect 4402 1758 4454 1761
rect 4538 1758 4574 1761
rect -26 1752 -23 1758
rect -26 1748 -22 1752
rect 46 1748 54 1751
rect 58 1748 110 1751
rect 114 1748 246 1751
rect 250 1748 278 1751
rect 282 1748 374 1751
rect 434 1748 454 1751
rect 602 1748 710 1751
rect 730 1748 830 1751
rect 834 1748 846 1751
rect 1002 1748 1006 1751
rect 1034 1748 1086 1751
rect 1258 1748 1278 1751
rect 1306 1748 1326 1751
rect 1422 1751 1425 1758
rect 1422 1748 1446 1751
rect 1450 1748 1502 1751
rect 1546 1748 1598 1751
rect 1602 1748 1782 1751
rect 1786 1748 2006 1751
rect 2010 1748 2054 1751
rect 2178 1748 2230 1751
rect 2234 1748 2262 1751
rect 2266 1748 2270 1751
rect 2610 1748 2678 1751
rect 2682 1748 2718 1751
rect 2738 1748 2766 1751
rect 2822 1751 2825 1758
rect 2770 1748 2825 1751
rect 2862 1752 2865 1758
rect 3630 1752 3633 1758
rect 4318 1752 4321 1758
rect 4374 1752 4377 1758
rect 2970 1748 2974 1751
rect 2994 1748 2998 1751
rect 3042 1748 3126 1751
rect 3194 1748 3198 1751
rect 3282 1748 3318 1751
rect 3322 1748 3334 1751
rect 3434 1748 3502 1751
rect 3538 1748 3566 1751
rect 3578 1748 3606 1751
rect 3730 1748 3790 1751
rect 3794 1748 3830 1751
rect 3842 1748 3865 1751
rect 3874 1748 3910 1751
rect 3994 1748 4006 1751
rect 4114 1748 4134 1751
rect 4178 1748 4182 1751
rect 4234 1748 4278 1751
rect 4354 1748 4358 1751
rect 4402 1748 4406 1751
rect 4426 1748 4518 1751
rect 4522 1748 4590 1751
rect 74 1738 238 1741
rect 242 1738 254 1741
rect 262 1738 310 1741
rect 802 1738 806 1741
rect 1098 1738 1110 1741
rect 1246 1741 1249 1748
rect 1390 1742 1393 1748
rect 1246 1738 1262 1741
rect 1314 1738 1342 1741
rect 1586 1738 1774 1741
rect 1778 1738 1966 1741
rect 1970 1738 2030 1741
rect 2190 1738 2246 1741
rect 2258 1738 2262 1741
rect 2266 1738 2318 1741
rect 2322 1738 2358 1741
rect 2362 1738 2462 1741
rect 2466 1738 2470 1741
rect 2490 1738 2494 1741
rect 2498 1738 2614 1741
rect 2630 1738 2726 1741
rect 2730 1738 2814 1741
rect 2818 1738 2910 1741
rect 2938 1738 3094 1741
rect 3162 1738 3190 1741
rect 3194 1738 3198 1741
rect 3234 1738 3238 1741
rect 3266 1738 3294 1741
rect 3306 1738 3390 1741
rect 3394 1738 3406 1741
rect 3426 1738 3470 1741
rect 3498 1738 3518 1741
rect 3546 1738 3550 1741
rect 3554 1738 3622 1741
rect 3626 1738 3678 1741
rect 3834 1738 3838 1741
rect 3842 1738 3854 1741
rect 3862 1741 3865 1748
rect 3918 1742 3921 1748
rect 3982 1742 3985 1748
rect 3862 1738 3870 1741
rect 4146 1738 4174 1741
rect 4178 1738 4190 1741
rect 4250 1738 4254 1741
rect 4290 1738 4294 1741
rect 4298 1738 4350 1741
rect 4354 1738 4542 1741
rect 262 1732 265 1738
rect 314 1728 318 1731
rect 354 1728 366 1731
rect 674 1728 766 1731
rect 1078 1731 1081 1738
rect 1198 1732 1201 1738
rect 2190 1732 2193 1738
rect 2630 1732 2633 1738
rect 978 1728 1102 1731
rect 1122 1728 1182 1731
rect 1234 1728 1254 1731
rect 1346 1728 1358 1731
rect 1362 1728 1465 1731
rect 1666 1728 1710 1731
rect 1714 1728 1718 1731
rect 1730 1728 1798 1731
rect 1802 1728 1830 1731
rect 1834 1728 1878 1731
rect 1882 1728 2118 1731
rect 2122 1728 2142 1731
rect 2250 1728 2278 1731
rect 2298 1728 2326 1731
rect 2330 1728 2366 1731
rect 2498 1728 2518 1731
rect 2522 1728 2534 1731
rect 2594 1728 2622 1731
rect 2650 1728 2654 1731
rect 2658 1728 2702 1731
rect 2818 1728 2862 1731
rect 2902 1728 3062 1731
rect 3122 1728 3126 1731
rect 3130 1728 3169 1731
rect 3186 1728 3206 1731
rect 3338 1728 3366 1731
rect 3514 1728 3542 1731
rect 3570 1728 3574 1731
rect 3618 1728 3758 1731
rect 3762 1728 3878 1731
rect 3930 1728 3942 1731
rect 3962 1728 4046 1731
rect 4278 1728 4286 1731
rect 4378 1728 4486 1731
rect 4514 1728 4590 1731
rect 258 1718 286 1721
rect 674 1718 1454 1721
rect 1462 1721 1465 1728
rect 2902 1722 2905 1728
rect 1462 1718 1678 1721
rect 1862 1718 1870 1721
rect 1874 1718 1894 1721
rect 1986 1718 2078 1721
rect 2330 1718 2334 1721
rect 2346 1718 2358 1721
rect 2450 1718 2750 1721
rect 2754 1718 2798 1721
rect 2802 1718 2830 1721
rect 2834 1718 2854 1721
rect 3002 1718 3022 1721
rect 3166 1721 3169 1728
rect 3030 1718 3161 1721
rect 3166 1718 3478 1721
rect 3494 1721 3497 1728
rect 4278 1722 4281 1728
rect 3494 1718 3502 1721
rect 3510 1718 3694 1721
rect 3770 1718 3838 1721
rect 3850 1718 4046 1721
rect 4098 1718 4174 1721
rect 4290 1718 4310 1721
rect 4450 1718 4566 1721
rect 3030 1712 3033 1718
rect 322 1708 462 1711
rect 1146 1708 1158 1711
rect 1218 1708 1222 1711
rect 1690 1708 1974 1711
rect 2290 1708 2686 1711
rect 2690 1708 2718 1711
rect 2722 1708 2742 1711
rect 2746 1708 2758 1711
rect 2874 1708 2910 1711
rect 3018 1708 3022 1711
rect 3158 1711 3161 1718
rect 3158 1708 3222 1711
rect 3386 1708 3454 1711
rect 3510 1711 3513 1718
rect 3458 1708 3513 1711
rect 3522 1708 3534 1711
rect 3538 1708 3646 1711
rect 3650 1708 3654 1711
rect 3658 1708 3670 1711
rect 3674 1708 3702 1711
rect 3706 1708 3726 1711
rect 3730 1708 3742 1711
rect 3770 1708 3830 1711
rect 3962 1708 3974 1711
rect 4330 1708 4406 1711
rect 1000 1703 1002 1707
rect 1006 1703 1009 1707
rect 1014 1703 1016 1707
rect 2024 1703 2026 1707
rect 2030 1703 2033 1707
rect 2038 1703 2040 1707
rect 3048 1703 3050 1707
rect 3054 1703 3057 1707
rect 3062 1703 3064 1707
rect 4080 1703 4082 1707
rect 4086 1703 4089 1707
rect 4094 1703 4096 1707
rect 122 1698 654 1701
rect 794 1698 798 1701
rect 1138 1698 1654 1701
rect 1658 1698 1662 1701
rect 1706 1698 1982 1701
rect 2058 1698 2278 1701
rect 2282 1698 2358 1701
rect 2386 1698 2481 1701
rect 2490 1698 2582 1701
rect 2586 1698 2638 1701
rect 2642 1698 2806 1701
rect 2898 1698 2966 1701
rect 2978 1698 2982 1701
rect 3010 1698 3038 1701
rect 3146 1698 3166 1701
rect 3186 1698 3230 1701
rect 3234 1698 3358 1701
rect 3402 1698 3422 1701
rect 3442 1698 3550 1701
rect 3594 1698 3766 1701
rect 3770 1698 3814 1701
rect 3882 1698 3950 1701
rect 3954 1698 4054 1701
rect 4186 1698 4198 1701
rect 4242 1698 4246 1701
rect 4370 1698 4462 1701
rect 26 1688 206 1691
rect 278 1688 286 1691
rect 290 1688 350 1691
rect 746 1688 766 1691
rect 866 1688 1014 1691
rect 1018 1688 1158 1691
rect 1178 1688 1222 1691
rect 1234 1688 1286 1691
rect 1314 1688 1326 1691
rect 1346 1688 1534 1691
rect 1538 1688 1694 1691
rect 1818 1688 1894 1691
rect 2050 1688 2142 1691
rect 2154 1688 2166 1691
rect 2170 1688 2177 1691
rect 2182 1688 2262 1691
rect 2306 1688 2430 1691
rect 2434 1688 2438 1691
rect 2478 1691 2481 1698
rect 2478 1688 2518 1691
rect 2634 1688 2678 1691
rect 2730 1688 2790 1691
rect 2830 1688 2838 1691
rect 2854 1688 4182 1691
rect 4186 1688 4238 1691
rect 4242 1688 4334 1691
rect 4338 1688 4414 1691
rect 4418 1688 4502 1691
rect 2182 1682 2185 1688
rect 194 1678 198 1681
rect 234 1678 238 1681
rect 282 1678 286 1681
rect 394 1678 974 1681
rect 1130 1678 1177 1681
rect 1210 1678 1246 1681
rect 1306 1678 1310 1681
rect 1450 1678 1550 1681
rect 1602 1678 1606 1681
rect 1794 1678 1846 1681
rect 1970 1678 1974 1681
rect 1986 1678 2102 1681
rect 2106 1678 2110 1681
rect 2178 1678 2182 1681
rect 2226 1678 2246 1681
rect 2354 1678 2449 1681
rect 2458 1678 2470 1681
rect 2526 1681 2529 1688
rect 2474 1678 2529 1681
rect 2622 1681 2625 1688
rect 2694 1682 2697 1688
rect 2854 1682 2857 1688
rect 2570 1678 2654 1681
rect 2786 1678 2838 1681
rect 2986 1678 3030 1681
rect 3098 1678 3110 1681
rect 3114 1678 3134 1681
rect 3274 1678 3278 1681
rect 3410 1678 3414 1681
rect 3442 1678 3478 1681
rect 3498 1678 3542 1681
rect 3554 1678 3662 1681
rect 3666 1678 3686 1681
rect 3706 1678 3710 1681
rect 3786 1678 3806 1681
rect 3810 1678 3902 1681
rect 3926 1678 4110 1681
rect 4114 1678 4310 1681
rect 4358 1678 4366 1681
rect 4386 1678 4422 1681
rect 4594 1678 4598 1681
rect -26 1671 -22 1672
rect 30 1671 33 1678
rect -26 1668 33 1671
rect 50 1668 158 1671
rect 162 1668 214 1671
rect 218 1668 382 1671
rect 386 1668 438 1671
rect 442 1668 606 1671
rect 1054 1671 1057 1678
rect 1174 1672 1177 1678
rect 1318 1672 1321 1678
rect 1902 1672 1905 1678
rect 970 1668 1057 1671
rect 1242 1668 1254 1671
rect 1258 1668 1286 1671
rect 1362 1668 1598 1671
rect 1610 1668 1702 1671
rect 1706 1668 1750 1671
rect 1754 1668 1798 1671
rect 1834 1668 1878 1671
rect 1882 1668 1902 1671
rect 1938 1668 1950 1671
rect 1954 1668 1990 1671
rect 1994 1668 2094 1671
rect 2098 1668 2310 1671
rect 2314 1668 2382 1671
rect 2386 1668 2398 1671
rect 2402 1668 2422 1671
rect 2446 1671 2449 1678
rect 2918 1672 2921 1678
rect 2926 1672 2929 1678
rect 2934 1672 2937 1678
rect 2446 1668 2454 1671
rect 2458 1668 2486 1671
rect 2522 1668 2590 1671
rect 2626 1668 2630 1671
rect 2674 1668 2710 1671
rect 2946 1668 3078 1671
rect 3190 1671 3193 1678
rect 3926 1672 3929 1678
rect 4358 1672 4361 1678
rect 3186 1668 3193 1671
rect 3202 1668 3206 1671
rect 3210 1668 3246 1671
rect 3362 1668 3398 1671
rect 3482 1668 3630 1671
rect 3682 1668 3686 1671
rect 3706 1668 3710 1671
rect 4074 1668 4094 1671
rect 4154 1668 4198 1671
rect 4418 1668 4446 1671
rect 4458 1668 4494 1671
rect 4530 1668 4582 1671
rect 22 1658 30 1661
rect 34 1658 54 1661
rect 170 1658 198 1661
rect 202 1658 270 1661
rect 306 1658 326 1661
rect 330 1658 334 1661
rect 498 1659 534 1661
rect 494 1658 534 1659
rect 698 1658 718 1661
rect 722 1658 734 1661
rect 754 1658 769 1661
rect 858 1658 878 1661
rect 926 1661 929 1668
rect 1158 1662 1161 1668
rect 926 1658 934 1661
rect 1194 1658 1206 1661
rect 1418 1658 1574 1661
rect 1578 1658 1585 1661
rect 1626 1658 1630 1661
rect 1666 1658 1910 1661
rect 2074 1658 2110 1661
rect 2146 1658 2206 1661
rect 2210 1658 2246 1661
rect 2354 1658 2358 1661
rect 2394 1658 2470 1661
rect 2474 1658 2502 1661
rect 2538 1658 2614 1661
rect 2618 1658 2766 1661
rect 2770 1658 2790 1661
rect 2826 1658 2950 1661
rect 2978 1658 2982 1661
rect 3106 1658 3113 1661
rect 3122 1658 3150 1661
rect 3170 1658 3342 1661
rect 3394 1658 3398 1661
rect 3458 1658 3470 1661
rect 3514 1658 3542 1661
rect 3658 1658 3678 1661
rect 3722 1658 3766 1661
rect 3782 1661 3785 1668
rect 3958 1662 3961 1668
rect 3966 1662 3969 1668
rect 3770 1658 3785 1661
rect 3842 1658 3870 1661
rect 3890 1658 3926 1661
rect 3994 1658 4022 1661
rect 4026 1658 4046 1661
rect 4050 1658 4078 1661
rect 4082 1658 4118 1661
rect 4194 1658 4246 1661
rect 4370 1658 4417 1661
rect 4490 1658 4550 1661
rect 766 1652 769 1658
rect -26 1651 -22 1652
rect -26 1648 6 1651
rect 122 1648 422 1651
rect 426 1648 598 1651
rect 1130 1648 1254 1651
rect 1530 1648 1726 1651
rect 1730 1648 1750 1651
rect 1858 1648 1889 1651
rect 1954 1648 1990 1651
rect 2094 1648 2126 1651
rect 2130 1648 2238 1651
rect 2562 1648 2670 1651
rect 2698 1648 2806 1651
rect 2818 1648 2886 1651
rect 2962 1648 2966 1651
rect 2970 1648 3006 1651
rect 3018 1648 3102 1651
rect 3114 1648 3142 1651
rect 3202 1648 3318 1651
rect 3398 1651 3401 1658
rect 3526 1652 3529 1658
rect 4414 1652 4417 1658
rect 3398 1648 3494 1651
rect 3674 1648 3718 1651
rect 3858 1648 3937 1651
rect 186 1638 246 1641
rect 290 1638 310 1641
rect 326 1638 334 1641
rect 338 1638 366 1641
rect 570 1638 686 1641
rect 706 1638 726 1641
rect 730 1638 838 1641
rect 842 1638 870 1641
rect 1482 1638 1614 1641
rect 1618 1638 1662 1641
rect 1698 1638 1718 1641
rect 1738 1638 1758 1641
rect 1766 1641 1769 1648
rect 1762 1638 1769 1641
rect 1774 1641 1777 1648
rect 1886 1642 1889 1648
rect 2094 1642 2097 1648
rect 3838 1642 3841 1648
rect 3934 1642 3937 1648
rect 3950 1648 3982 1651
rect 4010 1648 4014 1651
rect 4058 1648 4150 1651
rect 4186 1648 4206 1651
rect 4234 1648 4398 1651
rect 4522 1648 4526 1651
rect 3950 1642 3953 1648
rect 1774 1638 1830 1641
rect 1994 1638 2078 1641
rect 2394 1638 3310 1641
rect 3314 1638 3326 1641
rect 3418 1638 3430 1641
rect 3442 1638 3678 1641
rect 3698 1638 3702 1641
rect 4250 1638 4294 1641
rect 4314 1638 4542 1641
rect 98 1628 390 1631
rect 658 1628 1382 1631
rect 2842 1628 2854 1631
rect 2866 1628 2870 1631
rect 3026 1628 3030 1631
rect 3042 1628 3094 1631
rect 3242 1628 3294 1631
rect 3306 1628 3654 1631
rect 4258 1628 4374 1631
rect 170 1618 198 1621
rect 730 1618 1446 1621
rect 1614 1621 1617 1628
rect 1458 1618 1617 1621
rect 1802 1618 2006 1621
rect 2010 1618 2054 1621
rect 2058 1618 2070 1621
rect 2402 1618 2430 1621
rect 2434 1618 2590 1621
rect 2594 1618 2630 1621
rect 2650 1618 2726 1621
rect 2994 1618 3030 1621
rect 3218 1618 3222 1621
rect 3314 1618 3454 1621
rect 3458 1618 3638 1621
rect 3742 1621 3745 1628
rect 3742 1618 4118 1621
rect 4122 1618 4134 1621
rect 4234 1618 4241 1621
rect 4238 1612 4241 1618
rect 194 1608 238 1611
rect 298 1608 398 1611
rect 778 1608 870 1611
rect 898 1608 982 1611
rect 986 1608 1494 1611
rect 1618 1608 1630 1611
rect 1634 1608 1742 1611
rect 2626 1608 2710 1611
rect 3026 1608 3046 1611
rect 4130 1608 4142 1611
rect 496 1603 498 1607
rect 502 1603 505 1607
rect 510 1603 512 1607
rect 1520 1603 1522 1607
rect 1526 1603 1529 1607
rect 1534 1603 1536 1607
rect 1886 1602 1889 1608
rect 2544 1603 2546 1607
rect 2550 1603 2553 1607
rect 2558 1603 2560 1607
rect 3568 1603 3570 1607
rect 3574 1603 3577 1607
rect 3582 1603 3584 1607
rect 762 1598 838 1601
rect 850 1598 910 1601
rect 1066 1598 1142 1601
rect 1346 1598 1366 1601
rect 1610 1598 1638 1601
rect 1914 1598 2150 1601
rect 2282 1598 2286 1601
rect 2466 1598 2502 1601
rect 2506 1598 2518 1601
rect 2658 1598 2766 1601
rect 2898 1598 2902 1601
rect 3034 1598 3046 1601
rect 3242 1598 3502 1601
rect 4010 1598 4142 1601
rect 4242 1598 4510 1601
rect 250 1588 398 1591
rect 434 1588 830 1591
rect 834 1588 958 1591
rect 1122 1588 1134 1591
rect 1138 1588 1702 1591
rect 1722 1588 1750 1591
rect 1754 1588 1926 1591
rect 1994 1588 2238 1591
rect 2250 1588 2390 1591
rect 2442 1588 2494 1591
rect 2542 1588 3190 1591
rect 3194 1588 3270 1591
rect 3394 1588 3510 1591
rect 3514 1588 3982 1591
rect 4082 1588 4254 1591
rect 4258 1588 4366 1591
rect 2542 1582 2545 1588
rect 234 1578 254 1581
rect 354 1578 374 1581
rect 418 1578 510 1581
rect 590 1578 598 1581
rect 614 1578 622 1581
rect 626 1578 742 1581
rect 778 1578 782 1581
rect 986 1578 1078 1581
rect 1370 1578 1409 1581
rect 1730 1578 1862 1581
rect 1874 1578 1886 1581
rect 1954 1578 2006 1581
rect 2010 1578 2294 1581
rect 2298 1578 2366 1581
rect 2370 1578 2542 1581
rect 2714 1578 2774 1581
rect 2834 1578 2846 1581
rect 3090 1578 3150 1581
rect 3154 1578 3310 1581
rect 3446 1578 3454 1581
rect 3458 1578 3574 1581
rect 3578 1578 3630 1581
rect 3722 1578 3926 1581
rect 4074 1578 4150 1581
rect 4282 1578 4294 1581
rect -26 1571 -22 1572
rect 126 1571 129 1578
rect 1406 1572 1409 1578
rect -26 1568 129 1571
rect 378 1568 534 1571
rect 538 1568 878 1571
rect 882 1568 918 1571
rect 930 1568 1326 1571
rect 1362 1568 1374 1571
rect 1538 1568 1550 1571
rect 1674 1568 1790 1571
rect 1834 1568 1966 1571
rect 2082 1568 2134 1571
rect 2138 1568 2526 1571
rect 2666 1568 2734 1571
rect 2738 1568 2822 1571
rect 2842 1568 2846 1571
rect 2930 1568 3070 1571
rect 3178 1568 3190 1571
rect 3354 1568 3494 1571
rect 3506 1568 3630 1571
rect 3690 1568 3894 1571
rect 4018 1568 4022 1571
rect 4166 1571 4169 1578
rect 4166 1568 4198 1571
rect 4226 1568 4230 1571
rect 4238 1571 4241 1578
rect 4238 1568 4326 1571
rect 4394 1568 4398 1571
rect 226 1558 230 1561
rect 242 1558 382 1561
rect 426 1558 438 1561
rect 466 1558 630 1561
rect 1002 1558 1022 1561
rect 1058 1558 1150 1561
rect 1154 1558 1158 1561
rect 1202 1558 1206 1561
rect 1274 1558 1318 1561
rect 1322 1558 1414 1561
rect 1574 1561 1577 1568
rect 1418 1558 1577 1561
rect 1814 1561 1817 1568
rect 2854 1562 2857 1568
rect 1642 1558 1769 1561
rect 1814 1558 1862 1561
rect 1874 1558 1950 1561
rect 1954 1558 2022 1561
rect 2250 1558 2278 1561
rect 2290 1558 2318 1561
rect 2370 1558 2398 1561
rect 2402 1558 2534 1561
rect 2586 1558 2646 1561
rect 2650 1558 2670 1561
rect 2738 1558 2750 1561
rect 2874 1558 2905 1561
rect 2954 1558 3030 1561
rect 3150 1561 3153 1568
rect 3106 1558 3153 1561
rect 3282 1558 3286 1561
rect 3318 1561 3321 1568
rect 3318 1558 3358 1561
rect 3362 1558 4254 1561
rect 4266 1558 4286 1561
rect 4298 1558 4422 1561
rect -26 1551 -22 1552
rect -26 1548 6 1551
rect 162 1548 174 1551
rect 218 1548 262 1551
rect 298 1548 302 1551
rect 394 1548 502 1551
rect 522 1548 542 1551
rect 562 1548 582 1551
rect 618 1548 766 1551
rect 790 1551 793 1558
rect 822 1551 825 1558
rect 1766 1552 1769 1558
rect 790 1548 825 1551
rect 1010 1548 1038 1551
rect 1042 1548 1046 1551
rect 1082 1548 1118 1551
rect 1226 1548 1358 1551
rect 1402 1548 1446 1551
rect 1458 1548 1654 1551
rect 1658 1548 1665 1551
rect 1794 1548 1814 1551
rect 1818 1548 1854 1551
rect 1858 1548 1926 1551
rect 1970 1548 1974 1551
rect 1978 1548 2126 1551
rect 2146 1548 2158 1551
rect 2202 1548 2214 1551
rect 2242 1548 2342 1551
rect 2386 1548 2414 1551
rect 2418 1548 2454 1551
rect 2458 1548 2478 1551
rect 2486 1548 2550 1551
rect 2570 1548 2598 1551
rect 2610 1548 2630 1551
rect 2666 1548 2670 1551
rect 2738 1548 2742 1551
rect 2794 1548 2806 1551
rect 2866 1548 2870 1551
rect 2890 1548 2894 1551
rect 2902 1551 2905 1558
rect 2902 1548 2966 1551
rect 3010 1548 3118 1551
rect 3158 1551 3161 1558
rect 3302 1552 3305 1558
rect 3138 1548 3174 1551
rect 3194 1548 3214 1551
rect 3282 1548 3286 1551
rect 3322 1548 3342 1551
rect 3350 1548 3374 1551
rect 3402 1548 3406 1551
rect 3498 1548 3518 1551
rect 3522 1548 3526 1551
rect 3530 1548 3590 1551
rect 3610 1548 3614 1551
rect 3626 1548 3654 1551
rect 3658 1548 3774 1551
rect 3786 1548 3942 1551
rect 3946 1548 3950 1551
rect 3978 1548 3990 1551
rect 3994 1548 4006 1551
rect 4066 1548 4102 1551
rect 4138 1548 4150 1551
rect 4154 1548 4166 1551
rect 4202 1548 4206 1551
rect 4242 1548 4318 1551
rect 4346 1548 4350 1551
rect 4402 1548 4406 1551
rect 4450 1548 4478 1551
rect 4490 1548 4510 1551
rect 26 1538 374 1541
rect 402 1538 425 1541
rect 442 1538 454 1541
rect 570 1538 590 1541
rect 674 1538 905 1541
rect 994 1538 1046 1541
rect 1054 1541 1057 1548
rect 1050 1538 1086 1541
rect 1214 1541 1217 1548
rect 1194 1538 1294 1541
rect 1402 1538 1486 1541
rect 1522 1538 1718 1541
rect 1750 1541 1753 1548
rect 2350 1542 2353 1548
rect 2486 1542 2489 1548
rect 3350 1542 3353 1548
rect 1730 1538 1766 1541
rect 1842 1538 1846 1541
rect 1874 1538 1878 1541
rect 1914 1538 1958 1541
rect 2034 1538 2078 1541
rect 2082 1538 2118 1541
rect 2202 1538 2230 1541
rect 2234 1538 2262 1541
rect 2274 1538 2278 1541
rect 2282 1538 2294 1541
rect 2394 1538 2398 1541
rect 2506 1538 2518 1541
rect 2578 1538 2590 1541
rect 2626 1538 2638 1541
rect 2642 1538 2894 1541
rect 2914 1538 2918 1541
rect 2978 1538 2998 1541
rect 3066 1538 3110 1541
rect 3146 1538 3222 1541
rect 3226 1538 3246 1541
rect 3298 1538 3326 1541
rect 3434 1538 3446 1541
rect 3474 1538 3534 1541
rect 3538 1538 3553 1541
rect 3570 1538 3622 1541
rect 3634 1538 3702 1541
rect 3850 1538 3862 1541
rect 3954 1538 3966 1541
rect 4046 1541 4049 1548
rect 4182 1542 4185 1548
rect 4230 1542 4233 1548
rect 4002 1538 4102 1541
rect 4258 1538 4278 1541
rect 4298 1538 4302 1541
rect 4370 1538 4470 1541
rect 4474 1538 4486 1541
rect 4538 1538 4561 1541
rect 422 1532 425 1538
rect 806 1532 809 1538
rect 902 1532 905 1538
rect 346 1528 366 1531
rect 458 1528 574 1531
rect 586 1528 718 1531
rect 970 1528 1006 1531
rect 1162 1528 1206 1531
rect 1326 1531 1329 1538
rect 1894 1532 1897 1538
rect 2998 1532 3001 1538
rect 1326 1528 1350 1531
rect 1474 1528 1542 1531
rect 1562 1528 1598 1531
rect 1602 1528 1606 1531
rect 1658 1528 1697 1531
rect 2106 1528 2310 1531
rect 2314 1528 2358 1531
rect 2474 1528 2726 1531
rect 2882 1528 2902 1531
rect 2906 1528 2942 1531
rect 3034 1528 3078 1531
rect 3082 1528 3086 1531
rect 3138 1528 3166 1531
rect 3262 1531 3265 1538
rect 3550 1532 3553 1538
rect 4558 1532 4561 1538
rect 3262 1528 3454 1531
rect 3466 1528 3502 1531
rect 3650 1528 3673 1531
rect 3914 1528 3942 1531
rect 4002 1528 4006 1531
rect 4058 1528 4070 1531
rect 4154 1528 4302 1531
rect 4354 1528 4390 1531
rect 4394 1528 4454 1531
rect 4570 1528 4574 1531
rect 1694 1522 1697 1528
rect 2278 1522 2281 1528
rect 3670 1522 3673 1528
rect 386 1518 470 1521
rect 722 1518 1070 1521
rect 1242 1518 1246 1521
rect 1498 1518 1566 1521
rect 1570 1518 1630 1521
rect 1634 1518 1678 1521
rect 2170 1518 2270 1521
rect 2338 1518 2430 1521
rect 2590 1518 2694 1521
rect 2714 1518 2750 1521
rect 2826 1518 2910 1521
rect 2918 1518 3086 1521
rect 3202 1518 3214 1521
rect 3946 1518 4006 1521
rect 4042 1518 4166 1521
rect 4178 1518 4182 1521
rect 4190 1518 4254 1521
rect 4282 1518 4286 1521
rect 558 1512 561 1518
rect 2590 1512 2593 1518
rect 250 1508 270 1511
rect 330 1508 334 1511
rect 370 1508 486 1511
rect 1026 1508 1054 1511
rect 1058 1508 1606 1511
rect 1698 1508 1710 1511
rect 1714 1508 1782 1511
rect 1906 1508 1982 1511
rect 2050 1508 2174 1511
rect 2194 1508 2198 1511
rect 2218 1508 2246 1511
rect 2290 1508 2302 1511
rect 2330 1508 2334 1511
rect 2394 1508 2502 1511
rect 2674 1508 2766 1511
rect 2918 1511 2921 1518
rect 2778 1508 2921 1511
rect 3114 1508 3334 1511
rect 3370 1508 3374 1511
rect 3418 1508 3790 1511
rect 3810 1508 3998 1511
rect 4002 1508 4062 1511
rect 4190 1511 4193 1518
rect 4130 1508 4193 1511
rect 4202 1508 4278 1511
rect 1000 1503 1002 1507
rect 1006 1503 1009 1507
rect 1014 1503 1016 1507
rect 2024 1503 2026 1507
rect 2030 1503 2033 1507
rect 2038 1503 2040 1507
rect 3048 1503 3050 1507
rect 3054 1503 3057 1507
rect 3062 1503 3064 1507
rect 4080 1503 4082 1507
rect 4086 1503 4089 1507
rect 4094 1503 4096 1507
rect 210 1498 350 1501
rect 1354 1498 1430 1501
rect 1482 1498 1502 1501
rect 1586 1498 1614 1501
rect 1626 1498 1790 1501
rect 1794 1498 1918 1501
rect 2106 1498 2350 1501
rect 2354 1498 2398 1501
rect 2770 1498 2878 1501
rect 3266 1498 3486 1501
rect 3738 1498 3766 1501
rect 3866 1498 3990 1501
rect 4138 1498 4206 1501
rect 4218 1498 4398 1501
rect 566 1492 569 1498
rect 210 1488 222 1491
rect 234 1488 254 1491
rect 354 1488 390 1491
rect 394 1488 430 1491
rect 882 1488 918 1491
rect 922 1488 1334 1491
rect 1386 1488 1438 1491
rect 1442 1488 1622 1491
rect 1650 1488 1702 1491
rect 1714 1488 1742 1491
rect 1778 1488 1918 1491
rect 1930 1488 1990 1491
rect 1994 1488 2054 1491
rect 2058 1488 2206 1491
rect 2242 1488 2414 1491
rect 2442 1488 2862 1491
rect 2874 1488 2878 1491
rect 2882 1488 2982 1491
rect 2994 1488 3038 1491
rect 3042 1488 3054 1491
rect 3058 1488 3142 1491
rect 3178 1488 3206 1491
rect 3250 1488 3382 1491
rect 3386 1488 3398 1491
rect 3402 1488 3406 1491
rect 3706 1488 3750 1491
rect 3770 1488 3774 1491
rect 3778 1488 3830 1491
rect 3834 1488 3878 1491
rect 3882 1488 3902 1491
rect 3906 1488 3918 1491
rect 4122 1488 4238 1491
rect 4266 1488 4294 1491
rect 4298 1488 4550 1491
rect 186 1478 302 1481
rect 306 1478 326 1481
rect 334 1481 337 1488
rect 334 1478 406 1481
rect 410 1478 414 1481
rect 418 1478 430 1481
rect 762 1478 886 1481
rect 906 1478 998 1481
rect 1154 1478 1166 1481
rect 1170 1478 1230 1481
rect 1250 1478 1270 1481
rect 1434 1478 1542 1481
rect 1658 1478 1662 1481
rect 1754 1478 1790 1481
rect 1938 1478 1974 1481
rect 1978 1478 2014 1481
rect 2018 1478 2086 1481
rect 2106 1478 2142 1481
rect 2274 1478 2286 1481
rect 2290 1478 2390 1481
rect 2498 1478 2606 1481
rect 2658 1478 2670 1481
rect 2746 1478 2750 1481
rect 2810 1478 2830 1481
rect 2842 1478 2846 1481
rect 2858 1478 2862 1481
rect 2946 1478 2966 1481
rect 2970 1478 3070 1481
rect 3074 1478 3118 1481
rect 3122 1478 3462 1481
rect 3682 1478 3721 1481
rect 3802 1478 3870 1481
rect 3998 1481 4001 1488
rect 3906 1478 3993 1481
rect 3998 1478 4022 1481
rect 4026 1478 4118 1481
rect 4250 1478 4262 1481
rect 4270 1478 4342 1481
rect -26 1471 -22 1472
rect 30 1471 33 1478
rect -26 1468 33 1471
rect 130 1468 214 1471
rect 242 1468 278 1471
rect 282 1468 297 1471
rect 410 1468 438 1471
rect 550 1471 553 1478
rect 1310 1472 1313 1478
rect 550 1468 622 1471
rect 818 1468 862 1471
rect 1026 1468 1110 1471
rect 1138 1468 1278 1471
rect 1326 1471 1329 1478
rect 1702 1472 1705 1478
rect 1326 1468 1446 1471
rect 1466 1468 1486 1471
rect 1514 1468 1558 1471
rect 1562 1468 1662 1471
rect 1906 1468 1918 1471
rect 1954 1468 1985 1471
rect 2074 1470 2150 1471
rect 2074 1468 2086 1470
rect 162 1458 278 1461
rect 294 1461 297 1468
rect 294 1458 350 1461
rect 534 1458 569 1461
rect 578 1458 598 1461
rect 602 1458 606 1461
rect 610 1458 790 1461
rect 810 1458 902 1461
rect 1002 1458 1038 1461
rect 1042 1458 1078 1461
rect 1094 1458 1102 1461
rect 1154 1458 1174 1461
rect 1194 1458 1206 1461
rect 1266 1458 1302 1461
rect 1322 1458 1350 1461
rect 1378 1458 1470 1461
rect 1538 1458 1566 1461
rect 1714 1458 1726 1461
rect 1766 1461 1769 1468
rect 1766 1458 1814 1461
rect 1882 1458 1958 1461
rect 1982 1461 1985 1468
rect 2090 1468 2150 1470
rect 2174 1471 2177 1478
rect 2174 1468 2206 1471
rect 2226 1468 2254 1471
rect 2322 1468 2337 1471
rect 2346 1468 2446 1471
rect 2466 1468 2470 1471
rect 2562 1468 2590 1471
rect 2610 1468 2902 1471
rect 2994 1468 3046 1471
rect 3058 1468 3062 1471
rect 3090 1468 3094 1471
rect 3114 1468 3126 1471
rect 3202 1468 3206 1471
rect 3234 1468 3238 1471
rect 3242 1468 3254 1471
rect 3322 1468 3518 1471
rect 3522 1468 3566 1471
rect 3614 1471 3617 1478
rect 3718 1472 3721 1478
rect 3990 1472 3993 1478
rect 3614 1468 3630 1471
rect 3650 1468 3654 1471
rect 3738 1468 3774 1471
rect 3778 1468 3782 1471
rect 3786 1468 3846 1471
rect 3914 1468 3982 1471
rect 3994 1468 4038 1471
rect 4066 1468 4110 1471
rect 4146 1468 4166 1471
rect 4234 1468 4238 1471
rect 4270 1471 4273 1478
rect 4382 1472 4385 1478
rect 4258 1468 4273 1471
rect 4338 1468 4374 1471
rect 4402 1468 4438 1471
rect 4466 1468 4486 1471
rect 4494 1471 4497 1478
rect 4494 1468 4542 1471
rect 4554 1468 4558 1471
rect 4578 1468 4582 1471
rect 1982 1458 2086 1461
rect 2090 1458 2102 1461
rect 2146 1458 2150 1461
rect 2162 1458 2190 1461
rect 2218 1458 2262 1461
rect 2266 1458 2326 1461
rect 2334 1461 2337 1468
rect 3302 1462 3305 1468
rect 2334 1458 2358 1461
rect 2394 1458 2502 1461
rect 2530 1458 2694 1461
rect 2706 1458 2710 1461
rect 2810 1458 2862 1461
rect 2882 1458 2886 1461
rect 2914 1458 3110 1461
rect 3114 1458 3118 1461
rect 3130 1458 3190 1461
rect 3194 1458 3206 1461
rect 3210 1458 3246 1461
rect 3250 1458 3273 1461
rect 158 1452 161 1458
rect 534 1452 537 1458
rect 566 1452 569 1458
rect 1622 1452 1625 1458
rect 2462 1452 2465 1458
rect 3270 1452 3273 1458
rect 3346 1458 3350 1461
rect 3394 1458 3398 1461
rect 3450 1458 3606 1461
rect 3618 1458 3670 1461
rect 3698 1458 3702 1461
rect 3714 1458 3726 1461
rect 3802 1458 3814 1461
rect 3818 1458 3878 1461
rect 3922 1458 3942 1461
rect 3970 1458 3974 1461
rect 4010 1458 4014 1461
rect 4026 1458 4030 1461
rect 4158 1458 4174 1461
rect 4242 1458 4246 1461
rect 4266 1458 4270 1461
rect 4314 1458 4318 1461
rect 4338 1458 4342 1461
rect 4378 1458 4414 1461
rect 4418 1458 4470 1461
rect 4474 1458 4502 1461
rect 4546 1458 4582 1461
rect 3278 1452 3281 1458
rect 3742 1452 3745 1458
rect -26 1451 -22 1452
rect -26 1448 6 1451
rect 262 1448 286 1451
rect 290 1448 358 1451
rect 602 1448 617 1451
rect 906 1448 926 1451
rect 934 1448 958 1451
rect 982 1448 990 1451
rect 994 1448 1046 1451
rect 1050 1448 1094 1451
rect 1178 1448 1190 1451
rect 1306 1448 1326 1451
rect 1682 1448 1830 1451
rect 1866 1448 1982 1451
rect 1986 1448 1990 1451
rect 2034 1448 2222 1451
rect 2266 1448 2310 1451
rect 2342 1448 2350 1451
rect 2482 1448 2486 1451
rect 2666 1448 2670 1451
rect 2690 1448 2806 1451
rect 2842 1448 2894 1451
rect 2898 1448 3006 1451
rect 3082 1448 3094 1451
rect 3198 1448 3225 1451
rect 3354 1448 3446 1451
rect 3498 1448 3510 1451
rect 3586 1448 3614 1451
rect 3958 1451 3961 1458
rect 4150 1452 4153 1458
rect 4158 1452 4161 1458
rect 3874 1448 3961 1451
rect 3994 1448 4006 1451
rect 4130 1448 4134 1451
rect 4170 1448 4294 1451
rect 4298 1448 4382 1451
rect 4410 1448 4422 1451
rect 4434 1448 4478 1451
rect 4514 1448 4550 1451
rect 262 1442 265 1448
rect 614 1442 617 1448
rect 934 1442 937 1448
rect 2342 1442 2345 1448
rect 3198 1442 3201 1448
rect 3222 1442 3225 1448
rect 4174 1442 4177 1448
rect 298 1438 446 1441
rect 450 1438 550 1441
rect 562 1438 566 1441
rect 986 1438 1038 1441
rect 1042 1438 1070 1441
rect 1202 1438 1262 1441
rect 1266 1438 1574 1441
rect 1706 1438 1798 1441
rect 1874 1438 1886 1441
rect 1978 1438 2030 1441
rect 2194 1438 2198 1441
rect 2210 1438 2230 1441
rect 2426 1438 2638 1441
rect 2674 1438 2726 1441
rect 2754 1438 2782 1441
rect 2830 1438 2849 1441
rect 2882 1438 2950 1441
rect 2954 1438 2966 1441
rect 2978 1438 2993 1441
rect 3082 1438 3086 1441
rect 3290 1438 3670 1441
rect 3674 1438 3998 1441
rect 4190 1438 4225 1441
rect 4338 1438 4358 1441
rect 4458 1438 4510 1441
rect 4562 1438 4566 1441
rect 1646 1432 1649 1438
rect 226 1428 334 1431
rect 466 1428 662 1431
rect 946 1428 1134 1431
rect 1290 1428 1638 1431
rect 1882 1428 2126 1431
rect 2406 1431 2409 1438
rect 2830 1432 2833 1438
rect 2846 1432 2849 1438
rect 2990 1432 2993 1438
rect 4190 1432 4193 1438
rect 4222 1432 4225 1438
rect 2130 1428 2630 1431
rect 2634 1428 2654 1431
rect 2706 1428 2774 1431
rect 3146 1428 3214 1431
rect 3418 1428 3750 1431
rect 3754 1428 4062 1431
rect 4498 1428 4550 1431
rect 482 1418 830 1421
rect 1314 1418 1318 1421
rect 1418 1418 1486 1421
rect 1490 1418 1550 1421
rect 1554 1418 1598 1421
rect 1602 1418 1646 1421
rect 1962 1418 2246 1421
rect 2250 1418 2358 1421
rect 2362 1418 2382 1421
rect 2386 1418 2694 1421
rect 2778 1418 2814 1421
rect 3130 1418 3161 1421
rect 3170 1418 3454 1421
rect 3554 1418 3614 1421
rect 3618 1418 3774 1421
rect 3786 1418 3814 1421
rect 4290 1418 4326 1421
rect 3158 1412 3161 1418
rect 4230 1412 4233 1418
rect 66 1408 262 1411
rect 1218 1408 1222 1411
rect 1226 1408 1270 1411
rect 1274 1408 1414 1411
rect 1874 1408 1958 1411
rect 2170 1408 2278 1411
rect 2370 1408 2438 1411
rect 2450 1408 2534 1411
rect 2650 1408 2790 1411
rect 2810 1408 2846 1411
rect 3210 1408 3238 1411
rect 3242 1408 3326 1411
rect 3346 1408 3518 1411
rect 3818 1408 4182 1411
rect 4466 1408 4478 1411
rect 496 1403 498 1407
rect 502 1403 505 1407
rect 510 1403 512 1407
rect 1520 1403 1522 1407
rect 1526 1403 1529 1407
rect 1534 1403 1536 1407
rect 2544 1403 2546 1407
rect 2550 1403 2553 1407
rect 2558 1403 2560 1407
rect 3568 1403 3570 1407
rect 3574 1403 3577 1407
rect 3582 1403 3584 1407
rect 74 1398 438 1401
rect 1770 1398 2102 1401
rect 2106 1398 2454 1401
rect 2458 1398 2486 1401
rect 2674 1398 2934 1401
rect 3154 1398 3430 1401
rect 3442 1398 3470 1401
rect 3786 1398 4158 1401
rect 4162 1398 4190 1401
rect 4202 1398 4254 1401
rect -26 1391 -22 1392
rect -26 1388 57 1391
rect 154 1388 190 1391
rect 194 1388 262 1391
rect 266 1388 462 1391
rect 898 1388 966 1391
rect 970 1388 1014 1391
rect 1018 1388 1142 1391
rect 1290 1388 1510 1391
rect 1722 1388 1798 1391
rect 1882 1388 1902 1391
rect 2174 1388 2182 1391
rect 2186 1388 2206 1391
rect 2214 1388 2430 1391
rect 2490 1388 2574 1391
rect 2602 1388 2638 1391
rect 2650 1388 2894 1391
rect 3114 1388 3166 1391
rect 3218 1388 3366 1391
rect 3370 1388 3486 1391
rect 3506 1388 3926 1391
rect 3946 1388 4054 1391
rect 4098 1388 4174 1391
rect 4178 1388 4190 1391
rect 4230 1388 4238 1391
rect 4242 1388 4246 1391
rect 4290 1388 4302 1391
rect 4306 1388 4518 1391
rect 54 1382 57 1388
rect 2214 1382 2217 1388
rect -26 1378 38 1381
rect 146 1378 390 1381
rect 598 1378 606 1381
rect 610 1378 718 1381
rect 930 1378 950 1381
rect 1146 1378 1590 1381
rect 1594 1378 1678 1381
rect 1746 1378 1814 1381
rect 1818 1378 2110 1381
rect 2114 1378 2214 1381
rect 2298 1378 2350 1381
rect 2354 1378 2478 1381
rect 2522 1378 2526 1381
rect 2530 1378 2542 1381
rect 2546 1378 2606 1381
rect 2730 1378 2734 1381
rect 2770 1378 2790 1381
rect 2826 1378 2862 1381
rect 2874 1378 2926 1381
rect 3066 1378 3086 1381
rect 3122 1378 3134 1381
rect 3198 1381 3201 1388
rect 4574 1382 4577 1388
rect 3170 1378 3262 1381
rect 3282 1378 3374 1381
rect 3474 1378 3566 1381
rect 3570 1378 3590 1381
rect 3594 1378 3670 1381
rect 3674 1378 3678 1381
rect 3682 1378 3710 1381
rect 3866 1378 3910 1381
rect 3930 1378 4390 1381
rect 4394 1378 4446 1381
rect -26 1372 -23 1378
rect -26 1368 -22 1372
rect 26 1368 86 1371
rect 322 1368 350 1371
rect 394 1368 782 1371
rect 906 1368 910 1371
rect 914 1368 974 1371
rect 1106 1368 1166 1371
rect 1234 1368 1246 1371
rect 1394 1368 1462 1371
rect 1466 1368 1470 1371
rect 1498 1368 1502 1371
rect 1554 1368 1598 1371
rect 1602 1368 1726 1371
rect 1866 1368 1870 1371
rect 1898 1368 1918 1371
rect 1994 1368 2014 1371
rect 2202 1368 2494 1371
rect 2594 1368 2614 1371
rect 2634 1368 2862 1371
rect 2866 1368 2966 1371
rect 2978 1368 3358 1371
rect 3378 1368 3430 1371
rect 3434 1368 3614 1371
rect 3730 1368 3758 1371
rect 3770 1368 3782 1371
rect 3874 1368 3974 1371
rect 3978 1368 4182 1371
rect 4222 1368 4246 1371
rect 4250 1368 4294 1371
rect 4298 1368 4334 1371
rect 4530 1368 4577 1371
rect 50 1358 174 1361
rect 178 1358 278 1361
rect 442 1358 478 1361
rect 778 1358 782 1361
rect 786 1358 846 1361
rect 954 1358 1022 1361
rect 1038 1361 1041 1368
rect 1038 1358 1054 1361
rect 1082 1358 1110 1361
rect 1162 1358 1174 1361
rect 1178 1358 1206 1361
rect 1250 1358 1254 1361
rect 1266 1358 1334 1361
rect 1382 1361 1385 1368
rect 1370 1358 1454 1361
rect 1482 1358 1542 1361
rect 1546 1358 1590 1361
rect 1594 1358 1758 1361
rect 1778 1358 1790 1361
rect 2070 1361 2073 1368
rect 1818 1358 2142 1361
rect 2146 1358 2182 1361
rect 2282 1358 2286 1361
rect 2306 1358 2342 1361
rect 2346 1358 2366 1361
rect 2386 1358 2390 1361
rect 2394 1358 2422 1361
rect 2434 1358 2462 1361
rect 2494 1361 2497 1368
rect 2494 1358 2526 1361
rect 2642 1358 2665 1361
rect 2738 1358 2742 1361
rect 2770 1358 2894 1361
rect 2946 1358 3126 1361
rect 3138 1358 3174 1361
rect 3178 1358 3185 1361
rect 3190 1358 3502 1361
rect 3538 1358 3582 1361
rect 3602 1358 3838 1361
rect 3842 1358 3878 1361
rect 3898 1358 3998 1361
rect 4002 1358 4006 1361
rect 4018 1358 4134 1361
rect 4222 1361 4225 1368
rect 4138 1358 4225 1361
rect 4234 1358 4270 1361
rect 4374 1361 4377 1368
rect 4354 1358 4406 1361
rect 4410 1358 4486 1361
rect 4494 1361 4497 1368
rect 4574 1362 4577 1368
rect 4494 1358 4518 1361
rect -26 1351 -22 1352
rect -26 1348 6 1351
rect 46 1348 54 1351
rect 58 1348 230 1351
rect 386 1348 574 1351
rect 678 1351 681 1358
rect 710 1351 713 1358
rect 2662 1352 2665 1358
rect 3190 1352 3193 1358
rect 678 1348 713 1351
rect 762 1348 766 1351
rect 1066 1348 1134 1351
rect 1162 1348 1174 1351
rect 1210 1348 1238 1351
rect 1494 1348 1502 1351
rect 1674 1348 1702 1351
rect 1746 1348 1758 1351
rect 1794 1348 1814 1351
rect 1850 1348 1886 1351
rect 1946 1348 2134 1351
rect 2138 1348 2150 1351
rect 2266 1348 2358 1351
rect 2402 1348 2414 1351
rect 2458 1348 2462 1351
rect 2498 1348 2510 1351
rect 2642 1348 2646 1351
rect 2754 1348 2782 1351
rect 2786 1348 2902 1351
rect 2954 1348 2974 1351
rect 3010 1348 3038 1351
rect 3066 1348 3070 1351
rect 3122 1348 3150 1351
rect 3186 1348 3190 1351
rect 3210 1348 3262 1351
rect 3386 1348 3422 1351
rect 3466 1348 3510 1351
rect 3530 1348 3558 1351
rect 3602 1348 3630 1351
rect 3738 1348 3830 1351
rect 3866 1348 3942 1351
rect 3994 1348 4022 1351
rect 4026 1348 4030 1351
rect 4058 1348 4166 1351
rect 4242 1348 4278 1351
rect 4322 1348 4470 1351
rect 4498 1348 4502 1351
rect 4562 1348 4566 1351
rect 310 1341 313 1348
rect 310 1338 470 1341
rect 498 1338 542 1341
rect 546 1338 558 1341
rect 562 1338 598 1341
rect 838 1341 841 1348
rect 694 1338 841 1341
rect 846 1341 849 1348
rect 846 1338 942 1341
rect 1002 1338 1038 1341
rect 1090 1338 1126 1341
rect 1290 1338 1310 1341
rect 1358 1341 1361 1348
rect 1494 1342 1497 1348
rect 3038 1342 3041 1348
rect 3334 1342 3337 1348
rect 1358 1338 1398 1341
rect 1418 1338 1462 1341
rect 1546 1338 1558 1341
rect 1634 1338 2134 1341
rect 2146 1338 2198 1341
rect 2318 1338 2366 1341
rect 2394 1338 2406 1341
rect 2474 1338 2598 1341
rect 2618 1338 2710 1341
rect 2722 1338 2934 1341
rect 3050 1338 3078 1341
rect 3282 1338 3286 1341
rect 3530 1338 3670 1341
rect 3674 1338 3734 1341
rect 3738 1338 3750 1341
rect 3778 1338 3854 1341
rect 3970 1338 4030 1341
rect 4046 1341 4049 1348
rect 4046 1338 4126 1341
rect 4218 1338 4230 1341
rect 4282 1338 4318 1341
rect 4434 1338 4454 1341
rect 4514 1338 4598 1341
rect 694 1332 697 1338
rect 2262 1332 2265 1338
rect 2318 1332 2321 1338
rect 2950 1332 2953 1338
rect 162 1328 326 1331
rect 562 1328 566 1331
rect 570 1328 606 1331
rect 842 1328 926 1331
rect 930 1328 942 1331
rect 1074 1328 1094 1331
rect 1122 1328 1158 1331
rect 1194 1328 1230 1331
rect 1234 1328 1310 1331
rect 1426 1328 1462 1331
rect 1562 1328 1566 1331
rect 1586 1328 1590 1331
rect 1666 1328 1694 1331
rect 1778 1328 1830 1331
rect 1890 1328 1934 1331
rect 1970 1328 1974 1331
rect 1978 1328 2006 1331
rect 2066 1328 2070 1331
rect 2074 1328 2214 1331
rect 2362 1328 2446 1331
rect 2458 1328 2510 1331
rect 2530 1328 2566 1331
rect 2666 1328 2670 1331
rect 2778 1328 2822 1331
rect 2842 1328 2846 1331
rect 2858 1328 2910 1331
rect 2930 1328 2934 1331
rect 3010 1328 3110 1331
rect 3114 1328 3126 1331
rect 3130 1328 3166 1331
rect 3294 1331 3297 1338
rect 3226 1328 3297 1331
rect 3314 1328 3526 1331
rect 3546 1328 3598 1331
rect 3618 1328 3697 1331
rect 3706 1328 3758 1331
rect 3762 1328 3782 1331
rect 3910 1331 3913 1338
rect 4342 1332 4345 1338
rect 3910 1328 3950 1331
rect 3962 1328 3966 1331
rect 3970 1328 4094 1331
rect 4098 1328 4150 1331
rect 4154 1328 4174 1331
rect 4178 1328 4206 1331
rect 4282 1328 4326 1331
rect 4402 1328 4582 1331
rect 218 1318 246 1321
rect 298 1318 358 1321
rect 442 1318 582 1321
rect 754 1318 862 1321
rect 1070 1321 1073 1328
rect 946 1318 1073 1321
rect 1106 1318 1254 1321
rect 1258 1318 1310 1321
rect 1606 1321 1609 1328
rect 1522 1318 1609 1321
rect 1846 1321 1849 1328
rect 1846 1318 1886 1321
rect 1906 1318 1918 1321
rect 1950 1321 1953 1328
rect 2646 1322 2649 1328
rect 3206 1322 3209 1328
rect 3694 1322 3697 1328
rect 1930 1318 1953 1321
rect 1994 1318 2006 1321
rect 2010 1318 2046 1321
rect 2050 1318 2150 1321
rect 2266 1318 2326 1321
rect 2682 1318 2726 1321
rect 2818 1318 3166 1321
rect 3170 1318 3174 1321
rect 3226 1318 3230 1321
rect 3282 1318 3318 1321
rect 3322 1318 3430 1321
rect 3486 1318 3558 1321
rect 3562 1318 3590 1321
rect 3610 1318 3638 1321
rect 3642 1318 3649 1321
rect 3722 1318 3798 1321
rect 3834 1318 3966 1321
rect 4018 1318 4046 1321
rect 4138 1318 4214 1321
rect 4234 1318 4278 1321
rect 4398 1321 4401 1328
rect 4282 1318 4401 1321
rect 1086 1312 1089 1318
rect 266 1308 302 1311
rect 370 1308 614 1311
rect 618 1308 654 1311
rect 818 1308 862 1311
rect 1402 1308 1406 1311
rect 1450 1308 1702 1311
rect 1730 1308 1750 1311
rect 1754 1308 1942 1311
rect 2370 1308 2438 1311
rect 2442 1308 2510 1311
rect 2650 1308 2702 1311
rect 2770 1308 2798 1311
rect 2834 1308 2838 1311
rect 2858 1308 2862 1311
rect 2890 1308 3038 1311
rect 3082 1308 3190 1311
rect 3298 1308 3334 1311
rect 3486 1311 3489 1318
rect 3338 1308 3489 1311
rect 3506 1308 3534 1311
rect 3538 1308 3590 1311
rect 3594 1308 3630 1311
rect 3634 1308 3686 1311
rect 3698 1308 3702 1311
rect 3802 1308 3942 1311
rect 3954 1308 4038 1311
rect 4042 1308 4062 1311
rect 4146 1308 4326 1311
rect 4362 1308 4366 1311
rect 1000 1303 1002 1307
rect 1006 1303 1009 1307
rect 1014 1303 1016 1307
rect 2024 1303 2026 1307
rect 2030 1303 2033 1307
rect 2038 1303 2040 1307
rect 26 1298 622 1301
rect 850 1298 894 1301
rect 898 1298 958 1301
rect 1026 1298 1046 1301
rect 1050 1298 1214 1301
rect 1226 1298 1238 1301
rect 1258 1298 1374 1301
rect 1378 1298 1414 1301
rect 1426 1298 1454 1301
rect 1458 1298 1582 1301
rect 1698 1298 1958 1301
rect 2250 1298 2262 1301
rect 2510 1301 2513 1308
rect 3048 1303 3050 1307
rect 3054 1303 3057 1307
rect 3062 1303 3064 1307
rect 4080 1303 4082 1307
rect 4086 1303 4089 1307
rect 4094 1303 4096 1307
rect 2510 1298 2870 1301
rect 2922 1298 2926 1301
rect 2978 1298 3006 1301
rect 3098 1298 3110 1301
rect 3130 1298 3142 1301
rect 3250 1298 3398 1301
rect 3410 1298 3486 1301
rect 3522 1298 3606 1301
rect 3682 1298 3686 1301
rect 3786 1298 3798 1301
rect 3850 1298 3870 1301
rect 3914 1298 3998 1301
rect 4170 1298 4278 1301
rect 4338 1298 4478 1301
rect 554 1288 590 1291
rect 594 1288 734 1291
rect 874 1288 990 1291
rect 1130 1288 1486 1291
rect 1658 1288 1678 1291
rect 1822 1288 1830 1291
rect 1834 1288 1862 1291
rect 1906 1288 1966 1291
rect 2106 1288 2126 1291
rect 2130 1288 2142 1291
rect 2346 1288 2446 1291
rect 2450 1288 2622 1291
rect 2630 1288 2638 1291
rect 2642 1288 2662 1291
rect 2674 1288 2678 1291
rect 2690 1288 2718 1291
rect 2754 1288 2766 1291
rect 2802 1288 2870 1291
rect 2874 1288 2942 1291
rect 2954 1288 2966 1291
rect 3010 1288 3134 1291
rect 3162 1288 3174 1291
rect 3242 1288 3294 1291
rect 3370 1288 3398 1291
rect 3402 1288 3422 1291
rect 3426 1288 3446 1291
rect 3622 1291 3625 1298
rect 3670 1292 3673 1298
rect 3482 1288 3654 1291
rect 3658 1288 3662 1291
rect 3690 1288 3718 1291
rect 3738 1288 3782 1291
rect 3842 1288 4118 1291
rect 4122 1288 4238 1291
rect 4242 1288 4254 1291
rect 4318 1291 4321 1298
rect 4318 1288 4406 1291
rect 194 1278 206 1281
rect 234 1278 270 1281
rect 282 1278 318 1281
rect 322 1278 358 1281
rect 426 1278 430 1281
rect 434 1278 478 1281
rect 794 1278 854 1281
rect 858 1278 910 1281
rect 1110 1281 1113 1288
rect 1090 1278 1113 1281
rect 1118 1281 1121 1288
rect 1118 1278 1198 1281
rect 1306 1278 1382 1281
rect 1410 1278 1414 1281
rect 1562 1278 1574 1281
rect 1618 1278 1630 1281
rect 1870 1281 1873 1288
rect 4590 1282 4593 1288
rect 1826 1278 1873 1281
rect 1882 1278 1886 1281
rect 1914 1278 1950 1281
rect 1978 1278 2110 1281
rect 2170 1278 2190 1281
rect 2218 1278 2246 1281
rect 2258 1278 2382 1281
rect 2386 1278 2494 1281
rect 2498 1278 2518 1281
rect 2618 1278 2678 1281
rect 2722 1278 2838 1281
rect 2842 1278 3030 1281
rect 3034 1278 3350 1281
rect 3354 1278 3590 1281
rect 3610 1278 3630 1281
rect 3634 1278 3742 1281
rect 3754 1278 3774 1281
rect 3802 1278 3822 1281
rect 3882 1278 3942 1281
rect 3962 1278 4014 1281
rect 4034 1278 4158 1281
rect 4162 1278 4350 1281
rect 4378 1278 4494 1281
rect 4522 1278 4534 1281
rect -26 1271 -22 1272
rect 30 1271 33 1278
rect -26 1268 33 1271
rect 162 1268 182 1271
rect 186 1268 230 1271
rect 258 1268 302 1271
rect 306 1268 334 1271
rect 370 1268 374 1271
rect 474 1268 558 1271
rect 590 1271 593 1278
rect 562 1268 593 1271
rect 702 1268 721 1271
rect 906 1268 910 1271
rect 950 1268 1086 1271
rect 1178 1268 1182 1271
rect 1210 1268 1398 1271
rect 1402 1268 1454 1271
rect 1466 1268 1638 1271
rect 1842 1268 1870 1271
rect 1898 1268 1902 1271
rect 1930 1268 1974 1271
rect 2034 1268 2054 1271
rect 2106 1268 2110 1271
rect 2118 1271 2121 1278
rect 2118 1268 2150 1271
rect 2218 1268 2230 1271
rect 2238 1270 2358 1271
rect 230 1262 233 1268
rect 702 1262 705 1268
rect 718 1262 721 1268
rect 950 1262 953 1268
rect 1206 1262 1209 1268
rect 2242 1268 2358 1270
rect 2362 1268 2390 1271
rect 2490 1268 2518 1271
rect 2546 1268 2550 1271
rect 2618 1268 2622 1271
rect 2730 1268 2734 1271
rect 2746 1268 2774 1271
rect 2786 1268 2902 1271
rect 2906 1268 2937 1271
rect 2962 1268 3014 1271
rect 3034 1268 3174 1271
rect 3234 1268 3238 1271
rect 3274 1268 3278 1271
rect 3306 1268 3310 1271
rect 3322 1268 3462 1271
rect 3466 1268 3486 1271
rect 3538 1268 3566 1271
rect 3610 1268 3622 1271
rect 3658 1268 3838 1271
rect 3874 1268 3950 1271
rect 3954 1268 3974 1271
rect 4034 1268 4062 1271
rect 4090 1268 4094 1271
rect 4138 1268 4150 1271
rect 4178 1268 4438 1271
rect 4466 1268 4486 1271
rect 4518 1268 4550 1271
rect 170 1258 190 1261
rect 194 1258 214 1261
rect 290 1258 302 1261
rect 330 1258 414 1261
rect 450 1258 486 1261
rect 1146 1258 1158 1261
rect 1290 1258 1534 1261
rect 1546 1258 1614 1261
rect 1618 1258 1625 1261
rect 1666 1258 1670 1261
rect 1706 1258 1718 1261
rect 1730 1258 1734 1261
rect 1746 1258 1750 1261
rect 1754 1258 1798 1261
rect 1866 1258 1910 1261
rect 1914 1258 1934 1261
rect 1938 1258 1990 1261
rect 2098 1258 2102 1261
rect 2122 1258 2150 1261
rect 2194 1258 2198 1261
rect 2290 1258 2318 1261
rect 2378 1258 2390 1261
rect 2466 1258 2494 1261
rect 2514 1258 2534 1261
rect 2658 1258 2662 1261
rect 2714 1258 2734 1261
rect 2738 1258 2798 1261
rect 2858 1258 2886 1261
rect 2898 1258 2902 1261
rect 2914 1258 2918 1261
rect 2934 1261 2937 1268
rect 2934 1258 2974 1261
rect 2994 1258 3038 1261
rect 3042 1258 3118 1261
rect 3146 1258 3150 1261
rect 3178 1258 3366 1261
rect 3394 1258 3398 1261
rect 3482 1258 3534 1261
rect 3538 1258 3545 1261
rect 3554 1258 3646 1261
rect 3674 1258 3678 1261
rect 3698 1258 3702 1261
rect 3762 1258 3774 1261
rect 3778 1258 3878 1261
rect 3890 1258 3918 1261
rect 3938 1258 3966 1261
rect 3986 1258 4049 1261
rect 4058 1258 4078 1261
rect 4082 1258 4110 1261
rect 4114 1258 4166 1261
rect 4258 1258 4262 1261
rect 4266 1258 4318 1261
rect 4362 1258 4366 1261
rect 4378 1258 4390 1261
rect 4518 1261 4521 1268
rect 4422 1258 4521 1261
rect 4554 1258 4558 1261
rect 446 1252 449 1258
rect 542 1252 545 1258
rect -26 1251 -22 1252
rect -26 1248 6 1251
rect 274 1248 342 1251
rect 602 1248 750 1251
rect 922 1248 1038 1251
rect 1058 1248 1222 1251
rect 1234 1248 1310 1251
rect 1362 1248 1366 1251
rect 1378 1248 1382 1251
rect 1402 1248 1470 1251
rect 1490 1248 1510 1251
rect 1594 1248 1606 1251
rect 1618 1248 1630 1251
rect 1650 1248 1654 1251
rect 1754 1248 1806 1251
rect 1842 1248 1918 1251
rect 1990 1251 1993 1258
rect 1990 1248 2022 1251
rect 2026 1248 2070 1251
rect 2230 1251 2233 1258
rect 2846 1252 2849 1258
rect 2926 1252 2929 1258
rect 2094 1248 2201 1251
rect 2230 1248 2238 1251
rect 2274 1248 2278 1251
rect 2314 1248 2318 1251
rect 2322 1248 2342 1251
rect 2378 1248 2422 1251
rect 2586 1248 2614 1251
rect 2706 1248 2710 1251
rect 2754 1248 2774 1251
rect 2786 1248 2814 1251
rect 2890 1248 2894 1251
rect 2942 1248 3054 1251
rect 3066 1248 3070 1251
rect 3082 1248 3094 1251
rect 3106 1248 3110 1251
rect 3146 1248 3158 1251
rect 3274 1248 3318 1251
rect 3406 1251 3409 1258
rect 3322 1248 3409 1251
rect 3470 1252 3473 1258
rect 4046 1252 4049 1258
rect 3482 1248 3486 1251
rect 3506 1248 3510 1251
rect 3554 1248 3566 1251
rect 3602 1248 3846 1251
rect 3922 1248 3966 1251
rect 4058 1248 4062 1251
rect 4106 1248 4142 1251
rect 4182 1251 4185 1258
rect 4422 1252 4425 1258
rect 4182 1248 4278 1251
rect 4298 1248 4302 1251
rect 4306 1248 4382 1251
rect 4514 1248 4518 1251
rect 586 1238 606 1241
rect 878 1241 881 1248
rect 2094 1242 2097 1248
rect 2198 1242 2201 1248
rect 878 1238 1022 1241
rect 1026 1238 1062 1241
rect 1154 1238 1182 1241
rect 1330 1238 1446 1241
rect 1530 1238 1590 1241
rect 1610 1238 1630 1241
rect 1714 1238 1897 1241
rect 1914 1238 1982 1241
rect 2422 1241 2425 1248
rect 2574 1242 2577 1248
rect 2862 1242 2865 1248
rect 2942 1242 2945 1248
rect 4462 1242 4465 1248
rect 2422 1238 2526 1241
rect 2530 1238 2558 1241
rect 2618 1238 2654 1241
rect 2690 1238 2830 1241
rect 2842 1238 2846 1241
rect 2954 1238 2998 1241
rect 3042 1238 3230 1241
rect 3234 1238 3366 1241
rect 3370 1238 3902 1241
rect 3962 1238 3990 1241
rect 4026 1238 4078 1241
rect 4170 1238 4406 1241
rect 4494 1241 4497 1248
rect 4494 1238 4542 1241
rect 1894 1232 1897 1238
rect 242 1228 510 1231
rect 682 1228 1246 1231
rect 1442 1228 1462 1231
rect 1482 1228 1614 1231
rect 1738 1228 1838 1231
rect 1930 1228 2222 1231
rect 2394 1228 2446 1231
rect 2642 1228 2734 1231
rect 2738 1228 2886 1231
rect 2922 1228 3030 1231
rect 3058 1228 3222 1231
rect 3258 1228 3318 1231
rect 3322 1228 3414 1231
rect 3426 1228 3430 1231
rect 3442 1228 3534 1231
rect 3546 1228 3625 1231
rect 3650 1228 3806 1231
rect 3890 1228 4046 1231
rect 4130 1228 4177 1231
rect 4194 1228 4206 1231
rect 4242 1228 4286 1231
rect 4290 1228 4334 1231
rect 4338 1228 4374 1231
rect 338 1218 806 1221
rect 986 1218 1286 1221
rect 1298 1218 1545 1221
rect 1666 1218 1798 1221
rect 1858 1218 1886 1221
rect 1926 1221 1929 1228
rect 3622 1222 3625 1228
rect 4174 1222 4177 1228
rect 1890 1218 1929 1221
rect 1954 1218 2006 1221
rect 2010 1218 2454 1221
rect 2522 1218 2702 1221
rect 2770 1218 2806 1221
rect 2810 1218 2894 1221
rect 2914 1218 2958 1221
rect 3010 1218 3094 1221
rect 3178 1218 3510 1221
rect 3634 1218 3726 1221
rect 3746 1218 3926 1221
rect 4026 1218 4169 1221
rect 4214 1221 4217 1228
rect 4202 1218 4217 1221
rect 4306 1218 4390 1221
rect 4402 1218 4502 1221
rect 578 1208 710 1211
rect 810 1208 1142 1211
rect 1298 1208 1502 1211
rect 1542 1211 1545 1218
rect 1542 1208 1678 1211
rect 1698 1208 1742 1211
rect 1978 1208 2110 1211
rect 2138 1208 2238 1211
rect 2242 1208 2302 1211
rect 2314 1208 2318 1211
rect 2698 1208 2710 1211
rect 2714 1208 2990 1211
rect 2994 1208 3366 1211
rect 3626 1208 3646 1211
rect 3658 1208 3678 1211
rect 3754 1208 3862 1211
rect 3970 1208 3974 1211
rect 4066 1208 4070 1211
rect 4166 1211 4169 1218
rect 4166 1208 4214 1211
rect 4330 1208 4510 1211
rect 496 1203 498 1207
rect 502 1203 505 1207
rect 510 1203 512 1207
rect 1520 1203 1522 1207
rect 1526 1203 1529 1207
rect 1534 1203 1536 1207
rect 2544 1203 2546 1207
rect 2550 1203 2553 1207
rect 2558 1203 2560 1207
rect 3568 1203 3570 1207
rect 3574 1203 3577 1207
rect 3582 1203 3584 1207
rect 4142 1202 4145 1208
rect 346 1198 446 1201
rect 546 1198 734 1201
rect 1098 1198 1118 1201
rect 1330 1198 1494 1201
rect 1722 1198 1926 1201
rect 1934 1198 2046 1201
rect 2194 1198 2262 1201
rect 2266 1198 2310 1201
rect 2338 1198 2438 1201
rect 2730 1198 2742 1201
rect 2794 1198 2982 1201
rect 3154 1198 3166 1201
rect 3218 1198 3294 1201
rect 3346 1198 3350 1201
rect 3362 1198 3398 1201
rect 3458 1198 3542 1201
rect 3618 1198 3654 1201
rect 3674 1198 4046 1201
rect 4154 1198 4294 1201
rect 4298 1198 4398 1201
rect 1198 1192 1201 1198
rect -26 1191 -22 1192
rect -26 1188 33 1191
rect 122 1188 334 1191
rect 410 1188 566 1191
rect 1370 1188 1430 1191
rect 1434 1188 1598 1191
rect 1602 1188 1686 1191
rect 1934 1191 1937 1198
rect 3014 1192 3017 1198
rect 1890 1188 1937 1191
rect 1946 1188 1990 1191
rect 2018 1188 2182 1191
rect 2186 1188 2214 1191
rect 2282 1188 2318 1191
rect 2418 1188 2462 1191
rect 2498 1188 2798 1191
rect 2834 1188 2878 1191
rect 2882 1188 2910 1191
rect 2970 1188 3006 1191
rect 3034 1188 3174 1191
rect 3210 1188 3214 1191
rect 3282 1188 3462 1191
rect 3482 1188 3486 1191
rect 3658 1188 3678 1191
rect 3730 1188 3734 1191
rect 3746 1188 3782 1191
rect 3794 1188 3806 1191
rect 3898 1188 3942 1191
rect 4066 1188 4110 1191
rect 4114 1188 4182 1191
rect 4186 1188 4374 1191
rect 4394 1188 4582 1191
rect 30 1182 33 1188
rect 74 1178 166 1181
rect 170 1178 286 1181
rect 290 1178 526 1181
rect 1442 1178 1606 1181
rect 1610 1178 1646 1181
rect 1650 1178 1670 1181
rect 1718 1181 1721 1188
rect 1674 1178 1721 1181
rect 1826 1178 1894 1181
rect 1998 1181 2001 1188
rect 1930 1178 2318 1181
rect 2338 1178 2350 1181
rect 2354 1178 2622 1181
rect 2626 1178 3774 1181
rect 3778 1178 3998 1181
rect 4026 1178 4150 1181
rect 4162 1178 4182 1181
rect 4210 1178 4222 1181
rect 4282 1178 4310 1181
rect 4354 1178 4446 1181
rect -26 1171 -22 1172
rect 54 1171 57 1178
rect -26 1168 57 1171
rect 330 1168 350 1171
rect 354 1168 406 1171
rect 718 1171 721 1178
rect 718 1168 742 1171
rect 762 1168 878 1171
rect 882 1168 918 1171
rect 1178 1168 1182 1171
rect 1250 1168 1262 1171
rect 1378 1168 1478 1171
rect 1610 1168 1702 1171
rect 1786 1168 1838 1171
rect 1874 1168 1902 1171
rect 1962 1168 2038 1171
rect 2326 1171 2329 1178
rect 2326 1168 2366 1171
rect 2490 1168 2678 1171
rect 2682 1168 2742 1171
rect 2786 1168 2814 1171
rect 2826 1168 2838 1171
rect 2858 1168 2862 1171
rect 2882 1168 2886 1171
rect 3018 1168 3254 1171
rect 3266 1168 3438 1171
rect 3442 1168 3470 1171
rect 3506 1168 3926 1171
rect 3970 1168 4070 1171
rect 4074 1168 4102 1171
rect 4106 1168 4254 1171
rect 4426 1168 4566 1171
rect 454 1162 457 1168
rect 50 1158 78 1161
rect 146 1158 302 1161
rect 306 1158 398 1161
rect 478 1161 481 1168
rect 654 1162 657 1168
rect 474 1158 481 1161
rect 498 1158 566 1161
rect 618 1158 638 1161
rect 706 1158 974 1161
rect 990 1161 993 1168
rect 1014 1161 1017 1168
rect 990 1158 1017 1161
rect 1034 1158 1062 1161
rect 1086 1161 1089 1168
rect 1086 1158 1094 1161
rect 1122 1158 1158 1161
rect 1234 1158 1262 1161
rect 1362 1158 1398 1161
rect 1410 1158 1438 1161
rect 1442 1158 1454 1161
rect 1498 1158 1542 1161
rect 1626 1158 1734 1161
rect 1802 1158 1934 1161
rect 1962 1158 2126 1161
rect 2170 1158 2246 1161
rect 2266 1158 2342 1161
rect 2426 1158 2454 1161
rect 2474 1158 2582 1161
rect 2586 1158 2622 1161
rect 2626 1158 2673 1161
rect 2754 1158 2926 1161
rect 2938 1158 2958 1161
rect 2998 1161 3001 1168
rect 4598 1162 4601 1168
rect 2998 1158 3030 1161
rect 3042 1158 3094 1161
rect 3114 1158 3118 1161
rect 3130 1158 3142 1161
rect 3186 1158 3190 1161
rect 3274 1158 3342 1161
rect 3354 1158 3358 1161
rect 3386 1158 3414 1161
rect 3418 1158 3438 1161
rect 3450 1158 3454 1161
rect 3490 1158 3526 1161
rect 3538 1158 3582 1161
rect 3594 1158 3686 1161
rect 3690 1158 3822 1161
rect 3834 1158 3905 1161
rect 3914 1158 3998 1161
rect 4010 1158 4014 1161
rect 4138 1158 4142 1161
rect 4210 1158 4270 1161
rect 4442 1158 4462 1161
rect 4490 1158 4518 1161
rect 4538 1158 4558 1161
rect 406 1152 409 1158
rect -26 1151 -22 1152
rect -26 1148 6 1151
rect 162 1148 209 1151
rect 442 1148 470 1151
rect 582 1151 585 1158
rect 562 1148 585 1151
rect 650 1148 670 1151
rect 698 1148 718 1151
rect 722 1148 758 1151
rect 762 1148 766 1151
rect 786 1148 790 1151
rect 794 1148 806 1151
rect 1058 1148 1062 1151
rect 1066 1148 1078 1151
rect 1082 1148 1134 1151
rect 1210 1148 1222 1151
rect 1290 1148 1302 1151
rect 1322 1148 1350 1151
rect 1410 1148 1433 1151
rect 1490 1148 1550 1151
rect 1734 1151 1737 1158
rect 2350 1152 2353 1158
rect 1734 1148 1742 1151
rect 1794 1148 1806 1151
rect 1810 1148 1814 1151
rect 1894 1148 1950 1151
rect 1970 1148 2046 1151
rect 2066 1148 2158 1151
rect 2170 1148 2270 1151
rect 2354 1148 2390 1151
rect 2394 1148 2398 1151
rect 2434 1148 2438 1151
rect 2482 1148 2486 1151
rect 2610 1148 2646 1151
rect 2670 1151 2673 1158
rect 3902 1152 3905 1158
rect 2670 1148 2758 1151
rect 2770 1148 2774 1151
rect 2802 1148 2918 1151
rect 2922 1148 3006 1151
rect 3042 1148 3046 1151
rect 3114 1148 3502 1151
rect 3522 1148 3646 1151
rect 3650 1148 3697 1151
rect 3738 1148 3742 1151
rect 3746 1148 3766 1151
rect 3850 1148 3886 1151
rect 3970 1148 4017 1151
rect 4042 1148 4166 1151
rect 4194 1148 4198 1151
rect 4290 1148 4310 1151
rect 4402 1148 4422 1151
rect 4434 1148 4438 1151
rect 206 1142 209 1148
rect 234 1138 398 1141
rect 450 1138 542 1141
rect 578 1138 606 1141
rect 902 1141 905 1148
rect 858 1138 905 1141
rect 1074 1138 1102 1141
rect 1106 1138 1142 1141
rect 1146 1138 1222 1141
rect 1246 1141 1249 1148
rect 1430 1142 1433 1148
rect 1686 1142 1689 1148
rect 1246 1138 1382 1141
rect 1530 1138 1662 1141
rect 1694 1141 1697 1148
rect 1694 1138 1766 1141
rect 1846 1141 1849 1148
rect 1878 1141 1881 1148
rect 1846 1138 1881 1141
rect 1894 1142 1897 1148
rect 1918 1138 1942 1141
rect 1946 1138 2086 1141
rect 2090 1138 2102 1141
rect 2122 1138 2214 1141
rect 2230 1138 2286 1141
rect 2402 1138 2406 1141
rect 2434 1138 2494 1141
rect 2514 1138 2558 1141
rect 2562 1138 2606 1141
rect 2626 1138 2630 1141
rect 2658 1138 2662 1141
rect 2698 1138 2878 1141
rect 2914 1138 2990 1141
rect 3018 1138 3094 1141
rect 3106 1138 3134 1141
rect 3138 1138 3150 1141
rect 3194 1138 3270 1141
rect 3282 1138 3286 1141
rect 3306 1138 3310 1141
rect 3330 1138 3406 1141
rect 3418 1138 3454 1141
rect 3474 1138 3510 1141
rect 3570 1138 3630 1141
rect 3634 1138 3686 1141
rect 3694 1141 3697 1148
rect 3790 1142 3793 1148
rect 4014 1142 4017 1148
rect 4262 1142 4265 1148
rect 3694 1138 3710 1141
rect 3714 1138 3758 1141
rect 3802 1138 3870 1141
rect 3874 1138 3910 1141
rect 4122 1138 4126 1141
rect 4154 1138 4222 1141
rect 4266 1138 4278 1141
rect 4314 1138 4334 1141
rect 4482 1138 4486 1141
rect 322 1128 326 1131
rect 530 1128 534 1131
rect 538 1128 830 1131
rect 906 1128 942 1131
rect 998 1128 1086 1131
rect 1090 1128 1118 1131
rect 1242 1128 1286 1131
rect 1298 1128 1406 1131
rect 1414 1131 1417 1138
rect 1918 1132 1921 1138
rect 1414 1128 1446 1131
rect 1458 1128 1646 1131
rect 1682 1128 1830 1131
rect 1950 1128 1958 1131
rect 1962 1128 1990 1131
rect 2002 1128 2022 1131
rect 2050 1128 2054 1131
rect 2118 1131 2121 1138
rect 2114 1128 2121 1131
rect 2230 1131 2233 1138
rect 2210 1128 2233 1131
rect 2242 1128 2246 1131
rect 2414 1131 2417 1138
rect 2314 1128 2417 1131
rect 2474 1128 2502 1131
rect 2570 1128 2574 1131
rect 2594 1128 2606 1131
rect 2610 1128 2646 1131
rect 2650 1128 2926 1131
rect 2930 1128 3118 1131
rect 3122 1128 3254 1131
rect 3258 1128 3294 1131
rect 3298 1128 3318 1131
rect 3334 1128 3342 1131
rect 3346 1128 3366 1131
rect 3454 1131 3457 1138
rect 3454 1128 3478 1131
rect 3482 1128 3502 1131
rect 3538 1128 3550 1131
rect 3562 1128 3574 1131
rect 3610 1128 3614 1131
rect 3634 1128 3678 1131
rect 3690 1128 3742 1131
rect 3770 1128 3782 1131
rect 3786 1128 3793 1131
rect 3834 1128 3870 1131
rect 3898 1128 3990 1131
rect 4074 1128 4110 1131
rect 4122 1128 4134 1131
rect 4154 1128 4158 1131
rect 4162 1128 4174 1131
rect 4234 1128 4238 1131
rect 4322 1128 4326 1131
rect 4482 1128 4558 1131
rect 26 1118 134 1121
rect 138 1118 350 1121
rect 402 1118 486 1121
rect 606 1118 622 1121
rect 998 1121 1001 1128
rect 946 1118 1001 1121
rect 1042 1118 1126 1121
rect 1234 1118 1358 1121
rect 1362 1118 1486 1121
rect 1638 1121 1641 1128
rect 1638 1118 1870 1121
rect 1922 1118 2073 1121
rect 2114 1118 2158 1121
rect 2234 1118 2398 1121
rect 2458 1118 2550 1121
rect 2554 1118 2638 1121
rect 2718 1118 2742 1121
rect 2906 1118 2934 1121
rect 2938 1118 2942 1121
rect 2950 1118 2974 1121
rect 2986 1118 2990 1121
rect 3002 1118 3014 1121
rect 3090 1118 3166 1121
rect 3210 1118 3278 1121
rect 3282 1118 3326 1121
rect 3530 1118 3582 1121
rect 3674 1118 3710 1121
rect 3750 1121 3753 1128
rect 3750 1118 3758 1121
rect 3786 1118 3966 1121
rect 3970 1118 4342 1121
rect 4346 1118 4590 1121
rect 306 1108 310 1111
rect 606 1111 609 1118
rect 418 1108 609 1111
rect 618 1108 670 1111
rect 1194 1108 1214 1111
rect 1242 1108 1342 1111
rect 1454 1108 1550 1111
rect 1618 1108 1678 1111
rect 1690 1108 1790 1111
rect 1818 1108 1870 1111
rect 1986 1108 2006 1111
rect 2070 1111 2073 1118
rect 2702 1112 2705 1118
rect 2718 1112 2721 1118
rect 2070 1108 2190 1111
rect 2418 1108 2438 1111
rect 2450 1108 2662 1111
rect 2950 1111 2953 1118
rect 2802 1108 2953 1111
rect 2962 1108 3038 1111
rect 3074 1108 3110 1111
rect 3146 1108 3238 1111
rect 3266 1108 3270 1111
rect 3306 1108 3382 1111
rect 3458 1108 3630 1111
rect 3666 1108 3774 1111
rect 4034 1108 4038 1111
rect 4218 1108 4382 1111
rect 4402 1108 4422 1111
rect 4426 1108 4502 1111
rect 678 1102 681 1108
rect 1000 1103 1002 1107
rect 1006 1103 1009 1107
rect 1014 1103 1016 1107
rect 298 1098 478 1101
rect 1122 1098 1158 1101
rect 1162 1098 1198 1101
rect 1202 1098 1302 1101
rect 1370 1098 1422 1101
rect 1454 1101 1457 1108
rect 2024 1103 2026 1107
rect 2030 1103 2033 1107
rect 2038 1103 2040 1107
rect 2358 1102 2361 1108
rect 3048 1103 3050 1107
rect 3054 1103 3057 1107
rect 3062 1103 3064 1107
rect 3846 1102 3849 1108
rect 3854 1102 3857 1108
rect 4080 1103 4082 1107
rect 4086 1103 4089 1107
rect 4094 1103 4096 1107
rect 4126 1102 4129 1108
rect 1426 1098 1457 1101
rect 1482 1098 1486 1101
rect 1546 1098 1614 1101
rect 1618 1098 1694 1101
rect 1782 1098 1945 1101
rect 1994 1098 1998 1101
rect 2306 1098 2326 1101
rect 2338 1098 2350 1101
rect 2370 1098 2470 1101
rect 2490 1098 2614 1101
rect 2626 1098 2782 1101
rect 3074 1098 3134 1101
rect 3142 1098 3174 1101
rect 3194 1098 3534 1101
rect 3538 1098 3542 1101
rect 3546 1098 3566 1101
rect 3698 1098 3710 1101
rect 3714 1098 3790 1101
rect 3922 1098 3942 1101
rect 3946 1098 4030 1101
rect 4258 1098 4302 1101
rect 4338 1098 4414 1101
rect 4434 1098 4494 1101
rect 1358 1092 1361 1098
rect 1782 1092 1785 1098
rect 122 1088 598 1091
rect 690 1088 702 1091
rect 706 1088 838 1091
rect 1050 1088 1126 1091
rect 1134 1088 1142 1091
rect 1146 1088 1238 1091
rect 1266 1088 1294 1091
rect 1362 1088 1430 1091
rect 1438 1088 1494 1091
rect 1514 1088 1654 1091
rect 1758 1088 1766 1091
rect 1770 1088 1782 1091
rect 1794 1088 1846 1091
rect 1942 1091 1945 1098
rect 2830 1092 2833 1098
rect 1942 1088 2134 1091
rect 2146 1088 2150 1091
rect 2406 1088 2670 1091
rect 2682 1088 2742 1091
rect 2850 1088 2886 1091
rect 2906 1088 2910 1091
rect 2930 1088 2942 1091
rect 2978 1088 3070 1091
rect 3142 1091 3145 1098
rect 3114 1088 3145 1091
rect 3162 1088 3630 1091
rect 3734 1088 3766 1091
rect 3786 1088 3854 1091
rect 3878 1088 3985 1091
rect 3994 1088 4150 1091
rect 4194 1088 4270 1091
rect 4330 1088 4350 1091
rect 4362 1088 4454 1091
rect 274 1078 454 1081
rect 458 1078 526 1081
rect 666 1078 702 1081
rect 706 1078 742 1081
rect 1026 1078 1062 1081
rect 1074 1078 1190 1081
rect 1194 1078 1382 1081
rect 1438 1081 1441 1088
rect 2406 1082 2409 1088
rect 3734 1082 3737 1088
rect 3878 1082 3881 1088
rect 3982 1082 3985 1088
rect 4486 1082 4489 1088
rect 1410 1078 1441 1081
rect 1450 1078 1558 1081
rect 1658 1078 1774 1081
rect 1850 1078 1886 1081
rect 1938 1078 1998 1081
rect 2058 1078 2158 1081
rect 2178 1078 2182 1081
rect 2218 1078 2270 1081
rect 2274 1078 2374 1081
rect 2498 1078 2502 1081
rect 2538 1078 2678 1081
rect 2714 1078 2774 1081
rect 2818 1078 2825 1081
rect 2834 1078 2934 1081
rect 2938 1078 3041 1081
rect 3178 1078 3262 1081
rect 3314 1078 3318 1081
rect 3362 1078 3398 1081
rect 3426 1078 3430 1081
rect 3434 1078 3454 1081
rect 3514 1078 3518 1081
rect 3542 1078 3590 1081
rect 3602 1078 3622 1081
rect 3770 1078 3798 1081
rect 3810 1078 3814 1081
rect 3906 1078 3926 1081
rect 4058 1078 4078 1081
rect 4114 1078 4134 1081
rect 4170 1078 4190 1081
rect 4218 1078 4278 1081
rect 4338 1078 4342 1081
rect 4418 1078 4454 1081
rect -26 1071 -22 1072
rect 30 1071 33 1078
rect 918 1072 921 1078
rect 2206 1072 2209 1078
rect -26 1068 33 1071
rect 50 1068 150 1071
rect 154 1068 270 1071
rect 306 1068 310 1071
rect 314 1068 414 1071
rect 418 1068 438 1071
rect 586 1068 681 1071
rect 922 1068 950 1071
rect 954 1068 1174 1071
rect 1218 1068 1230 1071
rect 1314 1068 1350 1071
rect 1354 1068 1446 1071
rect 1458 1068 1470 1071
rect 1642 1068 1718 1071
rect 1778 1068 1854 1071
rect 1906 1068 1990 1071
rect 2018 1068 2046 1071
rect 2050 1068 2070 1071
rect 2098 1068 2102 1071
rect 2162 1068 2182 1071
rect 2214 1071 2217 1078
rect 2814 1072 2817 1078
rect 2822 1072 2825 1078
rect 2214 1068 2246 1071
rect 2306 1068 2350 1071
rect 2374 1068 2390 1071
rect 2410 1068 2446 1071
rect 2514 1068 2590 1071
rect 2658 1068 2662 1071
rect 2690 1068 2718 1071
rect 2754 1068 2798 1071
rect 2830 1068 2894 1071
rect 2898 1068 2958 1071
rect 3002 1068 3006 1071
rect 3026 1068 3030 1071
rect 3038 1071 3041 1078
rect 3350 1072 3353 1078
rect 3038 1068 3198 1071
rect 3266 1068 3294 1071
rect 3330 1068 3334 1071
rect 3394 1068 3430 1071
rect 3474 1068 3486 1071
rect 3542 1071 3545 1078
rect 3638 1072 3641 1078
rect 4198 1072 4201 1078
rect 4294 1072 4297 1078
rect 4478 1072 4481 1078
rect 3538 1068 3545 1071
rect 3570 1068 3574 1071
rect 3610 1068 3614 1071
rect 3674 1068 3678 1071
rect 3706 1068 3734 1071
rect 3738 1068 3782 1071
rect 3794 1068 3838 1071
rect 3842 1068 3878 1071
rect 3882 1068 3918 1071
rect 3962 1068 3974 1071
rect 4042 1068 4094 1071
rect 4098 1068 4158 1071
rect 4242 1068 4254 1071
rect 4334 1068 4366 1071
rect 4402 1068 4422 1071
rect 4458 1068 4462 1071
rect 4482 1068 4534 1071
rect 678 1062 681 1068
rect 22 1058 30 1061
rect 34 1058 54 1061
rect 162 1058 230 1061
rect 234 1058 249 1061
rect 274 1058 310 1061
rect 354 1058 366 1061
rect 434 1058 438 1061
rect 550 1058 598 1061
rect 682 1059 750 1061
rect 1990 1062 1993 1068
rect 682 1058 753 1059
rect 938 1058 982 1061
rect 1178 1058 1190 1061
rect 1298 1058 1302 1061
rect 1322 1058 1382 1061
rect 1426 1058 1438 1061
rect 1482 1058 1486 1061
rect 1506 1058 1582 1061
rect 1586 1058 1630 1061
rect 1730 1058 1846 1061
rect 1930 1058 1950 1061
rect 1962 1058 1966 1061
rect 2090 1058 2094 1061
rect 2114 1058 2126 1061
rect 2130 1058 2206 1061
rect 2226 1058 2254 1061
rect 2330 1058 2334 1061
rect 2374 1061 2377 1068
rect 2614 1062 2617 1068
rect 2726 1062 2729 1068
rect 2346 1058 2377 1061
rect 2382 1058 2438 1061
rect 2442 1058 2454 1061
rect 2490 1058 2582 1061
rect 2658 1058 2694 1061
rect 2786 1058 2798 1061
rect 2802 1058 2806 1061
rect 2830 1061 2833 1068
rect 3014 1062 3017 1068
rect 3238 1062 3241 1068
rect 3502 1062 3505 1068
rect 3542 1062 3545 1068
rect 2818 1058 2833 1061
rect 2882 1058 2886 1061
rect 2918 1058 2926 1061
rect 2930 1058 3006 1061
rect 3034 1058 3038 1061
rect 3058 1058 3118 1061
rect 3122 1058 3126 1061
rect 3186 1058 3190 1061
rect 3210 1058 3214 1061
rect 3314 1058 3382 1061
rect 3410 1058 3465 1061
rect 3586 1058 3590 1061
rect 3658 1058 3694 1061
rect 3722 1058 3774 1061
rect 3778 1058 3862 1061
rect 3962 1058 3966 1061
rect 4014 1061 4017 1068
rect 3994 1058 4017 1061
rect 4050 1058 4062 1061
rect 4182 1061 4185 1068
rect 4334 1062 4337 1068
rect 4182 1058 4198 1061
rect 4338 1058 4438 1061
rect 4458 1058 4486 1061
rect 4510 1058 4534 1061
rect 246 1052 249 1058
rect 550 1052 553 1058
rect -26 1051 -22 1052
rect -26 1048 6 1051
rect 354 1048 438 1051
rect 674 1048 694 1051
rect 926 1048 958 1051
rect 1002 1048 1038 1051
rect 1274 1048 1326 1051
rect 1330 1048 1494 1051
rect 1602 1048 1622 1051
rect 1714 1048 1758 1051
rect 1762 1048 1774 1051
rect 1834 1048 1854 1051
rect 1858 1048 1998 1051
rect 2066 1048 2086 1051
rect 2102 1051 2105 1058
rect 2382 1052 2385 1058
rect 2102 1048 2150 1051
rect 2154 1048 2182 1051
rect 2210 1048 2222 1051
rect 2250 1048 2270 1051
rect 2322 1048 2382 1051
rect 2426 1048 2518 1051
rect 2526 1048 2558 1051
rect 2590 1051 2593 1058
rect 2694 1052 2697 1058
rect 2590 1048 2654 1051
rect 2702 1051 2705 1058
rect 2702 1048 2766 1051
rect 2874 1048 3094 1051
rect 3122 1048 3150 1051
rect 3270 1051 3273 1058
rect 3162 1048 3273 1051
rect 3338 1048 3358 1051
rect 3386 1048 3390 1051
rect 3450 1048 3454 1051
rect 3462 1051 3465 1058
rect 4510 1052 4513 1058
rect 3462 1048 3502 1051
rect 3666 1048 3670 1051
rect 3778 1048 3798 1051
rect 3826 1048 3830 1051
rect 3842 1048 3846 1051
rect 3850 1048 3918 1051
rect 3946 1048 3958 1051
rect 4010 1048 4046 1051
rect 4122 1048 4310 1051
rect 4338 1048 4390 1051
rect 4402 1048 4406 1051
rect 4442 1048 4446 1051
rect 926 1042 929 1048
rect 346 1038 614 1041
rect 970 1038 974 1041
rect 1306 1038 1342 1041
rect 1346 1038 1393 1041
rect 1466 1038 1646 1041
rect 1878 1038 2094 1041
rect 2106 1038 2166 1041
rect 2526 1041 2529 1048
rect 2186 1038 2529 1041
rect 2554 1038 2614 1041
rect 2702 1041 2705 1048
rect 2618 1038 2705 1041
rect 2770 1038 2790 1041
rect 2946 1038 2982 1041
rect 2994 1038 2998 1041
rect 3098 1038 3190 1041
rect 3218 1038 3222 1041
rect 3242 1038 3430 1041
rect 3490 1038 3494 1041
rect 3518 1041 3521 1048
rect 3702 1042 3705 1048
rect 3742 1042 3745 1048
rect 3518 1038 3694 1041
rect 3758 1041 3761 1048
rect 3758 1038 3918 1041
rect 3930 1038 4094 1041
rect 4106 1038 4438 1041
rect 4442 1038 4526 1041
rect 4546 1038 4558 1041
rect 1390 1032 1393 1038
rect 1878 1032 1881 1038
rect 358 1028 382 1031
rect 394 1028 694 1031
rect 914 1028 1030 1031
rect 1058 1028 1062 1031
rect 1146 1028 1302 1031
rect 1594 1028 1686 1031
rect 1690 1028 1694 1031
rect 1890 1028 2086 1031
rect 2090 1028 2198 1031
rect 2210 1028 2262 1031
rect 2282 1028 2478 1031
rect 2514 1028 2566 1031
rect 2766 1031 2769 1038
rect 2570 1028 2769 1031
rect 2906 1028 2950 1031
rect 2978 1028 3134 1031
rect 3138 1028 3993 1031
rect 4002 1028 4006 1031
rect 4018 1028 4198 1031
rect 4266 1028 4286 1031
rect 4294 1028 4302 1031
rect 4306 1028 4382 1031
rect 4442 1028 4550 1031
rect 4554 1028 4598 1031
rect 358 1022 361 1028
rect 394 1018 1086 1021
rect 1218 1018 1278 1021
rect 1414 1021 1417 1028
rect 1282 1018 1417 1021
rect 1770 1018 2646 1021
rect 2674 1018 2718 1021
rect 2778 1018 2846 1021
rect 2882 1018 2942 1021
rect 2954 1018 3270 1021
rect 3282 1018 3326 1021
rect 3354 1018 3454 1021
rect 3482 1018 3726 1021
rect 3730 1018 3750 1021
rect 3770 1018 3950 1021
rect 3990 1021 3993 1028
rect 3990 1018 4022 1021
rect 4026 1018 4182 1021
rect 4186 1018 4326 1021
rect 4330 1018 4350 1021
rect 4442 1018 4566 1021
rect 4382 1012 4385 1018
rect 218 1008 374 1011
rect 1562 1008 1830 1011
rect 2002 1008 2038 1011
rect 2178 1008 2286 1011
rect 2290 1008 2310 1011
rect 2322 1008 2454 1011
rect 2642 1008 2750 1011
rect 2754 1008 3070 1011
rect 3130 1008 3142 1011
rect 3170 1008 3206 1011
rect 3210 1008 3278 1011
rect 3282 1008 3470 1011
rect 3474 1008 3526 1011
rect 3746 1008 3838 1011
rect 3866 1008 4006 1011
rect 4138 1008 4190 1011
rect 4210 1008 4374 1011
rect 4394 1008 4454 1011
rect 496 1003 498 1007
rect 502 1003 505 1007
rect 510 1003 512 1007
rect 1520 1003 1522 1007
rect 1526 1003 1529 1007
rect 1534 1003 1536 1007
rect 2544 1003 2546 1007
rect 2550 1003 2553 1007
rect 2558 1003 2560 1007
rect 3568 1003 3570 1007
rect 3574 1003 3577 1007
rect 3582 1003 3584 1007
rect 210 998 222 1001
rect 226 998 278 1001
rect 282 998 326 1001
rect 978 998 1134 1001
rect 1170 998 1198 1001
rect 1714 998 1838 1001
rect 1842 998 1862 1001
rect 1890 998 1894 1001
rect 2010 998 2054 1001
rect 2170 998 2230 1001
rect 2242 998 2350 1001
rect 2634 998 2638 1001
rect 2658 998 2710 1001
rect 2746 998 2774 1001
rect 2938 998 2942 1001
rect 2978 998 2998 1001
rect 3002 998 3198 1001
rect 3226 998 3230 1001
rect 3250 998 3382 1001
rect 3390 998 3494 1001
rect 3530 998 3558 1001
rect 3666 998 3734 1001
rect 3754 998 3806 1001
rect 3986 998 4070 1001
rect 4170 998 4246 1001
rect 4258 998 4598 1001
rect 98 988 390 991
rect 422 988 574 991
rect 578 988 622 991
rect 870 988 1510 991
rect 1514 988 1854 991
rect 1858 988 1870 991
rect 1874 988 1902 991
rect 2178 988 2214 991
rect 2218 988 2398 991
rect 2402 988 2886 991
rect 2890 988 3062 991
rect 3246 991 3249 998
rect 3390 992 3393 998
rect 3066 988 3249 991
rect 3262 988 3334 991
rect 3342 988 3374 991
rect 4254 991 4257 998
rect 3490 988 4257 991
rect 4386 988 4390 991
rect 4410 988 4494 991
rect 422 982 425 988
rect 870 982 873 988
rect 2054 982 2057 988
rect 3262 982 3265 988
rect 3342 982 3345 988
rect 246 978 406 981
rect 1130 978 1366 981
rect 1378 978 1446 981
rect 1450 978 1486 981
rect 1674 978 1742 981
rect 1754 978 1782 981
rect 1814 978 2030 981
rect 2282 978 2478 981
rect 2506 978 2678 981
rect 2714 978 2782 981
rect 2814 978 2862 981
rect 2882 978 3254 981
rect 3330 978 3334 981
rect 3442 978 3550 981
rect 3554 978 4230 981
rect 4234 978 4470 981
rect 246 972 249 978
rect 454 971 457 978
rect 454 968 478 971
rect 654 971 657 978
rect 1814 972 1817 978
rect 498 968 657 971
rect 1050 968 1566 971
rect 1570 968 1702 971
rect 1706 968 1758 971
rect 1882 968 1886 971
rect 1938 968 1942 971
rect 2094 968 2142 971
rect 2250 968 2294 971
rect 2298 968 2318 971
rect 2322 968 2358 971
rect 2374 968 2505 971
rect 2514 968 2582 971
rect 2814 971 2817 978
rect 2586 968 2817 971
rect 2826 968 2838 971
rect 2862 971 2865 978
rect 2862 968 2910 971
rect 2978 968 3017 971
rect 3106 968 3150 971
rect 3154 968 3161 971
rect 3178 968 3182 971
rect 3202 968 3262 971
rect 3322 968 3390 971
rect 3398 971 3401 978
rect 3394 968 3401 971
rect 3434 968 3558 971
rect 3578 968 3646 971
rect 3682 968 3686 971
rect 3706 968 3726 971
rect 3738 968 3782 971
rect 3806 968 3865 971
rect 310 962 313 968
rect 146 958 278 961
rect 402 958 510 961
rect 514 958 558 961
rect 906 958 918 961
rect 954 958 974 961
rect 978 958 1014 961
rect 1018 958 1022 961
rect 1074 958 1078 961
rect 1146 958 1150 961
rect 1186 958 1198 961
rect 1218 958 1270 961
rect 1370 958 1438 961
rect 1442 958 1470 961
rect 1482 958 1542 961
rect 1674 958 1726 961
rect 1730 958 1798 961
rect 1846 961 1849 968
rect 2094 962 2097 968
rect 2374 962 2377 968
rect 1846 958 1878 961
rect 1890 958 1894 961
rect 1986 958 2014 961
rect 2210 958 2278 961
rect 2290 958 2366 961
rect 2426 958 2454 961
rect 2502 961 2505 968
rect 2502 958 2518 961
rect 2626 958 2630 961
rect 2674 958 2894 961
rect 2966 961 2969 968
rect 3014 962 3017 968
rect 3798 962 3801 968
rect 3806 962 3809 968
rect 3862 962 3865 968
rect 3938 968 4110 971
rect 4418 968 4446 971
rect 4458 968 4526 971
rect 4530 968 4537 971
rect 2966 958 2990 961
rect 3058 958 3078 961
rect 3090 958 3094 961
rect 3130 958 3350 961
rect 3354 958 3358 961
rect 3458 958 3542 961
rect 3550 958 3622 961
rect 3626 958 3633 961
rect 3642 958 3670 961
rect 3690 958 3766 961
rect 3874 958 3878 961
rect 3910 961 3913 968
rect 3890 958 3913 961
rect 4074 958 4134 961
rect 4286 961 4289 968
rect 4274 958 4289 961
rect 4362 958 4366 961
rect 4402 958 4417 961
rect 4434 958 4465 961
rect 4474 958 4486 961
rect 4490 958 4510 961
rect -26 951 -22 952
rect -26 948 6 951
rect 202 948 214 951
rect 266 948 286 951
rect 314 948 358 951
rect 370 948 390 951
rect 394 948 446 951
rect 474 948 630 951
rect 806 951 809 958
rect 706 948 809 951
rect 930 948 1054 951
rect 1166 951 1169 958
rect 2198 952 2201 958
rect 2406 952 2409 958
rect 2606 952 2609 958
rect 3406 952 3409 958
rect 1166 948 1190 951
rect 1226 948 1262 951
rect 1434 948 1478 951
rect 1490 948 1494 951
rect 1554 948 1590 951
rect 1618 948 1686 951
rect 1698 948 1766 951
rect 1826 948 1846 951
rect 1850 948 1918 951
rect 1922 948 2102 951
rect 2162 948 2174 951
rect 2202 948 2230 951
rect 2250 948 2374 951
rect 2514 948 2518 951
rect 2546 948 2550 951
rect 2578 948 2598 951
rect 2610 948 2790 951
rect 2802 948 2806 951
rect 2826 948 2870 951
rect 2890 948 2894 951
rect 2914 948 2974 951
rect 3002 948 3006 951
rect 3042 948 3206 951
rect 3226 948 3230 951
rect 3250 948 3262 951
rect 3266 948 3358 951
rect 3426 948 3526 951
rect 3550 951 3553 958
rect 3830 952 3833 958
rect 4318 952 4321 958
rect 4414 952 4417 958
rect 3538 948 3553 951
rect 3570 948 3622 951
rect 3626 948 3646 951
rect 3674 948 3678 951
rect 3730 948 3734 951
rect 3762 948 3766 951
rect 3850 948 3886 951
rect 3906 948 3950 951
rect 3978 948 3982 951
rect 3994 948 3998 951
rect 4090 948 4094 951
rect 4098 948 4118 951
rect 4138 948 4150 951
rect 4170 948 4174 951
rect 4194 948 4198 951
rect 4234 948 4238 951
rect 4258 948 4294 951
rect 4330 948 4350 951
rect 4462 951 4465 958
rect 4550 952 4553 958
rect 4462 948 4481 951
rect 1078 942 1081 948
rect 214 938 222 941
rect 226 938 289 941
rect 322 938 326 941
rect 330 938 406 941
rect 498 938 550 941
rect 618 938 742 941
rect 962 938 982 941
rect 986 938 990 941
rect 1158 941 1161 948
rect 1158 938 1222 941
rect 1234 938 1294 941
rect 1354 938 1606 941
rect 1666 938 1710 941
rect 1722 938 1766 941
rect 1834 938 1982 941
rect 2034 938 2126 941
rect 2154 938 2158 941
rect 2178 938 2182 941
rect 2194 938 2233 941
rect 2274 938 2278 941
rect 2338 938 2390 941
rect 2394 938 2398 941
rect 2414 941 2417 948
rect 2422 941 2425 948
rect 3782 942 3785 948
rect 4454 942 4457 948
rect 4478 942 4481 948
rect 4558 942 4561 948
rect 2414 938 2425 941
rect 2434 938 2678 941
rect 2682 938 2782 941
rect 2786 938 2806 941
rect 2866 938 2878 941
rect 2906 938 2910 941
rect 2922 938 2926 941
rect 2930 938 2950 941
rect 2962 938 2966 941
rect 2978 938 2998 941
rect 3050 938 3054 941
rect 3098 938 3102 941
rect 3106 938 3113 941
rect 3130 938 3158 941
rect 3170 938 3174 941
rect 3234 938 3238 941
rect 3322 938 3326 941
rect 3346 938 3350 941
rect 3378 938 3486 941
rect 3506 938 3518 941
rect 3546 938 3550 941
rect 3562 938 3598 941
rect 3602 938 3630 941
rect 3634 938 3686 941
rect 3698 938 3718 941
rect 3722 938 3750 941
rect 3802 938 3910 941
rect 3914 938 4014 941
rect 4034 938 4054 941
rect 4098 938 4102 941
rect 4114 938 4246 941
rect 4290 938 4310 941
rect 286 932 289 938
rect 1782 932 1785 938
rect 1982 932 1985 938
rect 2230 932 2233 938
rect 26 928 126 931
rect 130 928 182 931
rect 186 928 270 931
rect 370 928 382 931
rect 386 928 446 931
rect 450 928 518 931
rect 882 928 1158 931
rect 1170 928 1174 931
rect 1258 928 1374 931
rect 1418 928 1566 931
rect 1674 928 1742 931
rect 1818 928 1822 931
rect 1858 928 1886 931
rect 1930 928 1942 931
rect 2066 928 2070 931
rect 2082 928 2086 931
rect 2114 928 2158 931
rect 2406 931 2409 938
rect 2854 932 2857 938
rect 3262 932 3265 938
rect 2306 928 2337 931
rect 2406 928 2441 931
rect 2450 928 2454 931
rect 2486 928 2494 931
rect 2498 928 2518 931
rect 2586 928 2590 931
rect 2650 928 2670 931
rect 2694 928 2702 931
rect 2722 928 2806 931
rect 2862 928 2878 931
rect 2898 928 3094 931
rect 3098 928 3102 931
rect 3210 928 3222 931
rect 3282 928 3385 931
rect 3394 928 3398 931
rect 3402 928 3414 931
rect 3426 928 3430 931
rect 3442 928 3462 931
rect 3474 928 3478 931
rect 3498 928 3582 931
rect 3634 928 3654 931
rect 3674 928 3697 931
rect 3714 928 3774 931
rect 3850 928 3854 931
rect 3890 928 3894 931
rect 4026 928 4030 931
rect 4058 928 4118 931
rect 4306 928 4406 931
rect 4418 928 4502 931
rect 4550 931 4553 938
rect 4546 928 4553 931
rect 882 918 1281 921
rect 1290 918 1294 921
rect 1298 918 1398 921
rect 1466 918 1478 921
rect 1498 918 1678 921
rect 1694 918 1702 921
rect 1706 918 1726 921
rect 1738 918 1870 921
rect 1910 921 1913 928
rect 1910 918 1958 921
rect 1966 921 1969 928
rect 1966 918 1982 921
rect 1986 918 2110 921
rect 2138 918 2222 921
rect 2258 918 2326 921
rect 2334 921 2337 928
rect 2438 922 2441 928
rect 2862 922 2865 928
rect 2334 918 2406 921
rect 2450 918 2462 921
rect 2490 918 2502 921
rect 2538 918 2630 921
rect 2698 918 2742 921
rect 2778 918 2830 921
rect 2978 918 2990 921
rect 3010 918 3073 921
rect 3090 918 3094 921
rect 3238 921 3241 928
rect 3114 918 3241 921
rect 3338 918 3374 921
rect 3382 921 3385 928
rect 3614 922 3617 928
rect 3694 922 3697 928
rect 3382 918 3422 921
rect 3626 918 3630 921
rect 3746 918 3750 921
rect 3814 921 3817 928
rect 3770 918 3817 921
rect 3882 918 4030 921
rect 4050 918 4206 921
rect 4234 918 4310 921
rect 4314 918 4526 921
rect 4538 918 4574 921
rect 442 908 462 911
rect 602 908 798 911
rect 1178 908 1190 911
rect 1278 911 1281 918
rect 2766 912 2769 918
rect 1278 908 1470 911
rect 1474 908 1510 911
rect 1522 908 1590 911
rect 1634 908 1638 911
rect 1690 908 1838 911
rect 1946 908 1966 911
rect 2122 908 2225 911
rect 2234 908 2294 911
rect 2298 908 2470 911
rect 2474 908 2694 911
rect 2842 908 3030 911
rect 3070 911 3073 918
rect 4038 912 4041 918
rect 3070 908 3694 911
rect 3698 908 3966 911
rect 4186 908 4334 911
rect 4394 908 4478 911
rect 1000 903 1002 907
rect 1006 903 1009 907
rect 1014 903 1016 907
rect 2024 903 2026 907
rect 2030 903 2033 907
rect 2038 903 2040 907
rect 274 898 446 901
rect 450 898 622 901
rect 858 898 950 901
rect 1058 898 1118 901
rect 1154 898 1214 901
rect 1282 898 1398 901
rect 1402 898 1566 901
rect 1578 898 1630 901
rect 1874 898 1958 901
rect 2078 898 2206 901
rect 2222 901 2225 908
rect 3048 903 3050 907
rect 3054 903 3057 907
rect 3062 903 3064 907
rect 4080 903 4082 907
rect 4086 903 4089 907
rect 4094 903 4096 907
rect 2222 898 2278 901
rect 2354 898 2406 901
rect 2410 898 2601 901
rect 1638 892 1641 898
rect 678 888 966 891
rect 986 888 1142 891
rect 1162 888 1185 891
rect 1194 888 1254 891
rect 1274 888 1334 891
rect 1386 888 1462 891
rect 1482 888 1598 891
rect 1690 888 2001 891
rect 2078 891 2081 898
rect 2598 892 2601 898
rect 3226 898 3270 901
rect 3298 898 3310 901
rect 3346 898 3478 901
rect 3482 898 3638 901
rect 3650 898 3782 901
rect 3794 898 3806 901
rect 3850 898 4046 901
rect 4242 898 4262 901
rect 4274 898 4374 901
rect 4418 898 4486 901
rect 4522 898 4526 901
rect 2010 888 2081 891
rect 2122 888 2174 891
rect 2178 888 2302 891
rect 2378 888 2542 891
rect 2662 891 2665 898
rect 2602 888 2665 891
rect 2698 888 2710 891
rect 2754 888 2758 891
rect 2850 888 3046 891
rect 3050 888 3070 891
rect 3138 888 3198 891
rect 3218 888 3238 891
rect 3258 888 3270 891
rect 3290 888 3446 891
rect 3522 888 3534 891
rect 3610 888 3646 891
rect 3650 888 3662 891
rect 3714 888 3750 891
rect 3754 888 3774 891
rect 4002 888 4177 891
rect 678 882 681 888
rect 1182 882 1185 888
rect 186 878 222 881
rect 226 878 246 881
rect 434 878 646 881
rect 1090 878 1134 881
rect 1138 878 1166 881
rect 1290 878 1318 881
rect 1470 881 1473 888
rect 1998 882 2001 888
rect 1434 878 1473 881
rect 1594 878 1614 881
rect 1682 878 1686 881
rect 1762 878 1814 881
rect 1866 878 1926 881
rect 2050 878 2110 881
rect 2130 878 2134 881
rect 2226 878 2230 881
rect 2266 878 2294 881
rect 2298 878 2550 881
rect 2554 878 3302 881
rect 3306 878 3329 881
rect 3354 878 3358 881
rect 3362 878 3374 881
rect 3386 878 3390 881
rect 3462 881 3465 888
rect 3542 882 3545 888
rect 4174 882 4177 888
rect 4282 888 4553 891
rect 3394 878 3465 881
rect 3530 878 3534 881
rect 3570 878 3662 881
rect 3778 878 3822 881
rect 3826 878 3854 881
rect 3866 878 3926 881
rect 3938 878 3942 881
rect 3954 878 3982 881
rect 4026 878 4126 881
rect 4194 878 4198 881
rect 4210 878 4214 881
rect 4246 881 4249 888
rect 4550 882 4553 888
rect 4246 878 4281 881
rect -26 871 -22 872
rect 6 871 9 878
rect 934 872 937 878
rect -26 868 9 871
rect 134 868 153 871
rect 210 868 438 871
rect 674 868 694 871
rect 698 868 726 871
rect 730 868 742 871
rect 1034 868 1113 871
rect 1130 868 1142 871
rect 1194 868 1198 871
rect 1210 868 1214 871
rect 1286 871 1289 878
rect 1250 868 1289 871
rect 1298 868 1326 871
rect 1350 871 1353 878
rect 3326 872 3329 878
rect 3726 872 3729 878
rect 4278 872 4281 878
rect 4482 878 4486 881
rect 4570 878 4582 881
rect 1350 868 1374 871
rect 1378 868 1438 871
rect 1474 868 1478 871
rect 1618 868 1622 871
rect 1626 868 1638 871
rect 1698 868 1702 871
rect 1730 868 1758 871
rect 1762 868 1854 871
rect 2002 868 2022 871
rect 2026 870 2057 871
rect 2026 868 2054 870
rect 134 862 137 868
rect 150 862 153 868
rect 154 858 286 861
rect 378 858 486 861
rect 506 859 550 861
rect 502 858 550 859
rect 562 858 710 861
rect 714 859 822 861
rect 1110 862 1113 868
rect 1886 862 1889 868
rect 2154 868 2198 871
rect 2202 868 2254 871
rect 2274 868 2302 871
rect 2314 868 2318 871
rect 2346 868 2358 871
rect 2378 868 2382 871
rect 2394 868 2454 871
rect 2474 868 2478 871
rect 2506 868 2510 871
rect 2514 868 2574 871
rect 2642 868 2686 871
rect 2730 868 2766 871
rect 2770 868 2798 871
rect 2802 868 2886 871
rect 2890 868 2950 871
rect 2954 868 2958 871
rect 2970 868 2974 871
rect 2986 868 3014 871
rect 3026 868 3030 871
rect 3042 868 3046 871
rect 3138 868 3142 871
rect 3170 868 3174 871
rect 3210 868 3214 871
rect 3226 868 3254 871
rect 3298 868 3302 871
rect 3330 868 3350 871
rect 3354 868 3454 871
rect 3458 868 3558 871
rect 3562 868 3638 871
rect 3682 868 3694 871
rect 3738 868 3758 871
rect 3762 868 3790 871
rect 3810 868 3830 871
rect 3874 868 4110 871
rect 4178 868 4222 871
rect 4226 868 4238 871
rect 4326 871 4329 878
rect 4326 868 4366 871
rect 4434 868 4438 871
rect 714 858 825 859
rect 954 858 974 861
rect 1114 858 1166 861
rect 1234 858 1278 861
rect 1282 858 1326 861
rect 1466 858 1558 861
rect 1578 858 1630 861
rect 1738 858 1742 861
rect 1782 858 1790 861
rect 1938 858 1942 861
rect 2162 858 2166 861
rect 2194 858 2230 861
rect 2242 858 2422 861
rect 2426 858 2534 861
rect 2610 858 2638 861
rect 2722 858 2726 861
rect 2738 858 2742 861
rect 2770 858 2774 861
rect 2834 858 2846 861
rect 2858 858 2862 861
rect 2882 858 3102 861
rect 3110 861 3113 868
rect 4294 862 4297 868
rect 4318 862 4321 868
rect 3110 858 3126 861
rect 3130 858 3150 861
rect 3154 858 3166 861
rect 3170 858 3214 861
rect 3218 858 3270 861
rect 3314 858 3566 861
rect 3586 858 3590 861
rect 3650 858 3782 861
rect 3802 858 3822 861
rect 3826 858 3894 861
rect 3898 858 3942 861
rect 3946 858 3966 861
rect 3994 858 4062 861
rect 4066 858 4070 861
rect 4098 858 4198 861
rect 4202 858 4230 861
rect 4266 858 4270 861
rect 4282 858 4286 861
rect 4418 858 4422 861
rect 4474 858 4502 861
rect 4514 858 4518 861
rect 1782 852 1785 858
rect 2110 852 2113 858
rect 2126 852 2129 858
rect -26 851 -22 852
rect -26 848 30 851
rect 362 848 574 851
rect 666 848 702 851
rect 706 848 734 851
rect 978 848 1182 851
rect 1186 848 1190 851
rect 1226 848 1270 851
rect 1274 848 1278 851
rect 1322 848 1334 851
rect 1354 848 1398 851
rect 1418 848 1622 851
rect 1698 848 1729 851
rect 1738 848 1750 851
rect 1794 848 1814 851
rect 1954 848 2014 851
rect 2026 848 2046 851
rect 2186 848 2214 851
rect 2242 848 2358 851
rect 2370 848 2454 851
rect 2458 848 2494 851
rect 2498 848 2622 851
rect 2698 848 2742 851
rect 2750 848 2838 851
rect 2858 848 2862 851
rect 2866 848 2926 851
rect 2930 848 2982 851
rect 3066 848 3070 851
rect 3106 848 3110 851
rect 3130 848 3158 851
rect 3162 848 3286 851
rect 3302 848 3350 851
rect 3382 848 3390 851
rect 3402 848 3414 851
rect 3418 848 3502 851
rect 3586 848 3606 851
rect 3650 848 3654 851
rect 3662 848 3670 851
rect 3674 848 3686 851
rect 3786 848 3838 851
rect 3850 848 3889 851
rect 3914 848 3918 851
rect 3962 848 3966 851
rect 3986 848 4062 851
rect 4150 848 4158 851
rect 4194 848 4222 851
rect 4234 848 4249 851
rect 4290 848 4302 851
rect 4338 848 4382 851
rect 4458 848 4510 851
rect 1726 842 1729 848
rect 2230 842 2233 848
rect 378 838 558 841
rect 570 838 694 841
rect 1042 838 1214 841
rect 1426 838 1462 841
rect 1466 838 1534 841
rect 1594 838 1718 841
rect 1802 838 1814 841
rect 1818 838 1886 841
rect 1890 838 1910 841
rect 1914 838 2006 841
rect 2074 838 2102 841
rect 2146 838 2198 841
rect 2290 838 2310 841
rect 2338 838 2342 841
rect 2378 838 2414 841
rect 2450 838 2462 841
rect 2470 838 2478 841
rect 2530 838 2606 841
rect 2618 838 2662 841
rect 2666 838 2702 841
rect 2750 841 2753 848
rect 2730 838 2753 841
rect 2818 838 3150 841
rect 3162 838 3182 841
rect 3202 838 3206 841
rect 3222 838 3230 841
rect 3302 841 3305 848
rect 3886 842 3889 848
rect 3942 842 3945 848
rect 4246 842 4249 848
rect 4590 842 4593 848
rect 3234 838 3305 841
rect 3314 838 3414 841
rect 3426 838 3702 841
rect 3706 838 3766 841
rect 3818 838 3822 841
rect 3834 838 3870 841
rect 3958 838 3966 841
rect 3970 838 4006 841
rect 4034 838 4038 841
rect 4146 838 4198 841
rect 4298 838 4422 841
rect 4458 838 4518 841
rect 222 832 225 838
rect 338 828 726 831
rect 1906 828 1982 831
rect 1986 828 1990 831
rect 2066 828 2134 831
rect 2278 831 2281 838
rect 2278 828 2510 831
rect 2522 828 2822 831
rect 2962 828 3014 831
rect 3310 831 3313 838
rect 4214 832 4217 838
rect 3066 828 3313 831
rect 3410 828 3430 831
rect 3438 828 3454 831
rect 3546 828 3550 831
rect 3658 828 3782 831
rect 3810 828 3862 831
rect 3874 828 3990 831
rect 3994 828 4014 831
rect 4242 828 4326 831
rect 4370 828 4534 831
rect 122 818 774 821
rect 778 818 1102 821
rect 1330 818 1342 821
rect 1346 818 1510 821
rect 2074 818 2814 821
rect 2822 821 2825 828
rect 3438 822 3441 828
rect 2822 818 2958 821
rect 3026 818 3422 821
rect 3498 818 3510 821
rect 3554 818 3694 821
rect 3722 818 4182 821
rect 4210 818 4254 821
rect 4354 818 4430 821
rect 4442 818 4574 821
rect 650 808 758 811
rect 874 808 910 811
rect 1978 808 2174 811
rect 2250 808 2510 811
rect 2698 808 2710 811
rect 2730 808 2934 811
rect 2946 808 3158 811
rect 3170 808 3254 811
rect 3258 808 3478 811
rect 3514 808 3518 811
rect 3594 808 3630 811
rect 3706 808 3822 811
rect 3834 808 4046 811
rect 4242 808 4374 811
rect 496 803 498 807
rect 502 803 505 807
rect 510 803 512 807
rect 1520 803 1522 807
rect 1526 803 1529 807
rect 1534 803 1536 807
rect 2544 803 2546 807
rect 2550 803 2553 807
rect 2558 803 2560 807
rect 3568 803 3570 807
rect 3574 803 3577 807
rect 3582 803 3584 807
rect 74 798 318 801
rect 586 798 1078 801
rect 1882 798 1886 801
rect 1898 798 2054 801
rect 2122 798 2318 801
rect 2322 798 2382 801
rect 2386 798 2518 801
rect 2570 798 2582 801
rect 2626 798 2686 801
rect 2690 798 3166 801
rect 3234 798 3238 801
rect 3274 798 3350 801
rect 3410 798 3542 801
rect 3642 798 3686 801
rect 3814 798 3830 801
rect 3842 798 4134 801
rect 234 788 302 791
rect 962 788 1598 791
rect 1602 788 2294 791
rect 2354 788 2382 791
rect 2418 788 2614 791
rect 2706 788 2766 791
rect 2826 788 2894 791
rect 2938 788 2974 791
rect 2986 788 2990 791
rect 3086 788 3094 791
rect 3098 788 3214 791
rect 3218 788 3398 791
rect 3814 791 3817 798
rect 3522 788 3817 791
rect 3826 788 3830 791
rect 3914 788 3950 791
rect 3978 788 3982 791
rect 4050 788 4118 791
rect 4130 788 4286 791
rect 4306 788 4318 791
rect 566 781 569 788
rect 314 778 569 781
rect 1698 778 1806 781
rect 1810 778 2070 781
rect 2162 778 2166 781
rect 2382 781 2385 788
rect 2382 778 2502 781
rect 2538 778 2574 781
rect 2658 778 2846 781
rect 2850 778 3014 781
rect 3018 778 3054 781
rect 3058 778 4166 781
rect 4210 778 4214 781
rect 302 771 305 778
rect 678 772 681 778
rect 302 768 318 771
rect 562 768 630 771
rect 1162 768 1270 771
rect 1346 768 1366 771
rect 1490 768 1518 771
rect 1522 768 1550 771
rect 1634 768 1830 771
rect 1834 768 2014 771
rect 2018 768 2190 771
rect 2194 768 2262 771
rect 2314 768 2430 771
rect 2482 768 2566 771
rect 2594 768 2598 771
rect 2650 768 2750 771
rect 2786 768 2846 771
rect 2882 768 2926 771
rect 2934 768 3238 771
rect 3242 768 3246 771
rect 3298 768 3318 771
rect 3378 768 3502 771
rect 3570 768 3726 771
rect 4198 771 4201 778
rect 4010 768 4113 771
rect 4198 768 4206 771
rect 4262 771 4265 778
rect 4242 768 4265 771
rect 4382 771 4385 778
rect 4382 768 4414 771
rect 4426 768 4470 771
rect 4522 768 4542 771
rect 134 761 137 768
rect 134 758 142 761
rect 290 758 310 761
rect 434 758 446 761
rect 474 758 702 761
rect 714 758 766 761
rect 1210 758 1350 761
rect 1470 761 1473 768
rect 2934 762 2937 768
rect 4110 762 4113 768
rect 1378 758 1473 761
rect 1722 758 1753 761
rect 1778 758 1790 761
rect 1818 758 1822 761
rect 1902 758 1966 761
rect 2258 758 2358 761
rect 2362 758 2486 761
rect 2562 758 2614 761
rect 2642 758 2654 761
rect 2674 758 2726 761
rect 2810 758 2902 761
rect 2962 758 2966 761
rect 2978 758 3110 761
rect 3122 758 3134 761
rect 3186 758 3190 761
rect 3194 758 3214 761
rect 3226 758 3254 761
rect 3258 758 3302 761
rect 3306 758 3398 761
rect 3418 758 3422 761
rect 3442 758 3462 761
rect 3506 758 3678 761
rect 3722 758 3750 761
rect 3778 758 3782 761
rect 3834 758 3838 761
rect 3858 758 3886 761
rect 4010 758 4014 761
rect 4170 758 4238 761
rect 4242 758 4454 761
rect 366 752 369 758
rect 1566 752 1569 758
rect 146 748 174 751
rect 370 748 526 751
rect 578 748 582 751
rect 642 748 670 751
rect 754 748 870 751
rect 1098 748 1254 751
rect 1378 748 1422 751
rect 1606 751 1609 758
rect 1750 752 1753 758
rect 1902 752 1905 758
rect 1602 748 1609 751
rect 1658 748 1726 751
rect 1730 748 1742 751
rect 1770 748 1822 751
rect 1826 748 1846 751
rect 1930 748 1934 751
rect 1938 748 1974 751
rect 1978 748 1990 751
rect 2114 748 2126 751
rect 2146 748 2174 751
rect 2222 751 2225 758
rect 2486 752 2489 758
rect 2734 752 2737 758
rect 2202 748 2225 751
rect 2274 748 2278 751
rect 2314 748 2326 751
rect 2442 748 2470 751
rect 2530 748 2550 751
rect 2594 748 2662 751
rect 2682 748 2726 751
rect 2786 748 2790 751
rect 2866 748 2870 751
rect 2898 748 2926 751
rect 2938 748 2990 751
rect 3042 748 3198 751
rect 3210 748 3262 751
rect 3298 748 3342 751
rect 3362 748 3366 751
rect 3378 748 3382 751
rect 3430 751 3433 758
rect 3402 748 3433 751
rect 3466 748 3510 751
rect 3602 748 3606 751
rect 3618 748 3622 751
rect 3698 748 3702 751
rect 3746 748 3798 751
rect 3826 748 3958 751
rect 4010 748 4014 751
rect 1254 742 1257 748
rect 1878 742 1881 748
rect 2886 742 2889 748
rect 3278 742 3281 748
rect 3438 742 3441 748
rect 4022 742 4025 748
rect 4030 742 4033 751
rect 4162 748 4182 751
rect 4218 748 4438 751
rect 4442 748 4534 751
rect 4110 742 4113 748
rect 154 738 158 741
rect 162 738 182 741
rect 186 738 198 741
rect 202 738 206 741
rect 226 738 262 741
rect 322 738 358 741
rect 362 738 454 741
rect 458 738 502 741
rect 706 738 734 741
rect 738 738 750 741
rect 754 738 766 741
rect 1074 738 1150 741
rect 1154 738 1158 741
rect 1178 738 1246 741
rect 1346 738 1430 741
rect 1610 738 1622 741
rect 1650 738 1662 741
rect 1666 738 1678 741
rect 1770 738 1774 741
rect 1794 738 1830 741
rect 2106 738 2134 741
rect 2138 738 2150 741
rect 2154 738 2182 741
rect 2218 738 2238 741
rect 2242 738 2254 741
rect 2330 738 2334 741
rect 2354 738 2390 741
rect 2418 738 2622 741
rect 2666 738 2670 741
rect 2714 738 2734 741
rect 2794 738 2798 741
rect 2858 738 2862 741
rect 2938 738 2942 741
rect 3074 738 3102 741
rect 3106 738 3134 741
rect 3138 738 3150 741
rect 3186 738 3270 741
rect 3322 738 3390 741
rect 3426 738 3430 741
rect 3466 738 3558 741
rect 3578 738 3598 741
rect 3602 738 3726 741
rect 3754 738 3782 741
rect 3786 738 3798 741
rect 3802 738 3838 741
rect 3842 738 3910 741
rect 4066 738 4070 741
rect 4114 738 4142 741
rect 4146 738 4190 741
rect 4218 738 4246 741
rect 4266 738 4286 741
rect 4322 738 4358 741
rect 4386 738 4390 741
rect 4410 738 4438 741
rect 4474 738 4545 741
rect 2694 732 2697 738
rect 146 728 166 731
rect 202 728 302 731
rect 306 728 425 731
rect 1090 728 1198 731
rect 1202 728 1222 731
rect 1250 728 1342 731
rect 1506 728 1550 731
rect 1554 728 1574 731
rect 1674 728 1726 731
rect 1754 728 1854 731
rect 1858 728 2030 731
rect 2034 728 2166 731
rect 2170 728 2190 731
rect 2218 728 2238 731
rect 2290 728 2398 731
rect 2426 728 2438 731
rect 2458 728 2494 731
rect 2618 728 2662 731
rect 2810 728 2918 731
rect 2994 728 2998 731
rect 3030 731 3033 738
rect 3010 728 3033 731
rect 3042 728 3054 731
rect 3114 728 3118 731
rect 3122 728 3150 731
rect 3178 728 3206 731
rect 3226 728 3246 731
rect 3274 728 3286 731
rect 3346 728 3462 731
rect 3474 728 3622 731
rect 3642 728 3673 731
rect 3778 728 3854 731
rect 3926 731 3929 738
rect 4542 732 4545 738
rect 3922 728 4046 731
rect 4050 728 4054 731
rect 4130 728 4134 731
rect 4242 728 4294 731
rect 4354 728 4358 731
rect 4378 728 4385 731
rect 4402 728 4430 731
rect 4498 728 4526 731
rect 422 722 425 728
rect 1622 722 1625 728
rect 106 718 134 721
rect 186 718 230 721
rect 410 718 414 721
rect 434 718 750 721
rect 1026 718 1118 721
rect 1122 718 1214 721
rect 1290 718 1294 721
rect 1738 718 2054 721
rect 2058 718 2158 721
rect 2178 718 2182 721
rect 2510 721 2513 728
rect 3670 722 3673 728
rect 4342 722 4345 728
rect 4382 722 4385 728
rect 2510 718 2606 721
rect 2626 718 2694 721
rect 2810 718 2822 721
rect 2826 718 2862 721
rect 2938 718 3334 721
rect 3346 718 3478 721
rect 3490 718 3526 721
rect 3530 718 3590 721
rect 3594 718 3614 721
rect 3618 718 3670 721
rect 3698 718 3822 721
rect 3850 718 3854 721
rect 3898 718 4126 721
rect 4162 718 4294 721
rect 4482 718 4510 721
rect 4538 718 4574 721
rect 1398 712 1401 718
rect 178 708 342 711
rect 418 708 454 711
rect 458 708 558 711
rect 562 708 574 711
rect 586 708 638 711
rect 1034 708 1126 711
rect 1162 708 1174 711
rect 1210 708 1222 711
rect 1698 708 1734 711
rect 1738 708 1902 711
rect 1986 708 2006 711
rect 2122 708 2134 711
rect 2386 708 2414 711
rect 2498 708 2574 711
rect 2650 708 2678 711
rect 2802 708 2846 711
rect 2850 708 2894 711
rect 2914 708 3038 711
rect 3098 708 3134 711
rect 3146 708 3238 711
rect 3266 708 3294 711
rect 3330 708 3366 711
rect 3370 708 3438 711
rect 3442 708 3502 711
rect 3618 708 3798 711
rect 3834 708 3878 711
rect 4158 711 4161 718
rect 4106 708 4161 711
rect 4194 708 4462 711
rect 4466 708 4486 711
rect 4506 708 4542 711
rect 4546 708 4598 711
rect 1000 703 1002 707
rect 1006 703 1009 707
rect 1014 703 1016 707
rect 2024 703 2026 707
rect 2030 703 2033 707
rect 2038 703 2040 707
rect 2606 702 2609 708
rect 3048 703 3050 707
rect 3054 703 3057 707
rect 3062 703 3064 707
rect 3606 702 3609 708
rect 3806 702 3809 708
rect 4080 703 4082 707
rect 4086 703 4089 707
rect 4094 703 4096 707
rect 154 698 214 701
rect 410 698 438 701
rect 666 698 790 701
rect 1146 698 1238 701
rect 1306 698 1326 701
rect 1338 698 1398 701
rect 1442 698 1478 701
rect 1730 698 1798 701
rect 2122 698 2574 701
rect 2626 698 2734 701
rect 2746 698 2838 701
rect 2858 698 2982 701
rect 3138 698 3158 701
rect 3218 698 3230 701
rect 3238 698 3294 701
rect 3458 698 3478 701
rect 3506 698 3534 701
rect 4114 698 4166 701
rect 4314 698 4374 701
rect 4418 698 4422 701
rect 4426 698 4550 701
rect 1822 692 1825 698
rect 10 688 22 691
rect 26 688 126 691
rect 130 688 182 691
rect 226 688 294 691
rect 298 688 414 691
rect 634 688 654 691
rect 658 688 665 691
rect 674 688 830 691
rect 994 688 1014 691
rect 1050 688 1070 691
rect 1074 688 1182 691
rect 1290 688 1297 691
rect 1314 688 1630 691
rect 1682 688 1718 691
rect 1722 688 1766 691
rect 1770 688 1806 691
rect 1954 688 2014 691
rect 2018 688 2030 691
rect 2042 688 2046 691
rect 2370 688 2398 691
rect 2402 688 2422 691
rect 2498 688 2518 691
rect 2526 688 2622 691
rect 2690 688 2702 691
rect 2706 688 2718 691
rect 2778 688 2782 691
rect 2834 688 2910 691
rect 2922 688 3022 691
rect 3238 691 3241 698
rect 3162 688 3241 691
rect 3270 688 3582 691
rect 3662 688 3750 691
rect 3762 688 3814 691
rect 3818 688 3894 691
rect 3906 688 3990 691
rect 3994 688 4238 691
rect 4258 688 4289 691
rect 274 678 446 681
rect 450 678 478 681
rect 482 678 526 681
rect 538 678 550 681
rect 562 678 710 681
rect 1062 678 1190 681
rect 1242 678 1278 681
rect 206 671 209 678
rect 206 668 246 671
rect 250 668 278 671
rect 522 668 678 671
rect 682 668 790 671
rect 966 671 969 678
rect 1054 671 1057 678
rect 966 668 1057 671
rect 1062 672 1065 678
rect 1130 668 1198 671
rect 1294 671 1297 688
rect 1646 682 1649 688
rect 1306 678 1337 681
rect 1370 678 1382 681
rect 1690 678 1742 681
rect 1762 678 1782 681
rect 1786 678 1942 681
rect 1946 678 2014 681
rect 2018 678 2086 681
rect 2302 681 2305 688
rect 2302 678 2454 681
rect 2526 681 2529 688
rect 2514 678 2529 681
rect 2654 681 2657 688
rect 2654 678 2670 681
rect 2682 678 2718 681
rect 2722 678 2977 681
rect 3002 678 3006 681
rect 3030 681 3033 688
rect 3030 678 3070 681
rect 3142 681 3145 688
rect 3270 682 3273 688
rect 3662 682 3665 688
rect 4286 682 4289 688
rect 3082 678 3145 681
rect 3170 678 3174 681
rect 3370 678 3598 681
rect 3658 678 3662 681
rect 3714 678 3726 681
rect 3810 678 3902 681
rect 4034 678 4046 681
rect 4210 678 4262 681
rect 4366 681 4369 688
rect 4298 678 4446 681
rect 4562 678 4566 681
rect 1334 672 1337 678
rect 1294 668 1318 671
rect 1346 668 1358 671
rect 1494 671 1497 678
rect 1614 672 1617 678
rect 1466 668 1497 671
rect 1570 668 1606 671
rect 1634 668 1638 671
rect 1658 668 1734 671
rect 1858 668 1886 671
rect 2098 668 2174 671
rect 2194 668 2198 671
rect 2218 668 2222 671
rect 2274 668 2278 671
rect 2290 668 2294 671
rect 2346 668 2358 671
rect 2582 671 2585 678
rect 2974 672 2977 678
rect 3358 672 3361 678
rect 2554 668 2798 671
rect 2890 668 2934 671
rect 2982 668 3014 671
rect 3018 668 3062 671
rect 3066 668 3102 671
rect 3138 668 3206 671
rect 3226 668 3286 671
rect 3290 668 3326 671
rect 3426 668 3430 671
rect 3434 668 3478 671
rect 3602 668 3670 671
rect 3674 668 3718 671
rect 3722 668 3766 671
rect 3802 668 3854 671
rect 3858 668 3886 671
rect 3890 668 3950 671
rect 3962 668 4038 671
rect 4070 671 4073 678
rect 4070 668 4102 671
rect 4158 671 4161 678
rect 4154 668 4161 671
rect 4178 668 4182 671
rect 4234 668 4238 671
rect 4250 668 4254 671
rect 4346 668 4366 671
rect 4370 668 4374 671
rect 4498 668 4526 671
rect 90 659 142 661
rect 86 658 142 659
rect 186 658 238 661
rect 306 658 310 661
rect 370 658 478 661
rect 526 658 593 661
rect 706 658 750 661
rect 894 661 897 668
rect 810 658 897 661
rect 1122 658 1161 661
rect 1178 658 1206 661
rect 1422 661 1425 668
rect 1386 658 1425 661
rect 1578 658 1598 661
rect 1626 658 1630 661
rect 1642 658 1646 661
rect 1750 661 1753 668
rect 1846 662 1849 668
rect 1750 658 1774 661
rect 1850 658 1910 661
rect 2034 658 2070 661
rect 2106 658 2110 661
rect 2130 658 2142 661
rect 2146 658 2158 661
rect 2202 658 2278 661
rect 2282 658 2326 661
rect 2330 658 2430 661
rect 2490 658 2494 661
rect 2522 658 2566 661
rect 2634 658 2702 661
rect 2706 658 2726 661
rect 2786 658 2790 661
rect 2870 661 2873 668
rect 2818 658 2873 661
rect 2982 661 2985 668
rect 2930 658 2985 661
rect 3010 658 3070 661
rect 3106 658 3142 661
rect 3170 658 3182 661
rect 3266 658 3318 661
rect 3354 658 3382 661
rect 3386 658 3414 661
rect 3418 658 3510 661
rect 3546 658 3678 661
rect 3690 658 3798 661
rect 3986 658 3998 661
rect 4002 658 4054 661
rect 4186 658 4190 661
rect 4194 658 4278 661
rect 4314 658 4406 661
rect 4410 658 4422 661
rect 4490 658 4502 661
rect 4530 658 4590 661
rect 526 652 529 658
rect 590 652 593 658
rect 1158 652 1161 658
rect -26 651 -22 652
rect -26 648 6 651
rect 34 648 134 651
rect 162 648 190 651
rect 242 648 246 651
rect 318 648 326 651
rect 330 648 342 651
rect 346 648 401 651
rect 618 648 654 651
rect 658 648 686 651
rect 726 648 734 651
rect 738 648 750 651
rect 754 648 902 651
rect 1162 648 1302 651
rect 1410 648 1430 651
rect 1826 648 1870 651
rect 1890 648 1926 651
rect 1934 651 1937 658
rect 2006 652 2009 658
rect 1934 648 1950 651
rect 2066 648 2174 651
rect 2178 648 2230 651
rect 2298 648 2382 651
rect 2490 648 2606 651
rect 2610 648 2654 651
rect 2714 648 2750 651
rect 2770 648 2782 651
rect 2786 648 2822 651
rect 2830 648 3006 651
rect 3010 648 3046 651
rect 3274 648 3406 651
rect 3474 648 3486 651
rect 3610 648 3630 651
rect 3666 648 3670 651
rect 3722 648 3814 651
rect 3818 648 3838 651
rect 4002 648 4014 651
rect 4042 648 4102 651
rect 4122 648 4246 651
rect 4322 648 4438 651
rect 4458 648 4478 651
rect 286 641 289 648
rect 398 642 401 648
rect 266 638 342 641
rect 362 638 390 641
rect 410 638 526 641
rect 546 638 745 641
rect 1274 638 1390 641
rect 1718 641 1721 648
rect 2830 642 2833 648
rect 3126 642 3129 648
rect 3182 642 3185 648
rect 3398 642 3401 648
rect 1718 638 1766 641
rect 1874 638 2158 641
rect 2418 638 2494 641
rect 2618 638 2726 641
rect 2938 638 3022 641
rect 3026 638 3078 641
rect 3282 638 3286 641
rect 3482 638 3614 641
rect 3626 638 3726 641
rect 3738 638 3862 641
rect 3902 641 3905 648
rect 3866 638 3905 641
rect 3922 638 4118 641
rect 4122 638 4206 641
rect 4274 638 4310 641
rect 4354 638 4430 641
rect 4434 638 4494 641
rect 254 632 257 638
rect 742 632 745 638
rect 370 628 646 631
rect 658 628 670 631
rect 1274 628 1606 631
rect 1610 628 1862 631
rect 1882 628 1950 631
rect 2018 628 2094 631
rect 2298 628 4070 631
rect 4222 628 4334 631
rect 4354 628 4414 631
rect 170 618 254 621
rect 282 618 982 621
rect 1098 618 1102 621
rect 1138 618 1286 621
rect 1330 618 1558 621
rect 1562 618 1758 621
rect 1794 618 1798 621
rect 1866 618 1926 621
rect 2066 618 2150 621
rect 2242 618 2790 621
rect 2834 618 2870 621
rect 2946 618 2958 621
rect 2994 618 3182 621
rect 3226 618 3310 621
rect 3314 618 3334 621
rect 3402 618 3550 621
rect 3666 618 3822 621
rect 3858 618 3998 621
rect 4014 618 4022 621
rect 4026 618 4214 621
rect 4222 621 4225 628
rect 4218 618 4225 621
rect 4234 618 4398 621
rect 4402 618 4470 621
rect 4522 618 4574 621
rect 746 608 1150 611
rect 1938 608 2126 611
rect 2130 608 2238 611
rect 2258 608 2422 611
rect 2458 608 2478 611
rect 2482 608 2518 611
rect 2578 608 2910 611
rect 2954 608 3206 611
rect 3210 608 3334 611
rect 3682 608 3686 611
rect 3770 608 3934 611
rect 3938 608 3974 611
rect 4018 608 4142 611
rect 4146 608 4166 611
rect 4186 608 4382 611
rect 4386 608 4574 611
rect 496 603 498 607
rect 502 603 505 607
rect 510 603 512 607
rect 1520 603 1522 607
rect 1526 603 1529 607
rect 1534 603 1536 607
rect 2544 603 2546 607
rect 2550 603 2553 607
rect 2558 603 2560 607
rect 3568 603 3570 607
rect 3574 603 3577 607
rect 3582 603 3584 607
rect 394 598 422 601
rect 650 598 654 601
rect 762 598 894 601
rect 906 598 950 601
rect 1834 598 1902 601
rect 1906 598 1958 601
rect 1962 598 1974 601
rect 2442 598 2534 601
rect 2658 598 2662 601
rect 2666 598 2838 601
rect 2914 598 3022 601
rect 3082 598 3102 601
rect 3146 598 3190 601
rect 3194 598 3326 601
rect 3682 598 3790 601
rect 3866 598 3870 601
rect 3978 598 4206 601
rect 4210 598 4214 601
rect 4218 598 4486 601
rect 4490 598 4558 601
rect 2126 592 2129 598
rect 390 588 1126 591
rect 1490 588 1494 591
rect 2474 588 2606 591
rect 2666 588 2774 591
rect 3018 588 3030 591
rect 3242 588 3302 591
rect 3318 588 3446 591
rect 3454 588 3702 591
rect 4034 588 4062 591
rect 4074 588 4190 591
rect 4194 588 4318 591
rect 4458 588 4486 591
rect 390 582 393 588
rect 146 578 174 581
rect 658 578 1070 581
rect 1394 578 1398 581
rect 1470 581 1473 588
rect 2990 582 2993 588
rect 3318 582 3321 588
rect 3454 582 3457 588
rect 1402 578 1473 581
rect 1706 578 2086 581
rect 2138 578 2142 581
rect 2354 578 2462 581
rect 2466 578 2606 581
rect 2610 578 2630 581
rect 2730 578 2854 581
rect 2858 578 2902 581
rect 3002 578 3086 581
rect 3090 578 3094 581
rect 3130 578 3134 581
rect 3226 578 3238 581
rect 3602 578 3702 581
rect 3858 578 3878 581
rect 3930 578 4150 581
rect 4154 578 4222 581
rect 4242 578 4326 581
rect 4506 578 4561 581
rect -26 571 -22 572
rect 30 571 33 578
rect -26 568 33 571
rect 786 568 790 571
rect 798 568 846 571
rect 1002 568 1262 571
rect 1338 568 1382 571
rect 1386 568 1438 571
rect 1442 568 1470 571
rect 1514 568 1558 571
rect 1658 568 1702 571
rect 1794 568 1822 571
rect 1898 568 1910 571
rect 1914 568 2150 571
rect 2194 568 2254 571
rect 2266 568 2345 571
rect 2394 568 2430 571
rect 2434 568 2462 571
rect 2762 568 2814 571
rect 2818 568 2822 571
rect 2834 568 2870 571
rect 2906 568 2990 571
rect 3026 568 3374 571
rect 3394 568 3670 571
rect 3698 568 3702 571
rect 3714 568 3742 571
rect 3746 568 3838 571
rect 3858 568 4198 571
rect 4282 568 4302 571
rect 4390 571 4393 578
rect 4558 572 4561 578
rect 4314 568 4393 571
rect 4410 568 4462 571
rect 4466 568 4550 571
rect 258 558 326 561
rect 662 561 665 568
rect 798 562 801 568
rect 2342 562 2345 568
rect 642 558 694 561
rect 738 558 782 561
rect 830 558 838 561
rect 842 558 878 561
rect 902 558 998 561
rect 1130 558 1598 561
rect 1602 558 1654 561
rect 1738 558 1750 561
rect 1818 558 2014 561
rect 2026 558 2070 561
rect 2266 558 2270 561
rect 2278 558 2286 561
rect 2290 558 2318 561
rect 2378 558 2502 561
rect 2506 558 2574 561
rect 2590 561 2593 568
rect 2578 558 2593 561
rect 2602 558 2646 561
rect 2738 558 2742 561
rect 2746 558 2774 561
rect 3006 561 3009 568
rect 2970 558 3014 561
rect 3026 558 3046 561
rect 3106 558 3190 561
rect 3194 558 3198 561
rect 3210 558 3262 561
rect 3266 558 3270 561
rect 3418 558 3470 561
rect 3474 558 3494 561
rect 3498 558 3534 561
rect 3538 558 3542 561
rect 3594 558 3598 561
rect 3618 558 3622 561
rect 3670 561 3673 568
rect 3670 558 3766 561
rect 3770 558 3782 561
rect 3794 558 3830 561
rect 3874 558 3902 561
rect 3906 558 3958 561
rect 3970 558 4390 561
rect 4394 558 4526 561
rect 4558 561 4561 568
rect 4558 558 4574 561
rect -26 551 -22 552
rect -26 548 6 551
rect 114 548 278 551
rect 358 551 361 558
rect 902 552 905 558
rect 1694 552 1697 558
rect 2118 552 2121 558
rect 358 548 454 551
rect 530 548 742 551
rect 1138 548 1166 551
rect 1498 548 1518 551
rect 1522 548 1582 551
rect 1650 548 1694 551
rect 1698 548 1702 551
rect 1706 548 1718 551
rect 1722 548 1774 551
rect 1778 548 1782 551
rect 1874 548 1878 551
rect 1894 548 1982 551
rect 1986 548 1990 551
rect 2018 548 2118 551
rect 2702 551 2705 558
rect 2122 548 2705 551
rect 2802 548 2806 551
rect 2882 548 2886 551
rect 2954 548 2958 551
rect 3050 548 3070 551
rect 3122 548 3158 551
rect 3194 548 3246 551
rect 3274 548 3302 551
rect 3410 548 3422 551
rect 3482 548 3606 551
rect 3714 548 3734 551
rect 3782 548 3814 551
rect 3842 548 3854 551
rect 3986 548 4030 551
rect 4038 548 4046 551
rect 4050 548 4062 551
rect 4082 548 4086 551
rect 4122 548 4126 551
rect 4258 548 4286 551
rect 4290 548 4382 551
rect 4410 548 4438 551
rect 4442 548 4454 551
rect 4514 548 4518 551
rect 4554 548 4582 551
rect 310 541 313 548
rect 210 538 313 541
rect 454 541 457 548
rect 942 542 945 548
rect 454 538 577 541
rect 778 538 798 541
rect 802 538 902 541
rect 970 538 1102 541
rect 1106 538 1222 541
rect 1414 541 1417 548
rect 1226 538 1249 541
rect 1414 538 1422 541
rect 1426 538 1614 541
rect 1690 538 1718 541
rect 1722 538 1726 541
rect 1850 538 1862 541
rect 1894 541 1897 548
rect 3782 542 3785 548
rect 3822 542 3825 548
rect 4158 542 4161 548
rect 1866 538 1897 541
rect 2106 538 2110 541
rect 2266 538 2270 541
rect 2346 538 2374 541
rect 2386 538 2438 541
rect 2546 538 2582 541
rect 2586 538 2630 541
rect 2634 538 2638 541
rect 2658 538 2670 541
rect 2674 538 2734 541
rect 2778 538 2806 541
rect 2810 538 2846 541
rect 2874 538 2902 541
rect 2906 538 3038 541
rect 3042 538 3070 541
rect 3074 538 3094 541
rect 3122 538 3126 541
rect 3234 538 3238 541
rect 3258 538 3318 541
rect 3402 538 3406 541
rect 3458 538 3486 541
rect 3490 538 3502 541
rect 3546 538 3598 541
rect 3850 538 3934 541
rect 3938 538 3942 541
rect 3954 538 4038 541
rect 4058 538 4094 541
rect 4130 538 4134 541
rect 4198 538 4214 541
rect 4298 538 4478 541
rect 4570 538 4574 541
rect 574 532 577 538
rect 1246 532 1249 538
rect 1322 528 1326 531
rect 1330 528 1366 531
rect 1418 528 1478 531
rect 1490 528 1574 531
rect 1650 528 1654 531
rect 1786 528 1830 531
rect 1834 528 1838 531
rect 1842 528 1854 531
rect 1898 528 1910 531
rect 1938 528 1942 531
rect 1946 528 1974 531
rect 2054 531 2057 538
rect 2230 532 2233 538
rect 3110 532 3113 538
rect 4198 532 4201 538
rect 1994 528 2057 531
rect 2066 528 2070 531
rect 2178 528 2190 531
rect 2286 528 2385 531
rect 2410 528 2494 531
rect 2498 528 2534 531
rect 2578 528 2614 531
rect 2618 528 2638 531
rect 2790 528 2798 531
rect 2906 528 2982 531
rect 3186 528 3206 531
rect 3210 528 3350 531
rect 3354 528 3390 531
rect 3418 528 3430 531
rect 3586 528 3662 531
rect 3666 528 3718 531
rect 3802 528 3878 531
rect 3890 528 3918 531
rect 3930 528 3974 531
rect 3994 528 4022 531
rect 4058 528 4134 531
rect 4146 528 4158 531
rect 4250 528 4294 531
rect 4322 528 4374 531
rect 4378 528 4462 531
rect 4466 528 4510 531
rect 4538 528 4558 531
rect 1142 522 1145 528
rect 330 518 406 521
rect 410 518 862 521
rect 1218 518 1502 521
rect 1946 518 2006 521
rect 2010 518 2046 521
rect 2222 521 2225 528
rect 2286 522 2289 528
rect 2382 522 2385 528
rect 2222 518 2278 521
rect 2450 518 2526 521
rect 2546 518 2574 521
rect 2794 518 2886 521
rect 2938 518 2942 521
rect 2978 518 3174 521
rect 3194 518 3206 521
rect 3298 518 3358 521
rect 3726 521 3729 528
rect 3726 518 3934 521
rect 3946 518 3990 521
rect 3994 518 3998 521
rect 4070 518 4246 521
rect 4250 518 4262 521
rect 4274 518 4446 521
rect 1854 512 1857 518
rect 2598 512 2601 518
rect 3182 512 3185 518
rect 514 508 542 511
rect 562 508 590 511
rect 1386 508 1422 511
rect 1474 508 1550 511
rect 1554 508 1614 511
rect 1922 508 1934 511
rect 2082 508 2214 511
rect 2226 508 2254 511
rect 2274 508 2326 511
rect 2330 508 2414 511
rect 2474 508 2590 511
rect 2610 508 2630 511
rect 2634 508 2678 511
rect 2706 508 2822 511
rect 3346 508 3358 511
rect 3546 508 3758 511
rect 3810 508 3942 511
rect 4070 511 4073 518
rect 3954 508 4073 511
rect 4298 508 4366 511
rect 4434 508 4470 511
rect 1000 503 1002 507
rect 1006 503 1009 507
rect 1014 503 1016 507
rect 1430 502 1433 508
rect 2024 503 2026 507
rect 2030 503 2033 507
rect 2038 503 2040 507
rect 3048 503 3050 507
rect 3054 503 3057 507
rect 3062 503 3064 507
rect 3422 502 3425 508
rect 4080 503 4082 507
rect 4086 503 4089 507
rect 4094 503 4096 507
rect 202 498 270 501
rect 274 498 310 501
rect 338 498 598 501
rect 602 498 814 501
rect 1282 498 1342 501
rect 1346 498 1390 501
rect 1490 498 1654 501
rect 1674 498 1910 501
rect 2098 498 2190 501
rect 2242 498 2478 501
rect 2490 498 2502 501
rect 2514 498 2566 501
rect 2570 498 2606 501
rect 2610 498 2662 501
rect 2674 498 2710 501
rect 2722 498 2790 501
rect 2826 498 2942 501
rect 3090 498 3374 501
rect 3434 498 3470 501
rect 3634 498 3894 501
rect 3898 498 3910 501
rect 3914 498 3974 501
rect 3978 498 4006 501
rect 4018 498 4062 501
rect 4154 498 4158 501
rect 4162 498 4174 501
rect 4402 498 4414 501
rect 4458 498 4550 501
rect 266 488 294 491
rect 490 488 558 491
rect 674 488 710 491
rect 714 488 774 491
rect 778 488 942 491
rect 1210 488 1630 491
rect 2010 488 2030 491
rect 2050 488 2070 491
rect 2162 488 2166 491
rect 2170 488 2182 491
rect 2226 488 2238 491
rect 2242 488 2310 491
rect 2370 488 2406 491
rect 2418 488 2662 491
rect 2674 488 2686 491
rect 2698 488 2814 491
rect 2862 488 2870 491
rect 2874 488 2894 491
rect 3122 488 3249 491
rect 274 478 278 481
rect 538 478 630 481
rect 634 478 726 481
rect 882 478 934 481
rect 1418 478 1486 481
rect 1642 478 1646 481
rect 1666 478 1694 481
rect 1782 481 1785 488
rect 1738 478 1785 481
rect 1998 481 2001 488
rect 3246 482 3249 488
rect 3298 488 3310 491
rect 3398 491 3401 498
rect 3362 488 3401 491
rect 3410 488 3462 491
rect 3498 488 3502 491
rect 3506 488 3622 491
rect 3806 488 3814 491
rect 3858 488 3878 491
rect 3890 488 3982 491
rect 4002 488 4054 491
rect 4106 488 4174 491
rect 4178 488 4238 491
rect 4358 488 4366 491
rect 4370 488 4382 491
rect 4386 488 4414 491
rect 4418 488 4462 491
rect 1898 478 2001 481
rect 2066 478 2110 481
rect 2178 478 2358 481
rect 2386 478 2454 481
rect 2458 478 2470 481
rect 2474 478 2582 481
rect 2586 478 2718 481
rect 2762 478 2774 481
rect 2850 478 2918 481
rect 2954 478 3030 481
rect 3074 478 3126 481
rect 3178 478 3230 481
rect 3294 481 3297 488
rect 3742 482 3745 488
rect 3806 482 3809 488
rect 3258 478 3297 481
rect 3322 478 3438 481
rect 3458 478 3510 481
rect 3746 478 3758 481
rect 3834 478 3862 481
rect 3878 481 3881 488
rect 3878 478 3910 481
rect 3982 481 3985 488
rect 3982 478 4054 481
rect 4066 478 4126 481
rect 4202 478 4254 481
rect 4314 478 4326 481
rect 4354 478 4401 481
rect 4502 481 4505 488
rect 4426 478 4505 481
rect 4522 478 4542 481
rect 390 472 393 478
rect 226 468 246 471
rect 250 468 318 471
rect 482 468 566 471
rect 730 468 742 471
rect 898 468 950 471
rect 954 468 958 471
rect 1326 471 1329 478
rect 1034 468 1097 471
rect 1326 468 1334 471
rect 1382 471 1385 478
rect 1614 472 1617 478
rect 1790 472 1793 478
rect 1382 468 1510 471
rect 1634 468 1638 471
rect 1666 468 1718 471
rect 1722 468 1766 471
rect 1834 468 1886 471
rect 2022 471 2025 478
rect 2822 472 2825 478
rect 2022 468 2054 471
rect 2106 468 2118 471
rect 2158 468 2214 471
rect 2282 468 2342 471
rect 2354 468 2398 471
rect 2410 468 2414 471
rect 2458 468 2462 471
rect 2498 468 2502 471
rect 2514 468 2542 471
rect 2586 468 2606 471
rect 2658 468 2710 471
rect 2834 468 2838 471
rect 2858 468 2862 471
rect 2898 468 2902 471
rect 2950 471 2953 478
rect 4398 472 4401 478
rect 4574 472 4577 478
rect 2938 468 2953 471
rect 2962 468 2974 471
rect 3018 468 3086 471
rect 3090 468 3134 471
rect 3138 468 3174 471
rect 3298 468 3350 471
rect 3354 468 3422 471
rect 3434 468 3622 471
rect 3818 468 3846 471
rect 3882 468 3998 471
rect 4002 468 4006 471
rect 4010 468 4022 471
rect 4034 468 4038 471
rect 4058 468 4110 471
rect 4122 468 4142 471
rect 4338 468 4342 471
rect 4402 468 4574 471
rect 366 462 369 468
rect 1094 462 1097 468
rect 26 458 57 461
rect 90 458 166 461
rect 170 458 206 461
rect 258 458 262 461
rect 266 458 302 461
rect 306 458 366 461
rect 626 458 649 461
rect 682 458 694 461
rect 698 458 702 461
rect 794 458 798 461
rect 802 458 886 461
rect 1338 458 1438 461
rect 1442 458 1449 461
rect 1518 461 1521 468
rect 1458 458 1521 461
rect 1614 461 1617 468
rect 1766 462 1769 468
rect 1614 458 1670 461
rect 1674 458 1678 461
rect 1690 458 1718 461
rect 1722 458 1734 461
rect 1810 458 1814 461
rect 1850 458 1862 461
rect 1934 461 1937 468
rect 2158 462 2161 468
rect 1934 458 1966 461
rect 1978 458 1982 461
rect 2230 461 2233 468
rect 2782 462 2785 468
rect 3854 462 3857 468
rect 2230 458 2238 461
rect 2258 458 2294 461
rect 2362 458 2438 461
rect 2442 458 2582 461
rect 2602 458 2641 461
rect 2650 458 2758 461
rect 2882 458 2886 461
rect 2946 458 2966 461
rect 3034 458 3062 461
rect 3098 458 3254 461
rect 3274 458 3302 461
rect 3306 458 3342 461
rect 3346 458 3353 461
rect 3362 458 3430 461
rect 3442 458 3462 461
rect 3490 458 3558 461
rect 3562 458 3598 461
rect 3602 458 3646 461
rect 3650 458 3678 461
rect 3682 458 3710 461
rect 3714 458 3742 461
rect 3922 458 3942 461
rect 3962 458 4294 461
rect 4306 458 4318 461
rect 4322 458 4350 461
rect 4362 458 4398 461
rect 4466 458 4470 461
rect 4498 458 4518 461
rect 4538 458 4558 461
rect 54 452 57 458
rect 646 452 649 458
rect 1206 452 1209 458
rect 1606 452 1609 458
rect 2118 452 2121 458
rect -26 451 -22 452
rect -26 448 6 451
rect 58 448 126 451
rect 194 448 230 451
rect 242 448 294 451
rect 610 448 638 451
rect 690 448 702 451
rect 770 448 878 451
rect 1426 448 1438 451
rect 1650 448 1894 451
rect 1954 448 2006 451
rect 2010 448 2046 451
rect 2050 448 2070 451
rect 2122 448 2174 451
rect 2178 448 2198 451
rect 2202 448 2214 451
rect 2242 448 2262 451
rect 2266 448 2270 451
rect 2322 448 2622 451
rect 2626 448 2630 451
rect 2638 451 2641 458
rect 2638 448 2670 451
rect 2714 448 2718 451
rect 2802 448 2806 451
rect 2974 448 2982 451
rect 2986 448 3038 451
rect 3074 448 3110 451
rect 3130 448 3134 451
rect 3194 448 3222 451
rect 3234 448 3262 451
rect 3298 448 3302 451
rect 3458 448 3662 451
rect 3674 448 3678 451
rect 3690 448 3694 451
rect 3698 448 3782 451
rect 3934 448 3950 451
rect 3970 448 4206 451
rect 4282 448 4422 451
rect 4426 448 4457 451
rect 4466 448 4510 451
rect 4514 448 4534 451
rect 130 438 286 441
rect 302 441 305 448
rect 298 438 350 441
rect 582 441 585 448
rect 702 442 705 448
rect 582 438 590 441
rect 674 438 678 441
rect 894 441 897 448
rect 2942 442 2945 448
rect 2974 442 2977 448
rect 3406 442 3409 448
rect 3822 442 3825 448
rect 3830 442 3833 448
rect 3934 442 3937 448
rect 894 438 910 441
rect 986 438 1070 441
rect 1074 438 1110 441
rect 1170 438 1246 441
rect 1250 438 1294 441
rect 1754 438 2382 441
rect 2386 438 2598 441
rect 2602 438 2662 441
rect 2706 438 2734 441
rect 2738 438 2830 441
rect 2834 438 2878 441
rect 3026 438 3230 441
rect 3234 438 3310 441
rect 3314 438 3318 441
rect 3522 438 3526 441
rect 3706 438 3798 441
rect 3850 438 3913 441
rect 3958 441 3961 448
rect 4238 442 4241 448
rect 3958 438 4022 441
rect 4042 438 4182 441
rect 4186 438 4190 441
rect 4314 438 4318 441
rect 4322 438 4366 441
rect 4370 438 4438 441
rect 4454 441 4457 448
rect 4454 438 4478 441
rect 4554 438 4558 441
rect 242 428 273 431
rect 354 428 406 431
rect 698 428 702 431
rect 706 428 710 431
rect 1170 428 1438 431
rect 1442 428 1454 431
rect 1466 428 1598 431
rect 1602 428 1854 431
rect 1874 428 1878 431
rect 2010 428 2014 431
rect 2194 428 2414 431
rect 2426 428 2430 431
rect 2506 428 2534 431
rect 2546 428 2622 431
rect 2754 428 2806 431
rect 2970 428 3014 431
rect 3042 428 3670 431
rect 3722 428 3902 431
rect 3910 431 3913 438
rect 3910 428 4334 431
rect 270 422 273 428
rect 378 418 606 421
rect 626 418 1305 421
rect 1322 418 1350 421
rect 1546 418 1686 421
rect 1802 418 2118 421
rect 2234 418 2526 421
rect 2530 418 2702 421
rect 2770 418 3102 421
rect 3162 418 3198 421
rect 3506 418 3606 421
rect 3706 418 3758 421
rect 3770 418 4310 421
rect 4314 418 4337 421
rect 1302 412 1305 418
rect 266 408 486 411
rect 2018 408 2094 411
rect 2346 408 2478 411
rect 2650 408 2734 411
rect 2738 408 2750 411
rect 2922 408 3102 411
rect 3170 408 3238 411
rect 3738 408 3742 411
rect 3746 408 3814 411
rect 3850 408 3934 411
rect 3946 408 3958 411
rect 3962 408 4174 411
rect 4218 408 4262 411
rect 4334 411 4337 418
rect 4334 408 4390 411
rect 4394 408 4518 411
rect 496 403 498 407
rect 502 403 505 407
rect 510 403 512 407
rect 1520 403 1522 407
rect 1526 403 1529 407
rect 1534 403 1536 407
rect 1822 402 1825 408
rect 2544 403 2546 407
rect 2550 403 2553 407
rect 2558 403 2560 407
rect 3568 403 3570 407
rect 3574 403 3577 407
rect 3582 403 3584 407
rect 202 398 286 401
rect 330 398 374 401
rect 866 398 1134 401
rect 1370 398 1398 401
rect 1402 398 1454 401
rect 2082 398 2318 401
rect 2330 398 2502 401
rect 2578 398 2678 401
rect 3082 398 3086 401
rect 3186 398 3198 401
rect 3210 398 3302 401
rect 3602 398 3606 401
rect 3614 398 3678 401
rect 3682 398 3950 401
rect 3970 398 3974 401
rect 4010 398 4038 401
rect 4050 398 4174 401
rect 4210 398 4334 401
rect 250 388 406 391
rect 410 388 462 391
rect 466 388 590 391
rect 610 388 1102 391
rect 1506 388 1526 391
rect 1762 388 2774 391
rect 3614 391 3617 398
rect 2818 388 3617 391
rect 3666 388 4278 391
rect 78 378 222 381
rect 562 378 590 381
rect 642 378 734 381
rect 738 378 742 381
rect 794 378 1006 381
rect 1010 378 1294 381
rect 1450 378 1494 381
rect 1498 378 1670 381
rect 1698 378 1934 381
rect 1986 378 2110 381
rect 2114 378 2190 381
rect 2194 378 2286 381
rect 2450 378 2558 381
rect 2562 378 2590 381
rect 2634 378 2654 381
rect 2666 378 2766 381
rect 2970 378 3150 381
rect 3162 378 3198 381
rect 3346 378 3374 381
rect 3378 378 3390 381
rect 3962 378 4070 381
rect 4074 378 4230 381
rect 78 372 81 378
rect 130 368 142 371
rect 146 368 310 371
rect 326 371 329 378
rect 3806 372 3809 378
rect 326 368 350 371
rect 426 368 622 371
rect 906 368 934 371
rect 1770 368 1806 371
rect 1938 368 1942 371
rect 2074 368 2142 371
rect 2178 368 2265 371
rect 26 358 46 361
rect 118 361 121 368
rect 118 358 222 361
rect 226 358 414 361
rect 482 358 657 361
rect 690 358 806 361
rect 810 358 902 361
rect 1606 361 1609 368
rect 1418 358 1609 361
rect 1710 358 1713 368
rect 1726 362 1729 368
rect 1746 358 1750 361
rect 1794 358 1814 361
rect 1818 358 1870 361
rect 1874 358 1910 361
rect 1934 361 1937 368
rect 1934 358 1974 361
rect 1998 361 2001 368
rect 2262 362 2265 368
rect 2466 368 2654 371
rect 2682 368 2710 371
rect 2730 368 2734 371
rect 3162 368 3270 371
rect 3274 368 3398 371
rect 3450 368 3518 371
rect 3522 368 3606 371
rect 3690 368 3718 371
rect 3818 368 3926 371
rect 4026 368 4062 371
rect 4066 368 4150 371
rect 4170 368 4246 371
rect 4258 368 4270 371
rect 1998 358 2054 361
rect 2130 358 2134 361
rect 2154 358 2158 361
rect 2218 358 2246 361
rect 2302 361 2305 368
rect 2302 358 2326 361
rect 2394 358 2398 361
rect 2446 361 2449 368
rect 2418 358 2449 361
rect 2466 358 2502 361
rect 2506 358 2742 361
rect 2746 358 2750 361
rect 2786 358 2814 361
rect 2822 361 2825 368
rect 4438 362 4441 368
rect 2822 358 2830 361
rect 2850 358 2862 361
rect 3026 358 3030 361
rect 3162 358 3262 361
rect 3298 358 3382 361
rect 3386 358 3406 361
rect 3410 358 3462 361
rect 3538 358 3558 361
rect 3642 358 3718 361
rect 3770 358 3966 361
rect 4018 358 4118 361
rect 4242 358 4246 361
rect 4306 358 4318 361
rect 4502 361 4505 368
rect 4502 358 4566 361
rect 42 348 70 351
rect 178 348 190 351
rect 234 348 249 351
rect 258 348 273 351
rect 314 348 318 351
rect 346 348 470 351
rect 562 348 566 351
rect 654 351 657 358
rect 2350 352 2353 358
rect 578 348 649 351
rect 654 348 745 351
rect 754 348 1174 351
rect 1178 348 1206 351
rect 1230 348 1310 351
rect 1570 348 1590 351
rect 1706 348 1726 351
rect 1730 348 1814 351
rect 1850 348 1854 351
rect 1890 348 1926 351
rect 1930 348 1998 351
rect 2010 348 2302 351
rect 2394 348 2438 351
rect 2442 348 2446 351
rect 2490 348 2494 351
rect 2498 348 2574 351
rect 2594 348 2622 351
rect 2626 348 2662 351
rect 2690 348 2694 351
rect 2706 348 2822 351
rect 2826 348 2830 351
rect 2854 348 2878 351
rect 2914 348 3094 351
rect 3142 351 3145 358
rect 3974 352 3977 358
rect 3142 348 3150 351
rect 3170 348 3174 351
rect 3242 348 3446 351
rect 3450 348 3486 351
rect 3522 348 3630 351
rect 3650 348 3654 351
rect 3722 348 3726 351
rect 3738 348 3774 351
rect 3898 348 3953 351
rect 3994 348 3998 351
rect 4050 348 4150 351
rect 4226 348 4230 351
rect 4250 348 4254 351
rect 4258 348 4270 351
rect 4282 348 4286 351
rect 4314 348 4350 351
rect 4386 348 4406 351
rect 4410 348 4446 351
rect 4498 348 4526 351
rect 4530 348 4550 351
rect 4570 348 4582 351
rect 106 338 126 341
rect 202 338 238 341
rect 246 341 249 348
rect 270 342 273 348
rect 646 342 649 348
rect 742 342 745 348
rect 1230 342 1233 348
rect 1438 342 1441 348
rect 246 338 262 341
rect 314 338 350 341
rect 410 338 430 341
rect 762 338 766 341
rect 770 338 854 341
rect 1138 338 1230 341
rect 1562 338 1574 341
rect 1646 341 1649 348
rect 1578 338 1649 341
rect 1730 338 1734 341
rect 1810 338 1822 341
rect 1842 338 1846 341
rect 1882 338 1926 341
rect 1930 338 1942 341
rect 1962 338 2014 341
rect 2082 338 2102 341
rect 2350 341 2353 348
rect 2462 342 2465 348
rect 2106 338 2353 341
rect 2394 338 2417 341
rect 2470 341 2473 348
rect 2854 342 2857 348
rect 2470 338 2478 341
rect 2538 338 2630 341
rect 2682 338 2694 341
rect 2738 338 2742 341
rect 2770 338 2798 341
rect 2818 338 2822 341
rect 2890 338 2934 341
rect 2978 338 2982 341
rect 3150 341 3153 348
rect 2994 338 3222 341
rect 3226 338 3246 341
rect 3282 338 3286 341
rect 3694 341 3697 348
rect 3950 342 3953 348
rect 3306 338 3697 341
rect 3762 338 3838 341
rect 3954 338 3974 341
rect 3982 341 3985 348
rect 3982 338 3990 341
rect 4022 341 4025 348
rect 4022 338 4046 341
rect 4058 338 4062 341
rect 4106 338 4142 341
rect 4194 338 4534 341
rect 26 328 174 331
rect 238 331 241 338
rect 238 328 382 331
rect 386 328 438 331
rect 474 328 590 331
rect 618 328 790 331
rect 1470 331 1473 338
rect 2414 332 2417 338
rect 1470 328 1502 331
rect 1506 328 1577 331
rect 1586 328 1638 331
rect 1642 328 1662 331
rect 1682 328 1846 331
rect 1858 328 1878 331
rect 1922 328 1982 331
rect 2010 328 2182 331
rect 2186 328 2214 331
rect 2218 328 2230 331
rect 2258 328 2369 331
rect 2638 331 2641 338
rect 2490 328 2641 331
rect 2726 331 2729 338
rect 2726 328 3022 331
rect 3042 328 3086 331
rect 3090 328 3150 331
rect 3306 328 3358 331
rect 3394 328 3398 331
rect 3426 328 3438 331
rect 3506 328 3550 331
rect 3626 328 3662 331
rect 3674 328 3678 331
rect 3682 328 3710 331
rect 3742 331 3745 338
rect 3918 332 3921 338
rect 4542 332 4545 338
rect 3742 328 3790 331
rect 3794 328 3814 331
rect 3842 328 3854 331
rect 3946 328 3982 331
rect 3994 328 4006 331
rect 4018 328 4070 331
rect 4074 328 4081 331
rect 4098 328 4182 331
rect 4190 328 4214 331
rect 4234 328 4238 331
rect 4250 328 4254 331
rect 4282 328 4286 331
rect 4314 328 4361 331
rect 4394 328 4422 331
rect 4426 328 4478 331
rect 4490 328 4494 331
rect 1574 322 1577 328
rect 2326 322 2329 328
rect 2366 322 2369 328
rect 3406 322 3409 328
rect 4190 322 4193 328
rect 4358 322 4361 328
rect 10 318 30 321
rect 34 318 54 321
rect 58 318 126 321
rect 258 318 406 321
rect 602 318 662 321
rect 666 318 726 321
rect 730 318 870 321
rect 874 318 1014 321
rect 1074 318 1078 321
rect 1274 318 1374 321
rect 1530 318 1553 321
rect 1610 318 1662 321
rect 1698 318 1910 321
rect 1922 318 2126 321
rect 2138 318 2150 321
rect 2170 318 2174 321
rect 2410 318 2446 321
rect 2514 318 2718 321
rect 2730 318 2766 321
rect 2786 318 2790 321
rect 2810 318 2814 321
rect 2842 318 2846 321
rect 3010 318 3073 321
rect 3090 318 3094 321
rect 3138 318 3366 321
rect 3458 318 3462 321
rect 3490 318 3694 321
rect 3738 318 3822 321
rect 3858 318 3910 321
rect 3994 318 4110 321
rect 4202 318 4286 321
rect 1390 312 1393 318
rect 170 308 214 311
rect 218 308 326 311
rect 546 308 566 311
rect 570 308 702 311
rect 1426 308 1542 311
rect 1550 311 1553 318
rect 1550 308 1734 311
rect 1762 308 1870 311
rect 1874 308 1950 311
rect 2050 308 2102 311
rect 2162 308 2254 311
rect 2266 308 2318 311
rect 2322 308 2374 311
rect 2610 308 2614 311
rect 2634 308 2678 311
rect 2698 308 2710 311
rect 2818 308 2966 311
rect 3070 311 3073 318
rect 3070 308 3110 311
rect 3178 308 3254 311
rect 3266 308 3398 311
rect 3570 308 3590 311
rect 3618 308 3710 311
rect 3818 308 3910 311
rect 3914 308 3998 311
rect 4026 308 4070 311
rect 4202 308 4222 311
rect 4250 308 4374 311
rect 4378 308 4414 311
rect 4450 308 4558 311
rect 1000 303 1002 307
rect 1006 303 1009 307
rect 1014 303 1016 307
rect 2024 303 2026 307
rect 2030 303 2033 307
rect 2038 303 2040 307
rect 3048 303 3050 307
rect 3054 303 3057 307
rect 3062 303 3064 307
rect 4080 303 4082 307
rect 4086 303 4089 307
rect 4094 303 4096 307
rect 210 298 302 301
rect 314 298 382 301
rect 410 298 486 301
rect 490 298 646 301
rect 650 298 678 301
rect 682 298 702 301
rect 842 298 958 301
rect 1138 298 1550 301
rect 1554 298 1598 301
rect 1650 298 1654 301
rect 1754 298 2014 301
rect 2058 298 2086 301
rect 2146 298 2222 301
rect 2266 298 2358 301
rect 2610 298 2710 301
rect 3138 298 3190 301
rect 3210 298 3246 301
rect 3298 298 3302 301
rect 3514 298 3566 301
rect 3578 298 3694 301
rect 3754 298 3878 301
rect 3882 298 4030 301
rect 4042 298 4070 301
rect 4130 298 4342 301
rect 4354 298 4414 301
rect 4450 298 4470 301
rect 4474 298 4518 301
rect 298 288 390 291
rect 458 288 502 291
rect 754 288 846 291
rect 874 288 1062 291
rect 1170 288 1262 291
rect 1482 288 1510 291
rect 1514 288 1694 291
rect 1746 288 1766 291
rect 1826 288 2006 291
rect 2114 288 2142 291
rect 2154 288 2294 291
rect 2298 288 2305 291
rect 2330 288 2390 291
rect 2458 288 2494 291
rect 2594 288 2662 291
rect 2766 288 2774 291
rect 2778 288 3102 291
rect 3106 288 3414 291
rect 3442 288 3510 291
rect 3554 288 3614 291
rect 3618 288 3625 291
rect 3834 288 3862 291
rect 3866 288 3894 291
rect 3898 288 3950 291
rect 3970 288 4038 291
rect 4054 288 4102 291
rect 4286 288 4294 291
rect 4298 288 4318 291
rect 4322 288 4350 291
rect 4362 288 4478 291
rect 218 278 278 281
rect 282 278 286 281
rect 290 278 318 281
rect 322 278 374 281
rect 498 278 526 281
rect 582 281 585 288
rect 546 278 585 281
rect 594 278 622 281
rect 858 278 1017 281
rect 1034 278 1038 281
rect 1106 278 1326 281
rect 1330 278 1358 281
rect 1722 278 1782 281
rect 1914 278 2286 281
rect 2298 278 2342 281
rect 2362 278 2390 281
rect 2414 281 2417 288
rect 2414 278 2486 281
rect 2498 278 2534 281
rect 2618 278 2630 281
rect 2754 278 2758 281
rect 2770 278 2774 281
rect 2938 278 2982 281
rect 2986 278 3038 281
rect 3042 278 3078 281
rect 3386 278 3390 281
rect 3450 278 3454 281
rect 3474 278 3494 281
rect 3526 281 3529 288
rect 3506 278 3529 281
rect 3542 282 3545 288
rect 4054 282 4057 288
rect 3554 278 3598 281
rect 3602 278 3646 281
rect 3650 278 3654 281
rect 3666 278 3670 281
rect 3706 278 3718 281
rect 3946 278 3958 281
rect 3970 278 3974 281
rect 4110 281 4113 288
rect 4206 282 4209 288
rect 4486 282 4489 288
rect 4110 278 4182 281
rect 4218 278 4222 281
rect 4518 281 4521 288
rect 4514 278 4521 281
rect 158 271 161 278
rect 122 268 161 271
rect 210 268 294 271
rect 298 268 310 271
rect 478 271 481 278
rect 418 268 630 271
rect 818 268 910 271
rect 914 268 934 271
rect 938 268 966 271
rect 1014 271 1017 278
rect 1014 268 1062 271
rect 1298 268 1310 271
rect 1314 268 1390 271
rect 1394 268 1494 271
rect 1582 271 1585 278
rect 1498 268 1585 271
rect 1670 272 1673 278
rect 1674 268 1742 271
rect 1834 268 1838 271
rect 1850 268 1918 271
rect 1938 268 1942 271
rect 1962 268 2022 271
rect 2026 268 2070 271
rect 2138 268 2166 271
rect 2170 268 2190 271
rect 2194 268 2217 271
rect 2234 268 2262 271
rect 2266 268 2414 271
rect 2538 268 2590 271
rect 2602 268 2638 271
rect 2698 268 2702 271
rect 2746 268 2782 271
rect 2866 268 2870 271
rect 2874 268 2894 271
rect 2898 268 2942 271
rect 2946 268 2958 271
rect 3034 268 3086 271
rect 3122 268 3150 271
rect 3154 268 3190 271
rect 3194 268 3222 271
rect 3238 271 3241 278
rect 3742 272 3745 278
rect 3238 268 3350 271
rect 3354 268 3374 271
rect 3410 268 3422 271
rect 3442 268 3454 271
rect 3458 268 3502 271
rect 3506 268 3678 271
rect 3682 268 3686 271
rect 3818 268 3830 271
rect 3850 268 3862 271
rect 3898 268 4110 271
rect 4114 268 4150 271
rect 4154 268 4502 271
rect 130 258 158 261
rect 266 258 270 261
rect 306 258 350 261
rect 410 258 430 261
rect 458 258 478 261
rect 602 258 606 261
rect 618 258 646 261
rect 706 258 782 261
rect 802 258 886 261
rect 890 258 918 261
rect 922 258 974 261
rect 1018 258 1030 261
rect 1050 258 1078 261
rect 1090 258 1110 261
rect 1134 261 1137 268
rect 1166 261 1169 268
rect 2214 262 2217 268
rect 1134 258 1169 261
rect 1234 258 1278 261
rect 1282 258 1342 261
rect 1610 258 1614 261
rect 1730 258 1758 261
rect 1834 258 1894 261
rect 1914 258 1998 261
rect 2002 258 2038 261
rect 2098 258 2110 261
rect 2114 258 2158 261
rect 2162 258 2166 261
rect 2282 258 2294 261
rect 2330 258 2342 261
rect 2386 258 2406 261
rect 2426 258 2446 261
rect 2454 261 2457 268
rect 2450 258 2457 261
rect 2474 258 2598 261
rect 2606 258 2614 261
rect 2686 261 2689 268
rect 3710 262 3713 268
rect 2674 258 2689 261
rect 2802 258 2838 261
rect 2842 258 2870 261
rect 2890 258 2934 261
rect 3194 258 3198 261
rect 3210 258 3222 261
rect 3226 258 3257 261
rect 3346 258 3350 261
rect 3354 258 3390 261
rect 3394 258 3590 261
rect 3594 258 3678 261
rect 3722 258 3782 261
rect 3826 258 3926 261
rect 3938 258 3942 261
rect 3954 258 3998 261
rect 4002 258 4014 261
rect 4042 258 4086 261
rect 4106 258 4134 261
rect 4218 258 4222 261
rect 4226 258 4270 261
rect 4314 258 4318 261
rect 4354 258 4382 261
rect 4410 258 4422 261
rect 246 252 249 258
rect -26 251 -22 252
rect -26 248 6 251
rect 186 248 190 251
rect 202 248 246 251
rect 314 248 358 251
rect 378 248 494 251
rect 550 251 553 258
rect 550 248 630 251
rect 634 248 726 251
rect 834 248 846 251
rect 926 248 934 251
rect 938 248 950 251
rect 970 248 1038 251
rect 1042 248 1102 251
rect 1782 251 1785 258
rect 1442 248 1785 251
rect 1946 248 1958 251
rect 2086 251 2089 258
rect 1994 248 2174 251
rect 2194 248 2198 251
rect 2234 248 2238 251
rect 2354 248 2390 251
rect 2442 248 2446 251
rect 2506 248 2510 251
rect 2546 248 2566 251
rect 2602 248 2622 251
rect 2662 251 2665 258
rect 3254 252 3257 258
rect 4390 252 4393 258
rect 2662 248 2718 251
rect 2746 248 2750 251
rect 2754 248 2822 251
rect 2878 248 2886 251
rect 2890 248 2902 251
rect 2930 248 2934 251
rect 2970 248 2998 251
rect 3082 248 3222 251
rect 3266 248 3854 251
rect 3858 248 4078 251
rect 4094 248 4166 251
rect 4298 248 4358 251
rect 130 238 238 241
rect 250 238 278 241
rect 282 238 294 241
rect 298 238 342 241
rect 354 238 358 241
rect 362 238 558 241
rect 798 241 801 248
rect 798 238 814 241
rect 894 241 897 248
rect 2950 242 2953 248
rect 894 238 1118 241
rect 1810 238 1982 241
rect 2114 238 2238 241
rect 2258 238 2526 241
rect 2530 238 2638 241
rect 2642 238 2670 241
rect 2690 238 2710 241
rect 2842 238 2910 241
rect 2970 238 3014 241
rect 3314 238 3318 241
rect 3338 238 3414 241
rect 3418 238 3470 241
rect 3474 238 3558 241
rect 3562 238 3590 241
rect 3618 238 3758 241
rect 3786 238 3838 241
rect 3842 238 3870 241
rect 3946 238 3974 241
rect 4058 238 4062 241
rect 4094 241 4097 248
rect 4082 238 4097 241
rect 4162 238 4238 241
rect 4258 238 4286 241
rect 4290 238 4454 241
rect 206 228 214 231
rect 218 228 230 231
rect 338 228 774 231
rect 778 228 1230 231
rect 1458 228 2126 231
rect 2266 228 2310 231
rect 2314 228 2318 231
rect 2322 228 2334 231
rect 2338 228 2510 231
rect 2522 228 2582 231
rect 2626 228 2942 231
rect 2946 228 2982 231
rect 2986 228 3054 231
rect 3058 228 3118 231
rect 3346 228 3374 231
rect 3378 228 3574 231
rect 3690 228 3742 231
rect 3774 228 4126 231
rect 4154 228 4166 231
rect 4186 228 4414 231
rect 154 218 318 221
rect 322 218 542 221
rect 882 218 982 221
rect 1058 218 1398 221
rect 1402 218 1430 221
rect 1858 218 2649 221
rect 2666 218 2798 221
rect 2938 218 3078 221
rect 3090 218 3302 221
rect 3482 218 3486 221
rect 3506 218 3510 221
rect 3518 218 3662 221
rect 3774 221 3777 228
rect 3722 218 3777 221
rect 3786 218 3862 221
rect 3906 218 3918 221
rect 3962 218 4022 221
rect 4026 218 4078 221
rect 4098 218 4342 221
rect 4410 218 4494 221
rect 314 208 422 211
rect 666 208 1094 211
rect 1098 208 1166 211
rect 1890 208 1894 211
rect 1930 208 2206 211
rect 2210 208 2246 211
rect 2282 208 2358 211
rect 2442 208 2494 211
rect 2646 211 2649 218
rect 3518 212 3521 218
rect 2646 208 3518 211
rect 3682 208 3774 211
rect 3786 208 3910 211
rect 3986 208 4038 211
rect 4042 208 4054 211
rect 4066 208 4214 211
rect 4258 208 4518 211
rect 496 203 498 207
rect 502 203 505 207
rect 510 203 512 207
rect 1520 203 1522 207
rect 1526 203 1529 207
rect 1534 203 1536 207
rect 74 198 222 201
rect 362 198 462 201
rect 538 198 614 201
rect 722 198 1318 201
rect 1938 198 1974 201
rect 1978 198 2286 201
rect 2358 201 2361 208
rect 2544 203 2546 207
rect 2550 203 2553 207
rect 2558 203 2560 207
rect 3568 203 3570 207
rect 3574 203 3577 207
rect 3582 203 3584 207
rect 2358 198 2462 201
rect 2642 198 2790 201
rect 2802 198 2862 201
rect 3026 198 3062 201
rect 3066 198 3126 201
rect 3250 198 3438 201
rect 3474 198 3486 201
rect 3498 198 3558 201
rect 3626 198 3774 201
rect 3802 198 3854 201
rect 3858 198 4086 201
rect 4226 198 4246 201
rect 4266 198 4486 201
rect 4490 198 4542 201
rect 26 188 94 191
rect 98 188 150 191
rect 250 188 366 191
rect 462 191 465 198
rect 462 188 678 191
rect 682 188 702 191
rect 1242 188 1454 191
rect 1458 188 1526 191
rect 1650 188 1870 191
rect 1922 188 2262 191
rect 2298 188 2398 191
rect 2462 191 2465 198
rect 2462 188 2590 191
rect 2594 188 2630 191
rect 2674 188 2862 191
rect 2874 188 2886 191
rect 2978 188 2982 191
rect 2986 188 3078 191
rect 3154 188 3670 191
rect 3674 188 3734 191
rect 3762 188 3782 191
rect 3890 188 4054 191
rect 4058 188 4118 191
rect 4146 188 4446 191
rect 2358 182 2361 188
rect 210 178 238 181
rect 266 178 326 181
rect 394 178 558 181
rect 562 178 569 181
rect 706 178 758 181
rect 962 178 1030 181
rect 1042 178 1046 181
rect 1074 178 1142 181
rect 1146 178 1174 181
rect 1290 178 2046 181
rect 2050 178 2102 181
rect 2130 178 2166 181
rect 2194 178 2350 181
rect 2402 178 2478 181
rect 2482 178 2662 181
rect 2858 178 3550 181
rect 3554 178 3630 181
rect 3658 178 3918 181
rect 3938 178 3958 181
rect 4050 178 4305 181
rect 4322 178 4382 181
rect 226 168 294 171
rect 514 168 574 171
rect 866 168 942 171
rect 946 168 1078 171
rect 1106 168 1326 171
rect 1330 168 1910 171
rect 2094 168 2366 171
rect 2370 168 2574 171
rect 2578 168 2734 171
rect 2746 168 2758 171
rect 2770 168 2878 171
rect 2882 168 2926 171
rect 2954 168 2958 171
rect 2978 168 2982 171
rect 3130 168 3158 171
rect 3234 168 3238 171
rect 3290 168 3318 171
rect 3322 168 3334 171
rect 3362 168 3806 171
rect 3818 168 3990 171
rect 3994 168 4006 171
rect 4066 168 4142 171
rect 4154 168 4230 171
rect 4234 168 4294 171
rect 4302 171 4305 178
rect 4302 168 4369 171
rect 242 158 270 161
rect 274 158 350 161
rect 390 161 393 168
rect 390 158 422 161
rect 582 161 585 168
rect 2094 162 2097 168
rect 3110 162 3113 168
rect 4366 162 4369 168
rect 434 158 622 161
rect 634 158 902 161
rect 930 158 934 161
rect 1002 158 1182 161
rect 1202 158 1214 161
rect 1794 158 1846 161
rect 1850 158 1854 161
rect 1946 158 2094 161
rect 2138 158 2150 161
rect 2206 158 2214 161
rect 2218 158 2270 161
rect 2274 158 2350 161
rect 2354 158 2414 161
rect 2418 158 2686 161
rect 2698 158 2790 161
rect 2794 158 2918 161
rect 2922 158 2990 161
rect 3026 158 3030 161
rect 3042 158 3094 161
rect 3194 158 3238 161
rect 3258 158 3262 161
rect 3270 158 3278 161
rect 3298 158 3318 161
rect 3338 158 3366 161
rect 3370 158 3454 161
rect 3458 158 3646 161
rect 3682 158 3686 161
rect 3698 158 3702 161
rect 3714 158 3782 161
rect 3790 158 3798 161
rect 3802 158 3846 161
rect 3850 158 3934 161
rect 3946 158 3950 161
rect 4042 158 4094 161
rect 4098 158 4110 161
rect 4162 158 4174 161
rect 4250 158 4302 161
rect 4306 158 4318 161
rect 4510 161 4513 168
rect 4474 158 4513 161
rect 166 151 169 158
rect 222 151 225 158
rect 950 152 953 158
rect 90 148 137 151
rect 166 148 225 151
rect 234 148 254 151
rect 346 148 366 151
rect 562 148 606 151
rect 610 148 646 151
rect 858 148 950 151
rect 954 148 1086 151
rect 1818 148 1878 151
rect 1882 148 1998 151
rect 2002 148 2062 151
rect 2066 148 2118 151
rect 2122 148 2166 151
rect 2170 148 2182 151
rect 2186 148 2198 151
rect 2242 148 2310 151
rect 2378 148 2382 151
rect 2402 148 2470 151
rect 2474 148 2542 151
rect 2546 148 2553 151
rect 2610 148 2614 151
rect 2690 148 2702 151
rect 2730 148 2742 151
rect 2754 148 2758 151
rect 2770 148 2774 151
rect 2794 148 2846 151
rect 2850 148 2862 151
rect 2866 148 2942 151
rect 2946 148 3134 151
rect 3138 148 3166 151
rect 3170 148 3174 151
rect 3178 148 3198 151
rect 3202 148 3350 151
rect 3354 148 3478 151
rect 3482 148 3510 151
rect 3522 148 3526 151
rect 3538 148 3606 151
rect 3610 148 3702 151
rect 3778 148 3790 151
rect 3794 148 3822 151
rect 3838 148 3854 151
rect 3874 148 3894 151
rect 3898 148 4030 151
rect 4034 148 4134 151
rect 4154 148 4158 151
rect 4190 151 4193 158
rect 4170 148 4193 151
rect 4198 152 4201 158
rect 4218 148 4230 151
rect 4370 148 4374 151
rect 4402 148 4438 151
rect 4454 151 4457 158
rect 4542 152 4545 158
rect 4442 148 4457 151
rect 4506 148 4510 151
rect 134 142 137 148
rect 326 141 329 148
rect 406 141 409 148
rect 326 138 409 141
rect 490 138 526 141
rect 578 138 598 141
rect 618 138 638 141
rect 706 138 718 141
rect 882 138 1102 141
rect 1178 138 1206 141
rect 1562 138 1630 141
rect 1662 141 1665 148
rect 1678 141 1681 148
rect 1634 138 1681 141
rect 1694 142 1697 148
rect 3838 142 3841 148
rect 4206 142 4209 148
rect 4342 142 4345 148
rect 1714 138 1897 141
rect 1986 138 2078 141
rect 2178 138 2302 141
rect 2310 138 2318 141
rect 2322 138 2366 141
rect 2386 138 2414 141
rect 2426 138 2430 141
rect 2466 138 2710 141
rect 2714 138 2774 141
rect 2802 138 2806 141
rect 2946 138 2950 141
rect 3002 138 3014 141
rect 3042 138 3126 141
rect 3186 138 3214 141
rect 3226 138 3230 141
rect 3234 138 3422 141
rect 3426 138 3438 141
rect 3466 138 3534 141
rect 3546 138 3566 141
rect 3578 138 3590 141
rect 3658 138 3718 141
rect 3738 138 3742 141
rect 3762 138 3830 141
rect 3858 138 3886 141
rect 3922 138 3934 141
rect 3946 138 3966 141
rect 3978 138 3982 141
rect 3994 138 4022 141
rect 4042 138 4118 141
rect 4122 138 4145 141
rect 4154 138 4158 141
rect 4274 138 4294 141
rect 4418 138 4470 141
rect 4538 138 4542 141
rect 1774 132 1777 138
rect 1894 132 1897 138
rect 554 128 622 131
rect 714 128 878 131
rect 1114 128 1158 131
rect 1162 128 1270 131
rect 1978 128 2078 131
rect 2154 128 2222 131
rect 2298 128 2326 131
rect 2370 128 2374 131
rect 2386 128 2438 131
rect 2442 128 2470 131
rect 2594 128 2598 131
rect 2618 128 2633 131
rect 2642 128 2646 131
rect 2722 128 2854 131
rect 2946 128 3534 131
rect 3546 128 3550 131
rect 3562 128 3598 131
rect 3714 128 3766 131
rect 3778 128 3886 131
rect 3910 131 3913 138
rect 3906 128 3913 131
rect 3930 128 3942 131
rect 3946 128 3950 131
rect 3986 128 4014 131
rect 4018 128 4054 131
rect 4114 128 4118 131
rect 4142 131 4145 138
rect 4358 132 4361 138
rect 4142 128 4166 131
rect 4178 128 4334 131
rect 4346 128 4350 131
rect 4362 128 4406 131
rect 4434 128 4438 131
rect 4442 128 4526 131
rect 2630 122 2633 128
rect 3606 122 3609 128
rect 18 118 22 121
rect 26 118 54 121
rect 602 118 790 121
rect 846 118 1014 121
rect 1074 118 1134 121
rect 1402 118 1406 121
rect 1522 118 1798 121
rect 1882 118 1982 121
rect 2002 118 2150 121
rect 2210 118 2486 121
rect 2490 118 2518 121
rect 2522 118 2558 121
rect 2602 118 2606 121
rect 2642 118 3270 121
rect 3274 118 3278 121
rect 3298 118 3366 121
rect 3378 118 3462 121
rect 3474 118 3590 121
rect 3698 118 4318 121
rect 4322 118 4422 121
rect 4530 118 4598 121
rect 846 112 849 118
rect 778 108 846 111
rect 898 108 974 111
rect 1202 108 1390 111
rect 1394 108 1462 111
rect 1570 108 1590 111
rect 1954 108 2006 111
rect 2082 108 2222 111
rect 2226 108 2278 111
rect 2378 108 2406 111
rect 2426 108 2454 111
rect 2458 108 2494 111
rect 2578 108 2774 111
rect 2794 108 2806 111
rect 2810 108 2830 111
rect 2922 108 3038 111
rect 3138 108 3174 111
rect 3226 108 3262 111
rect 3274 108 3310 111
rect 3314 108 3366 111
rect 3386 108 3438 111
rect 3450 108 3518 111
rect 3530 108 3558 111
rect 3578 108 3750 111
rect 3778 108 3782 111
rect 3786 108 3798 111
rect 3810 108 3870 111
rect 3890 108 3902 111
rect 3914 108 4070 111
rect 4106 108 4118 111
rect 4130 108 4190 111
rect 4194 108 4230 111
rect 4242 108 4270 111
rect 4314 108 4326 111
rect 4354 108 4478 111
rect 1000 103 1002 107
rect 1006 103 1009 107
rect 1014 103 1016 107
rect 2024 103 2026 107
rect 2030 103 2033 107
rect 2038 103 2040 107
rect 3048 103 3050 107
rect 3054 103 3057 107
rect 3062 103 3064 107
rect 4080 103 4082 107
rect 4086 103 4089 107
rect 4094 103 4096 107
rect 738 98 838 101
rect 842 98 918 101
rect 2050 98 2134 101
rect 2138 98 2198 101
rect 2274 98 2638 101
rect 2698 98 2726 101
rect 2738 98 2814 101
rect 2882 98 2910 101
rect 2930 98 2934 101
rect 2962 98 2974 101
rect 3162 98 3230 101
rect 3234 98 3270 101
rect 3282 98 3430 101
rect 3450 98 3582 101
rect 3594 98 3662 101
rect 3674 98 4006 101
rect 4050 98 4070 101
rect 4114 98 4302 101
rect 4338 98 4430 101
rect 226 88 230 91
rect 362 88 446 91
rect 450 88 686 91
rect 698 88 782 91
rect 938 88 958 91
rect 962 88 1718 91
rect 1890 88 2062 91
rect 2066 88 2158 91
rect 2162 88 2214 91
rect 2218 88 2294 91
rect 2298 88 2422 91
rect 2434 88 2462 91
rect 2534 88 2630 91
rect 2634 88 2662 91
rect 2666 88 3086 91
rect 3090 88 3278 91
rect 3306 88 3398 91
rect 3402 88 3598 91
rect 3602 88 3846 91
rect 3882 88 3998 91
rect 4074 88 4102 91
rect 4162 88 4182 91
rect 4210 88 4270 91
rect 4282 88 4286 91
rect 4314 88 4454 91
rect 4458 88 4478 91
rect 98 78 262 81
rect 410 78 574 81
rect 578 78 654 81
rect 658 78 774 81
rect 810 78 870 81
rect 874 78 934 81
rect 938 78 1110 81
rect 1922 78 1982 81
rect 1986 78 1998 81
rect 2122 78 2182 81
rect 2194 78 2281 81
rect 2290 78 2350 81
rect 2354 78 2358 81
rect 2430 81 2433 88
rect 2394 78 2433 81
rect 2470 81 2473 88
rect 2534 82 2537 88
rect 4190 82 4193 88
rect 2470 78 2502 81
rect 2506 78 2534 81
rect 2626 78 2630 81
rect 2650 78 2670 81
rect 2682 78 2766 81
rect 2770 78 3070 81
rect 3082 78 3102 81
rect 3106 78 3142 81
rect 3162 78 3166 81
rect 3170 78 3198 81
rect 3210 78 3254 81
rect 3266 78 3310 81
rect 3330 78 3342 81
rect 3346 78 3390 81
rect 3394 78 3422 81
rect 3426 78 3430 81
rect 3442 78 3622 81
rect 3706 78 3718 81
rect 3746 78 3750 81
rect 3770 78 3774 81
rect 3794 78 3798 81
rect 3866 78 3878 81
rect 3914 78 3918 81
rect 3930 78 3934 81
rect 3998 78 4134 81
rect 4250 78 4262 81
rect 4274 78 4294 81
rect 4310 81 4313 88
rect 4534 82 4537 88
rect 4310 78 4334 81
rect 4346 78 4374 81
rect 4378 78 4430 81
rect 4450 78 4470 81
rect 186 68 278 71
rect 946 68 958 71
rect 1818 68 1830 71
rect 1874 68 2270 71
rect 2278 71 2281 78
rect 3838 72 3841 78
rect 3894 72 3897 78
rect 2278 68 2366 71
rect 2402 68 2406 71
rect 2426 68 2510 71
rect 2522 68 2526 71
rect 2570 68 2574 71
rect 2594 68 2790 71
rect 2818 68 2822 71
rect 2842 68 2849 71
rect 2858 68 2878 71
rect 2962 68 2990 71
rect 3002 68 3286 71
rect 3290 68 3366 71
rect 3370 68 3438 71
rect 3442 68 3462 71
rect 3482 68 3502 71
rect 3530 68 3550 71
rect 3602 68 3630 71
rect 3642 68 3670 71
rect 3722 68 3822 71
rect 3910 68 3918 71
rect 3922 68 3950 71
rect 3958 71 3961 78
rect 3974 71 3977 78
rect 3958 68 3977 71
rect 3998 72 4001 78
rect 4034 68 4038 71
rect 4050 68 4054 71
rect 4130 68 4142 71
rect 4178 68 4182 71
rect 4258 68 4262 71
rect 4274 68 4318 71
rect 4394 68 4398 71
rect 4402 68 4438 71
rect 4530 68 4550 71
rect 118 61 121 68
rect 118 58 198 61
rect 354 59 398 61
rect 402 59 486 61
rect 354 58 486 59
rect 578 58 582 61
rect 622 58 630 61
rect 634 59 678 61
rect 682 59 742 61
rect 634 58 742 59
rect 794 58 822 61
rect 826 59 870 61
rect 874 59 894 61
rect 826 58 894 59
rect 1198 61 1201 68
rect 1198 58 1294 61
rect 1614 61 1617 68
rect 3862 62 3865 68
rect 1514 58 1617 61
rect 1798 58 1806 61
rect 1826 58 1846 61
rect 1914 58 2070 61
rect 2090 58 2118 61
rect 2138 58 2150 61
rect 2202 58 2238 61
rect 2242 58 2310 61
rect 2314 58 2326 61
rect 2330 58 2750 61
rect 2754 58 2782 61
rect 2786 58 2934 61
rect 2986 58 3009 61
rect 3026 58 3030 61
rect 3042 58 3046 61
rect 3074 58 3342 61
rect 3346 58 3382 61
rect 3434 58 3454 61
rect 3458 58 3478 61
rect 3490 58 3494 61
rect 3498 58 3526 61
rect 3530 58 3574 61
rect 3706 58 3726 61
rect 3802 58 3806 61
rect 3906 58 3910 61
rect 3922 58 3926 61
rect 3946 58 3966 61
rect 4026 58 4030 61
rect 4130 58 4134 61
rect 4162 58 4342 61
rect 4366 61 4369 68
rect 4366 58 4422 61
rect 4426 58 4470 61
rect 4482 58 4566 61
rect 1046 52 1049 58
rect 1798 52 1801 58
rect 3006 52 3009 58
rect -26 51 -22 52
rect -26 48 6 51
rect 2010 48 2014 51
rect 2018 48 2062 51
rect 2074 48 2142 51
rect 2146 48 2190 51
rect 2242 48 2246 51
rect 2258 48 2286 51
rect 2458 48 2702 51
rect 2706 48 2870 51
rect 2914 48 2958 51
rect 2978 48 2982 51
rect 3018 48 3022 51
rect 3046 48 3054 51
rect 3058 48 3110 51
rect 3122 48 3126 51
rect 3154 48 3174 51
rect 3178 48 3214 51
rect 3242 48 3246 51
rect 3258 48 3270 51
rect 3274 48 3278 51
rect 3290 48 3294 51
rect 3306 48 3310 51
rect 3410 48 3598 51
rect 3610 48 3614 51
rect 3618 48 3694 51
rect 3782 51 3785 58
rect 3854 52 3857 58
rect 3762 48 3785 51
rect 3810 48 3814 51
rect 3834 48 3846 51
rect 3938 48 3942 51
rect 3970 48 3974 51
rect 3994 48 4070 51
rect 4186 48 4190 51
rect 4226 48 4230 51
rect 4282 48 4342 51
rect 4346 48 4382 51
rect 4386 48 4414 51
rect 4418 48 4494 51
rect 4506 48 4574 51
rect 2042 38 2102 41
rect 2334 41 2337 48
rect 2334 38 2486 41
rect 2490 38 3414 41
rect 3418 38 3654 41
rect 3658 38 3790 41
rect 3798 41 3801 48
rect 3798 38 4014 41
rect 4050 38 4198 41
rect 4306 38 4374 41
rect 4378 38 4406 41
rect 4554 38 4574 41
rect 3110 28 3118 31
rect 3122 28 3318 31
rect 3334 28 3342 31
rect 3346 28 3774 31
rect 3850 28 3886 31
rect 3954 28 4046 31
rect 4058 28 4089 31
rect 4142 28 4150 31
rect 4154 28 4366 31
rect 4386 28 4494 31
rect 3082 18 3726 21
rect 3730 18 3910 21
rect 3954 18 3969 21
rect 4050 18 4078 21
rect 4086 21 4089 28
rect 4086 18 4166 21
rect 4170 18 4222 21
rect 786 8 790 11
rect 1034 8 1038 11
rect 3682 8 3958 11
rect 3966 11 3969 18
rect 3966 8 4262 11
rect 496 3 498 7
rect 502 3 505 7
rect 510 3 512 7
rect 1520 3 1522 7
rect 1526 3 1529 7
rect 1534 3 1536 7
rect 2544 3 2546 7
rect 2550 3 2553 7
rect 2558 3 2560 7
rect 3568 3 3570 7
rect 3574 3 3577 7
rect 3582 3 3584 7
<< m4contact >>
rect 498 4403 502 4407
rect 506 4403 509 4407
rect 509 4403 510 4407
rect 1522 4403 1526 4407
rect 1530 4403 1533 4407
rect 1533 4403 1534 4407
rect 2546 4403 2550 4407
rect 2554 4403 2557 4407
rect 2557 4403 2558 4407
rect 3570 4403 3574 4407
rect 3578 4403 3581 4407
rect 3581 4403 3582 4407
rect 3758 4398 3762 4402
rect 3822 4398 3826 4402
rect 4014 4398 4018 4402
rect 4054 4398 4058 4402
rect 4158 4398 4162 4402
rect 4374 4398 4378 4402
rect 1998 4388 2002 4392
rect 3942 4388 3946 4392
rect 3998 4388 4002 4392
rect 4022 4388 4026 4392
rect 4366 4388 4370 4392
rect 3494 4368 3498 4372
rect 3766 4368 3770 4372
rect 3918 4368 3922 4372
rect 4190 4368 4194 4372
rect 790 4358 794 4362
rect 1758 4358 1762 4362
rect 2678 4358 2682 4362
rect 3422 4358 3426 4362
rect 4062 4358 4066 4362
rect 4142 4358 4146 4362
rect 4214 4358 4218 4362
rect 4438 4358 4442 4362
rect 2526 4348 2530 4352
rect 3070 4348 3074 4352
rect 3550 4348 3554 4352
rect 3694 4348 3698 4352
rect 3798 4348 3802 4352
rect 3934 4348 3938 4352
rect 3974 4348 3978 4352
rect 4166 4348 4170 4352
rect 4358 4348 4362 4352
rect 4398 4348 4402 4352
rect 4446 4348 4450 4352
rect 4494 4348 4498 4352
rect 4526 4348 4530 4352
rect 4582 4348 4586 4352
rect 2302 4338 2306 4342
rect 3238 4338 3242 4342
rect 3366 4338 3370 4342
rect 3486 4338 3490 4342
rect 3494 4338 3498 4342
rect 3686 4338 3690 4342
rect 3958 4338 3962 4342
rect 4110 4338 4114 4342
rect 4334 4338 4338 4342
rect 4350 4338 4354 4342
rect 4406 4338 4410 4342
rect 4462 4338 4466 4342
rect 4510 4338 4514 4342
rect 614 4328 618 4332
rect 790 4328 794 4332
rect 934 4328 938 4332
rect 2422 4328 2426 4332
rect 2814 4328 2818 4332
rect 3262 4328 3266 4332
rect 3494 4328 3498 4332
rect 3702 4328 3706 4332
rect 4102 4328 4106 4332
rect 4118 4328 4122 4332
rect 4350 4328 4354 4332
rect 4358 4328 4362 4332
rect 4422 4328 4426 4332
rect 4558 4328 4562 4332
rect 678 4318 682 4322
rect 1766 4318 1770 4322
rect 2662 4318 2666 4322
rect 3678 4318 3682 4322
rect 3686 4318 3690 4322
rect 3806 4318 3810 4322
rect 3958 4318 3962 4322
rect 3990 4318 3994 4322
rect 4054 4318 4058 4322
rect 4142 4318 4146 4322
rect 4174 4318 4178 4322
rect 334 4308 338 4312
rect 934 4308 938 4312
rect 3654 4308 3658 4312
rect 3718 4308 3722 4312
rect 4302 4308 4306 4312
rect 4310 4308 4314 4312
rect 4518 4308 4522 4312
rect 4550 4308 4554 4312
rect 1002 4303 1006 4307
rect 1010 4303 1013 4307
rect 1013 4303 1014 4307
rect 2026 4303 2030 4307
rect 2034 4303 2037 4307
rect 2037 4303 2038 4307
rect 3050 4303 3054 4307
rect 3058 4303 3061 4307
rect 3061 4303 3062 4307
rect 4082 4303 4086 4307
rect 4090 4303 4093 4307
rect 4093 4303 4094 4307
rect 350 4298 354 4302
rect 3278 4298 3282 4302
rect 3670 4298 3674 4302
rect 3742 4298 3746 4302
rect 3750 4298 3754 4302
rect 3814 4298 3818 4302
rect 4454 4298 4458 4302
rect 958 4288 962 4292
rect 2078 4288 2082 4292
rect 2270 4288 2274 4292
rect 3494 4288 3498 4292
rect 3902 4288 3906 4292
rect 4102 4288 4106 4292
rect 4574 4288 4578 4292
rect 4430 4278 4434 4282
rect 4454 4278 4458 4282
rect 4534 4278 4538 4282
rect 302 4268 306 4272
rect 534 4268 538 4272
rect 870 4268 874 4272
rect 1558 4268 1562 4272
rect 1814 4268 1818 4272
rect 2110 4268 2114 4272
rect 2286 4268 2290 4272
rect 2334 4268 2338 4272
rect 2534 4268 2538 4272
rect 2846 4268 2850 4272
rect 3990 4268 3994 4272
rect 1102 4258 1106 4262
rect 1206 4258 1210 4262
rect 1358 4258 1362 4262
rect 1366 4258 1370 4262
rect 1486 4258 1490 4262
rect 2006 4258 2010 4262
rect 2166 4258 2170 4262
rect 2406 4258 2410 4262
rect 3734 4258 3738 4262
rect 3750 4258 3754 4262
rect 3766 4258 3770 4262
rect 3782 4258 3786 4262
rect 3790 4258 3794 4262
rect 3814 4258 3818 4262
rect 3862 4258 3866 4262
rect 4006 4258 4010 4262
rect 4302 4258 4306 4262
rect 4350 4258 4354 4262
rect 4478 4258 4482 4262
rect 4566 4258 4570 4262
rect 518 4248 522 4252
rect 534 4248 538 4252
rect 710 4248 714 4252
rect 814 4248 818 4252
rect 942 4248 946 4252
rect 1246 4248 1250 4252
rect 2150 4248 2154 4252
rect 2278 4248 2282 4252
rect 2502 4248 2506 4252
rect 2646 4248 2650 4252
rect 3702 4248 3706 4252
rect 4190 4248 4194 4252
rect 4278 4248 4282 4252
rect 4294 4248 4298 4252
rect 4382 4248 4386 4252
rect 958 4238 962 4242
rect 1462 4238 1466 4242
rect 1982 4238 1986 4242
rect 2478 4238 2482 4242
rect 2662 4238 2666 4242
rect 3422 4238 3426 4242
rect 4134 4238 4138 4242
rect 4350 4238 4354 4242
rect 4478 4238 4482 4242
rect 470 4228 474 4232
rect 3622 4228 3626 4232
rect 3830 4228 3834 4232
rect 3918 4228 3922 4232
rect 4126 4228 4130 4232
rect 4254 4228 4258 4232
rect 4318 4228 4322 4232
rect 270 4218 274 4222
rect 1494 4218 1498 4222
rect 3718 4218 3722 4222
rect 3758 4218 3762 4222
rect 4566 4218 4570 4222
rect 2318 4208 2322 4212
rect 2534 4208 2538 4212
rect 2678 4208 2682 4212
rect 3326 4208 3330 4212
rect 4102 4208 4106 4212
rect 4142 4208 4146 4212
rect 4550 4208 4554 4212
rect 498 4203 502 4207
rect 506 4203 509 4207
rect 509 4203 510 4207
rect 1522 4203 1526 4207
rect 1530 4203 1533 4207
rect 1533 4203 1534 4207
rect 2546 4203 2550 4207
rect 2554 4203 2557 4207
rect 2557 4203 2558 4207
rect 3570 4203 3574 4207
rect 3578 4203 3581 4207
rect 3581 4203 3582 4207
rect 838 4198 842 4202
rect 3966 4198 3970 4202
rect 702 4188 706 4192
rect 1126 4188 1130 4192
rect 2238 4188 2242 4192
rect 2286 4188 2290 4192
rect 2414 4188 2418 4192
rect 2678 4188 2682 4192
rect 2766 4188 2770 4192
rect 3158 4188 3162 4192
rect 4430 4188 4434 4192
rect 1934 4178 1938 4182
rect 2798 4178 2802 4182
rect 4414 4178 4418 4182
rect 1254 4168 1258 4172
rect 2414 4168 2418 4172
rect 2510 4168 2514 4172
rect 2686 4168 2690 4172
rect 3694 4168 3698 4172
rect 4022 4168 4026 4172
rect 4142 4168 4146 4172
rect 4158 4168 4162 4172
rect 4334 4168 4338 4172
rect 4558 4168 4562 4172
rect 382 4158 386 4162
rect 702 4158 706 4162
rect 726 4158 730 4162
rect 1302 4158 1306 4162
rect 1446 4158 1450 4162
rect 1790 4158 1794 4162
rect 2206 4158 2210 4162
rect 2222 4158 2226 4162
rect 2430 4158 2434 4162
rect 2526 4158 2530 4162
rect 3662 4158 3666 4162
rect 4118 4158 4122 4162
rect 630 4148 634 4152
rect 798 4148 802 4152
rect 1406 4148 1410 4152
rect 1694 4148 1698 4152
rect 1766 4148 1770 4152
rect 1846 4148 1850 4152
rect 2254 4148 2258 4152
rect 2334 4148 2338 4152
rect 2342 4148 2346 4152
rect 2726 4148 2730 4152
rect 3982 4148 3986 4152
rect 4062 4148 4066 4152
rect 4590 4148 4594 4152
rect 334 4138 338 4142
rect 542 4138 546 4142
rect 854 4138 858 4142
rect 1046 4138 1050 4142
rect 1918 4138 1922 4142
rect 2814 4138 2818 4142
rect 3430 4138 3434 4142
rect 246 4128 250 4132
rect 990 4128 994 4132
rect 1966 4128 1970 4132
rect 2086 4128 2090 4132
rect 3302 4128 3306 4132
rect 3918 4128 3922 4132
rect 574 4118 578 4122
rect 718 4118 722 4122
rect 2350 4118 2354 4122
rect 2654 4118 2658 4122
rect 2662 4118 2666 4122
rect 4438 4118 4442 4122
rect 4598 4118 4602 4122
rect 1974 4108 1978 4112
rect 2238 4108 2242 4112
rect 2910 4108 2914 4112
rect 3070 4108 3074 4112
rect 3942 4108 3946 4112
rect 4102 4108 4106 4112
rect 4470 4108 4474 4112
rect 1002 4103 1006 4107
rect 1010 4103 1013 4107
rect 1013 4103 1014 4107
rect 2026 4103 2030 4107
rect 2034 4103 2037 4107
rect 2037 4103 2038 4107
rect 3050 4103 3054 4107
rect 3058 4103 3061 4107
rect 3061 4103 3062 4107
rect 4082 4103 4086 4107
rect 4090 4103 4093 4107
rect 4093 4103 4094 4107
rect 2358 4098 2362 4102
rect 2854 4098 2858 4102
rect 3358 4098 3362 4102
rect 3814 4098 3818 4102
rect 4294 4098 4298 4102
rect 4454 4098 4458 4102
rect 470 4088 474 4092
rect 1766 4088 1770 4092
rect 4110 4088 4114 4092
rect 4134 4088 4138 4092
rect 174 4078 178 4082
rect 2110 4078 2114 4082
rect 2446 4078 2450 4082
rect 2470 4078 2474 4082
rect 2638 4078 2642 4082
rect 2654 4078 2658 4082
rect 3038 4078 3042 4082
rect 3262 4078 3266 4082
rect 3662 4078 3666 4082
rect 3910 4078 3914 4082
rect 4118 4078 4122 4082
rect 4470 4078 4474 4082
rect 4534 4078 4538 4082
rect 238 4068 242 4072
rect 334 4068 338 4072
rect 830 4068 834 4072
rect 1838 4068 1842 4072
rect 2590 4068 2594 4072
rect 2622 4068 2626 4072
rect 3430 4068 3434 4072
rect 4134 4068 4138 4072
rect 4142 4068 4146 4072
rect 4230 4068 4234 4072
rect 4326 4068 4330 4072
rect 4358 4068 4362 4072
rect 1494 4058 1498 4062
rect 1502 4058 1506 4062
rect 1782 4058 1786 4062
rect 1918 4058 1922 4062
rect 2334 4058 2338 4062
rect 2710 4058 2714 4062
rect 2830 4058 2834 4062
rect 2894 4058 2898 4062
rect 4486 4058 4490 4062
rect 334 4048 338 4052
rect 486 4048 490 4052
rect 2494 4048 2498 4052
rect 2510 4048 2514 4052
rect 2614 4048 2618 4052
rect 854 4038 858 4042
rect 1102 4038 1106 4042
rect 1926 4038 1930 4042
rect 2006 4038 2010 4042
rect 2302 4038 2306 4042
rect 2390 4038 2394 4042
rect 4366 4048 4370 4052
rect 3998 4038 4002 4042
rect 4046 4038 4050 4042
rect 4350 4038 4354 4042
rect 4374 4038 4378 4042
rect 1846 4028 1850 4032
rect 3734 4028 3738 4032
rect 3982 4028 3986 4032
rect 4558 4028 4562 4032
rect 358 4018 362 4022
rect 1102 4018 1106 4022
rect 1486 4018 1490 4022
rect 2222 4018 2226 4022
rect 2806 4018 2810 4022
rect 3998 4018 4002 4022
rect 246 4008 250 4012
rect 486 4008 490 4012
rect 2446 4008 2450 4012
rect 2702 4008 2706 4012
rect 3030 4008 3034 4012
rect 3622 4008 3626 4012
rect 4062 4008 4066 4012
rect 4166 4008 4170 4012
rect 498 4003 502 4007
rect 506 4003 509 4007
rect 509 4003 510 4007
rect 1522 4003 1526 4007
rect 1530 4003 1533 4007
rect 1533 4003 1534 4007
rect 2546 4003 2550 4007
rect 2554 4003 2557 4007
rect 2557 4003 2558 4007
rect 3570 4003 3574 4007
rect 3578 4003 3581 4007
rect 3581 4003 3582 4007
rect 1398 3998 1402 4002
rect 2566 3998 2570 4002
rect 2750 3998 2754 4002
rect 2830 3998 2834 4002
rect 3806 3998 3810 4002
rect 174 3988 178 3992
rect 302 3988 306 3992
rect 1774 3988 1778 3992
rect 1958 3988 1962 3992
rect 1982 3988 1986 3992
rect 2118 3988 2122 3992
rect 3270 3988 3274 3992
rect 174 3978 178 3982
rect 1918 3978 1922 3982
rect 2422 3978 2426 3982
rect 3406 3978 3410 3982
rect 3790 3978 3794 3982
rect 4022 3978 4026 3982
rect 4214 3978 4218 3982
rect 646 3968 650 3972
rect 838 3968 842 3972
rect 2110 3968 2114 3972
rect 2830 3968 2834 3972
rect 3110 3968 3114 3972
rect 4430 3968 4434 3972
rect 486 3958 490 3962
rect 838 3958 842 3962
rect 1518 3958 1522 3962
rect 1806 3958 1810 3962
rect 1910 3958 1914 3962
rect 2174 3958 2178 3962
rect 2198 3958 2202 3962
rect 2630 3958 2634 3962
rect 342 3948 346 3952
rect 422 3948 426 3952
rect 1270 3948 1274 3952
rect 3854 3958 3858 3962
rect 3894 3958 3898 3962
rect 3902 3958 3906 3962
rect 4254 3958 4258 3962
rect 4478 3958 4482 3962
rect 4598 3958 4602 3962
rect 1662 3948 1666 3952
rect 1998 3948 2002 3952
rect 2182 3948 2186 3952
rect 2926 3948 2930 3952
rect 638 3938 642 3942
rect 766 3938 770 3942
rect 798 3938 802 3942
rect 2766 3938 2770 3942
rect 3606 3948 3610 3952
rect 3726 3948 3730 3952
rect 3870 3948 3874 3952
rect 3886 3948 3890 3952
rect 3974 3948 3978 3952
rect 4414 3948 4418 3952
rect 4558 3948 4562 3952
rect 3230 3938 3234 3942
rect 3430 3938 3434 3942
rect 3622 3938 3626 3942
rect 3814 3938 3818 3942
rect 3966 3938 3970 3942
rect 4366 3938 4370 3942
rect 4438 3938 4442 3942
rect 4470 3938 4474 3942
rect 478 3928 482 3932
rect 1302 3928 1306 3932
rect 1966 3928 1970 3932
rect 2382 3928 2386 3932
rect 2622 3928 2626 3932
rect 3590 3928 3594 3932
rect 3838 3928 3842 3932
rect 4286 3928 4290 3932
rect 446 3918 450 3922
rect 2086 3918 2090 3922
rect 3198 3918 3202 3922
rect 3814 3918 3818 3922
rect 3934 3918 3938 3922
rect 4294 3918 4298 3922
rect 270 3908 274 3912
rect 1918 3908 1922 3912
rect 2270 3908 2274 3912
rect 2718 3908 2722 3912
rect 3870 3908 3874 3912
rect 4070 3908 4074 3912
rect 4534 3908 4538 3912
rect 1002 3903 1006 3907
rect 1010 3903 1013 3907
rect 1013 3903 1014 3907
rect 2026 3903 2030 3907
rect 2034 3903 2037 3907
rect 2037 3903 2038 3907
rect 3050 3903 3054 3907
rect 3058 3903 3061 3907
rect 3061 3903 3062 3907
rect 4082 3903 4086 3907
rect 4090 3903 4093 3907
rect 4093 3903 4094 3907
rect 1110 3898 1114 3902
rect 2574 3898 2578 3902
rect 2814 3898 2818 3902
rect 3590 3898 3594 3902
rect 574 3888 578 3892
rect 934 3888 938 3892
rect 1494 3888 1498 3892
rect 1502 3888 1506 3892
rect 2406 3888 2410 3892
rect 3814 3888 3818 3892
rect 4230 3888 4234 3892
rect 4550 3888 4554 3892
rect 422 3878 426 3882
rect 718 3878 722 3882
rect 2246 3878 2250 3882
rect 2390 3878 2394 3882
rect 2494 3878 2498 3882
rect 2710 3878 2714 3882
rect 2902 3878 2906 3882
rect 3494 3878 3498 3882
rect 4422 3878 4426 3882
rect 342 3868 346 3872
rect 1494 3868 1498 3872
rect 2086 3868 2090 3872
rect 2174 3868 2178 3872
rect 2494 3868 2498 3872
rect 2502 3868 2506 3872
rect 2870 3868 2874 3872
rect 382 3858 386 3862
rect 838 3858 842 3862
rect 1406 3858 1410 3862
rect 2902 3858 2906 3862
rect 3790 3868 3794 3872
rect 3918 3868 3922 3872
rect 3934 3868 3938 3872
rect 3950 3868 3954 3872
rect 4046 3868 4050 3872
rect 4406 3868 4410 3872
rect 3294 3858 3298 3862
rect 3302 3858 3306 3862
rect 3518 3858 3522 3862
rect 4374 3858 4378 3862
rect 4398 3858 4402 3862
rect 4526 3858 4530 3862
rect 4558 3858 4562 3862
rect 1966 3848 1970 3852
rect 2502 3848 2506 3852
rect 2542 3848 2546 3852
rect 2566 3848 2570 3852
rect 3078 3848 3082 3852
rect 3430 3848 3434 3852
rect 3870 3848 3874 3852
rect 4550 3848 4554 3852
rect 1030 3838 1034 3842
rect 1478 3838 1482 3842
rect 1958 3838 1962 3842
rect 2006 3838 2010 3842
rect 2238 3838 2242 3842
rect 2870 3838 2874 3842
rect 3710 3838 3714 3842
rect 4438 3838 4442 3842
rect 2278 3828 2282 3832
rect 4270 3828 4274 3832
rect 966 3818 970 3822
rect 2110 3818 2114 3822
rect 2374 3818 2378 3822
rect 4334 3818 4338 3822
rect 2758 3808 2762 3812
rect 3174 3808 3178 3812
rect 4598 3808 4602 3812
rect 498 3803 502 3807
rect 506 3803 509 3807
rect 509 3803 510 3807
rect 1522 3803 1526 3807
rect 1530 3803 1533 3807
rect 1533 3803 1534 3807
rect 2546 3803 2550 3807
rect 2554 3803 2557 3807
rect 2557 3803 2558 3807
rect 3570 3803 3574 3807
rect 3578 3803 3581 3807
rect 3581 3803 3582 3807
rect 478 3798 482 3802
rect 1278 3798 1282 3802
rect 1918 3798 1922 3802
rect 2302 3798 2306 3802
rect 2534 3798 2538 3802
rect 2830 3798 2834 3802
rect 3006 3798 3010 3802
rect 238 3788 242 3792
rect 614 3788 618 3792
rect 1398 3788 1402 3792
rect 2118 3788 2122 3792
rect 2366 3788 2370 3792
rect 3278 3788 3282 3792
rect 1382 3778 1386 3782
rect 3230 3778 3234 3782
rect 3790 3778 3794 3782
rect 3854 3778 3858 3782
rect 3894 3778 3898 3782
rect 566 3768 570 3772
rect 2350 3768 2354 3772
rect 2366 3768 2370 3772
rect 2534 3768 2538 3772
rect 3910 3768 3914 3772
rect 4358 3768 4362 3772
rect 2254 3758 2258 3762
rect 2526 3758 2530 3762
rect 3342 3758 3346 3762
rect 4070 3758 4074 3762
rect 4294 3758 4298 3762
rect 4318 3758 4322 3762
rect 710 3748 714 3752
rect 1062 3748 1066 3752
rect 406 3738 410 3742
rect 774 3738 778 3742
rect 1902 3748 1906 3752
rect 2054 3748 2058 3752
rect 2718 3748 2722 3752
rect 3094 3748 3098 3752
rect 4054 3748 4058 3752
rect 4262 3748 4266 3752
rect 4350 3748 4354 3752
rect 4382 3748 4386 3752
rect 4598 3748 4602 3752
rect 1398 3738 1402 3742
rect 2070 3738 2074 3742
rect 2534 3738 2538 3742
rect 2998 3738 3002 3742
rect 766 3728 770 3732
rect 2358 3728 2362 3732
rect 2662 3728 2666 3732
rect 4286 3728 4290 3732
rect 4438 3728 4442 3732
rect 4470 3728 4474 3732
rect 4566 3728 4570 3732
rect 2342 3718 2346 3722
rect 3798 3718 3802 3722
rect 4414 3718 4418 3722
rect 4582 3718 4586 3722
rect 1022 3708 1026 3712
rect 1846 3708 1850 3712
rect 2334 3708 2338 3712
rect 2606 3708 2610 3712
rect 2734 3708 2738 3712
rect 3110 3708 3114 3712
rect 3398 3708 3402 3712
rect 1002 3703 1006 3707
rect 1010 3703 1013 3707
rect 1013 3703 1014 3707
rect 2026 3703 2030 3707
rect 2034 3703 2037 3707
rect 2037 3703 2038 3707
rect 3050 3703 3054 3707
rect 3058 3703 3061 3707
rect 3061 3703 3062 3707
rect 4082 3703 4086 3707
rect 4090 3703 4093 3707
rect 4093 3703 4094 3707
rect 1798 3698 1802 3702
rect 1958 3698 1962 3702
rect 2270 3698 2274 3702
rect 2870 3698 2874 3702
rect 4118 3698 4122 3702
rect 358 3688 362 3692
rect 814 3688 818 3692
rect 1038 3688 1042 3692
rect 1110 3688 1114 3692
rect 2454 3688 2458 3692
rect 2694 3688 2698 3692
rect 2718 3688 2722 3692
rect 2742 3688 2746 3692
rect 3486 3688 3490 3692
rect 3494 3688 3498 3692
rect 4190 3688 4194 3692
rect 4326 3688 4330 3692
rect 166 3678 170 3682
rect 2326 3678 2330 3682
rect 2718 3678 2722 3682
rect 2766 3678 2770 3682
rect 2894 3678 2898 3682
rect 382 3668 386 3672
rect 2150 3668 2154 3672
rect 2734 3668 2738 3672
rect 2934 3668 2938 3672
rect 2950 3668 2954 3672
rect 3102 3668 3106 3672
rect 3118 3668 3122 3672
rect 3182 3668 3186 3672
rect 3206 3668 3210 3672
rect 3222 3668 3226 3672
rect 4102 3668 4106 3672
rect 4462 3668 4466 3672
rect 542 3658 546 3662
rect 910 3658 914 3662
rect 1054 3658 1058 3662
rect 1590 3658 1594 3662
rect 1846 3658 1850 3662
rect 1958 3658 1962 3662
rect 2134 3658 2138 3662
rect 2470 3658 2474 3662
rect 2710 3658 2714 3662
rect 2750 3658 2754 3662
rect 2846 3658 2850 3662
rect 2870 3658 2874 3662
rect 3550 3658 3554 3662
rect 3742 3658 3746 3662
rect 4030 3658 4034 3662
rect 4262 3658 4266 3662
rect 798 3648 802 3652
rect 1990 3648 1994 3652
rect 2270 3648 2274 3652
rect 2518 3648 2522 3652
rect 2558 3648 2562 3652
rect 2862 3648 2866 3652
rect 3014 3648 3018 3652
rect 3102 3648 3106 3652
rect 4190 3648 4194 3652
rect 4526 3648 4530 3652
rect 782 3638 786 3642
rect 1790 3638 1794 3642
rect 2014 3638 2018 3642
rect 2574 3638 2578 3642
rect 2838 3638 2842 3642
rect 4318 3638 4322 3642
rect 4334 3638 4338 3642
rect 4478 3638 4482 3642
rect 2102 3628 2106 3632
rect 2430 3628 2434 3632
rect 2590 3628 2594 3632
rect 3886 3628 3890 3632
rect 2134 3618 2138 3622
rect 2262 3618 2266 3622
rect 2990 3618 2994 3622
rect 3214 3618 3218 3622
rect 4374 3618 4378 3622
rect 3590 3608 3594 3612
rect 498 3603 502 3607
rect 506 3603 509 3607
rect 509 3603 510 3607
rect 1522 3603 1526 3607
rect 1530 3603 1533 3607
rect 1533 3603 1534 3607
rect 2546 3603 2550 3607
rect 2554 3603 2557 3607
rect 2557 3603 2558 3607
rect 3570 3603 3574 3607
rect 3578 3603 3581 3607
rect 3581 3603 3582 3607
rect 1798 3598 1802 3602
rect 2438 3598 2442 3602
rect 2494 3598 2498 3602
rect 2502 3598 2506 3602
rect 2590 3598 2594 3602
rect 3406 3598 3410 3602
rect 3774 3598 3778 3602
rect 2214 3588 2218 3592
rect 2766 3588 2770 3592
rect 3542 3588 3546 3592
rect 4222 3588 4226 3592
rect 406 3578 410 3582
rect 2838 3578 2842 3582
rect 3358 3578 3362 3582
rect 3470 3578 3474 3582
rect 2454 3568 2458 3572
rect 2486 3568 2490 3572
rect 2502 3568 2506 3572
rect 2630 3568 2634 3572
rect 2774 3568 2778 3572
rect 3094 3568 3098 3572
rect 3326 3568 3330 3572
rect 3814 3568 3818 3572
rect 3886 3568 3890 3572
rect 4430 3568 4434 3572
rect 462 3558 466 3562
rect 798 3558 802 3562
rect 2166 3558 2170 3562
rect 2390 3558 2394 3562
rect 2670 3558 2674 3562
rect 2718 3558 2722 3562
rect 3382 3558 3386 3562
rect 3430 3558 3434 3562
rect 3902 3558 3906 3562
rect 398 3548 402 3552
rect 1078 3548 1082 3552
rect 566 3538 570 3542
rect 1398 3548 1402 3552
rect 1494 3548 1498 3552
rect 1518 3548 1522 3552
rect 1814 3548 1818 3552
rect 1982 3548 1986 3552
rect 2638 3548 2642 3552
rect 2846 3548 2850 3552
rect 3486 3548 3490 3552
rect 3742 3548 3746 3552
rect 2310 3538 2314 3542
rect 2326 3538 2330 3542
rect 2414 3538 2418 3542
rect 2654 3538 2658 3542
rect 2894 3538 2898 3542
rect 3294 3538 3298 3542
rect 4214 3538 4218 3542
rect 4494 3538 4498 3542
rect 2006 3528 2010 3532
rect 2422 3528 2426 3532
rect 2478 3528 2482 3532
rect 726 3518 730 3522
rect 1950 3518 1954 3522
rect 2270 3518 2274 3522
rect 2390 3518 2394 3522
rect 2518 3518 2522 3522
rect 2870 3518 2874 3522
rect 3310 3518 3314 3522
rect 3334 3518 3338 3522
rect 3462 3518 3466 3522
rect 3886 3518 3890 3522
rect 1982 3508 1986 3512
rect 2350 3508 2354 3512
rect 2414 3508 2418 3512
rect 1002 3503 1006 3507
rect 1010 3503 1013 3507
rect 1013 3503 1014 3507
rect 2026 3503 2030 3507
rect 2034 3503 2037 3507
rect 2037 3503 2038 3507
rect 3050 3503 3054 3507
rect 3058 3503 3061 3507
rect 3061 3503 3062 3507
rect 4082 3503 4086 3507
rect 4090 3503 4093 3507
rect 4093 3503 4094 3507
rect 2654 3498 2658 3502
rect 2918 3498 2922 3502
rect 4070 3498 4074 3502
rect 4102 3498 4106 3502
rect 1022 3488 1026 3492
rect 1782 3488 1786 3492
rect 1918 3488 1922 3492
rect 1966 3488 1970 3492
rect 2230 3488 2234 3492
rect 2686 3488 2690 3492
rect 3502 3488 3506 3492
rect 470 3478 474 3482
rect 830 3478 834 3482
rect 2094 3478 2098 3482
rect 2910 3478 2914 3482
rect 3790 3478 3794 3482
rect 4318 3478 4322 3482
rect 1942 3468 1946 3472
rect 2022 3468 2026 3472
rect 2486 3468 2490 3472
rect 2646 3468 2650 3472
rect 2870 3468 2874 3472
rect 2942 3468 2946 3472
rect 3022 3468 3026 3472
rect 3830 3468 3834 3472
rect 230 3458 234 3462
rect 3078 3458 3082 3462
rect 3102 3458 3106 3462
rect 3142 3458 3146 3462
rect 3166 3458 3170 3462
rect 3214 3458 3218 3462
rect 3350 3458 3354 3462
rect 3366 3458 3370 3462
rect 3846 3458 3850 3462
rect 3942 3458 3946 3462
rect 4030 3458 4034 3462
rect 254 3448 258 3452
rect 462 3448 466 3452
rect 2798 3448 2802 3452
rect 2886 3448 2890 3452
rect 2934 3448 2938 3452
rect 3014 3448 3018 3452
rect 3462 3448 3466 3452
rect 3614 3448 3618 3452
rect 1590 3438 1594 3442
rect 2390 3438 2394 3442
rect 2686 3438 2690 3442
rect 2838 3438 2842 3442
rect 4510 3438 4514 3442
rect 1230 3428 1234 3432
rect 2366 3428 2370 3432
rect 2430 3428 2434 3432
rect 2670 3428 2674 3432
rect 2998 3428 3002 3432
rect 3598 3428 3602 3432
rect 2502 3418 2506 3422
rect 1806 3408 1810 3412
rect 2686 3408 2690 3412
rect 3038 3408 3042 3412
rect 3318 3408 3322 3412
rect 498 3403 502 3407
rect 506 3403 509 3407
rect 509 3403 510 3407
rect 1522 3403 1526 3407
rect 1530 3403 1533 3407
rect 1533 3403 1534 3407
rect 2546 3403 2550 3407
rect 2554 3403 2557 3407
rect 2557 3403 2558 3407
rect 3570 3403 3574 3407
rect 3578 3403 3581 3407
rect 3581 3403 3582 3407
rect 2214 3398 2218 3402
rect 2302 3398 2306 3402
rect 2830 3398 2834 3402
rect 3134 3398 3138 3402
rect 2254 3388 2258 3392
rect 2334 3388 2338 3392
rect 2430 3388 2434 3392
rect 2526 3388 2530 3392
rect 2678 3388 2682 3392
rect 2822 3388 2826 3392
rect 2838 3388 2842 3392
rect 3094 3388 3098 3392
rect 4110 3388 4114 3392
rect 4174 3388 4178 3392
rect 2446 3378 2450 3382
rect 2734 3378 2738 3382
rect 2894 3378 2898 3382
rect 2958 3378 2962 3382
rect 3110 3378 3114 3382
rect 3150 3378 3154 3382
rect 3190 3378 3194 3382
rect 3478 3378 3482 3382
rect 4494 3378 4498 3382
rect 2246 3368 2250 3372
rect 2318 3368 2322 3372
rect 2414 3368 2418 3372
rect 2518 3368 2522 3372
rect 2782 3368 2786 3372
rect 2814 3368 2818 3372
rect 1990 3358 1994 3362
rect 2110 3358 2114 3362
rect 2262 3358 2266 3362
rect 2934 3358 2938 3362
rect 2966 3358 2970 3362
rect 3006 3358 3010 3362
rect 3158 3358 3162 3362
rect 3166 3358 3170 3362
rect 3198 3358 3202 3362
rect 3278 3358 3282 3362
rect 3374 3358 3378 3362
rect 158 3348 162 3352
rect 470 3348 474 3352
rect 1134 3348 1138 3352
rect 1478 3348 1482 3352
rect 1766 3348 1770 3352
rect 2294 3348 2298 3352
rect 2374 3348 2378 3352
rect 2918 3348 2922 3352
rect 2990 3348 2994 3352
rect 3446 3348 3450 3352
rect 3534 3348 3538 3352
rect 3782 3348 3786 3352
rect 934 3338 938 3342
rect 2094 3338 2098 3342
rect 2406 3338 2410 3342
rect 2878 3338 2882 3342
rect 2974 3338 2978 3342
rect 3254 3338 3258 3342
rect 3286 3338 3290 3342
rect 4318 3338 4322 3342
rect 646 3328 650 3332
rect 726 3328 730 3332
rect 2374 3328 2378 3332
rect 2398 3328 2402 3332
rect 2526 3328 2530 3332
rect 2798 3328 2802 3332
rect 3126 3328 3130 3332
rect 3310 3328 3314 3332
rect 3318 3328 3322 3332
rect 438 3318 442 3322
rect 614 3318 618 3322
rect 798 3318 802 3322
rect 2126 3318 2130 3322
rect 2286 3318 2290 3322
rect 2366 3318 2370 3322
rect 2486 3318 2490 3322
rect 2550 3318 2554 3322
rect 2630 3318 2634 3322
rect 2694 3318 2698 3322
rect 2790 3318 2794 3322
rect 2830 3318 2834 3322
rect 2974 3318 2978 3322
rect 3070 3318 3074 3322
rect 3166 3318 3170 3322
rect 3206 3318 3210 3322
rect 3326 3318 3330 3322
rect 1686 3308 1690 3312
rect 2398 3308 2402 3312
rect 2702 3308 2706 3312
rect 2878 3308 2882 3312
rect 2910 3308 2914 3312
rect 3702 3308 3706 3312
rect 4502 3308 4506 3312
rect 1002 3303 1006 3307
rect 1010 3303 1013 3307
rect 1013 3303 1014 3307
rect 2026 3303 2030 3307
rect 2034 3303 2037 3307
rect 2037 3303 2038 3307
rect 3050 3303 3054 3307
rect 3058 3303 3061 3307
rect 3061 3303 3062 3307
rect 4082 3303 4086 3307
rect 4090 3303 4093 3307
rect 4093 3303 4094 3307
rect 742 3298 746 3302
rect 2342 3298 2346 3302
rect 2566 3298 2570 3302
rect 2886 3298 2890 3302
rect 2934 3298 2938 3302
rect 3102 3298 3106 3302
rect 3950 3298 3954 3302
rect 718 3288 722 3292
rect 1934 3288 1938 3292
rect 2014 3288 2018 3292
rect 2286 3288 2290 3292
rect 2534 3288 2538 3292
rect 2638 3288 2642 3292
rect 3022 3288 3026 3292
rect 3110 3288 3114 3292
rect 4390 3288 4394 3292
rect 494 3278 498 3282
rect 2182 3278 2186 3282
rect 2942 3278 2946 3282
rect 2982 3278 2986 3282
rect 3430 3278 3434 3282
rect 294 3268 298 3272
rect 318 3268 322 3272
rect 1934 3268 1938 3272
rect 2214 3268 2218 3272
rect 2254 3268 2258 3272
rect 2342 3268 2346 3272
rect 2670 3268 2674 3272
rect 2942 3268 2946 3272
rect 3262 3268 3266 3272
rect 3278 3268 3282 3272
rect 3302 3268 3306 3272
rect 3310 3268 3314 3272
rect 3398 3268 3402 3272
rect 4118 3268 4122 3272
rect 4214 3268 4218 3272
rect 366 3258 370 3262
rect 1862 3258 1866 3262
rect 2094 3258 2098 3262
rect 2262 3258 2266 3262
rect 2302 3258 2306 3262
rect 2598 3258 2602 3262
rect 2614 3258 2618 3262
rect 2910 3258 2914 3262
rect 2958 3258 2962 3262
rect 3694 3258 3698 3262
rect 4526 3258 4530 3262
rect 1350 3248 1354 3252
rect 1382 3248 1386 3252
rect 1774 3248 1778 3252
rect 2350 3248 2354 3252
rect 2390 3238 2394 3242
rect 2630 3238 2634 3242
rect 2966 3238 2970 3242
rect 4262 3238 4266 3242
rect 1342 3228 1346 3232
rect 1406 3228 1410 3232
rect 2798 3228 2802 3232
rect 3438 3228 3442 3232
rect 3454 3228 3458 3232
rect 806 3218 810 3222
rect 2822 3218 2826 3222
rect 2878 3218 2882 3222
rect 4102 3218 4106 3222
rect 766 3208 770 3212
rect 1102 3208 1106 3212
rect 1406 3208 1410 3212
rect 1478 3208 1482 3212
rect 2158 3208 2162 3212
rect 2326 3208 2330 3212
rect 3270 3208 3274 3212
rect 4326 3208 4330 3212
rect 498 3203 502 3207
rect 506 3203 509 3207
rect 509 3203 510 3207
rect 1522 3203 1526 3207
rect 1530 3203 1533 3207
rect 1533 3203 1534 3207
rect 2546 3203 2550 3207
rect 2554 3203 2557 3207
rect 2557 3203 2558 3207
rect 3570 3203 3574 3207
rect 3578 3203 3581 3207
rect 3581 3203 3582 3207
rect 1414 3198 1418 3202
rect 2286 3198 2290 3202
rect 2342 3198 2346 3202
rect 2350 3198 2354 3202
rect 2502 3198 2506 3202
rect 2574 3198 2578 3202
rect 3294 3198 3298 3202
rect 4406 3198 4410 3202
rect 2158 3188 2162 3192
rect 2854 3188 2858 3192
rect 3710 3188 3714 3192
rect 3958 3188 3962 3192
rect 2270 3178 2274 3182
rect 2806 3178 2810 3182
rect 2838 3178 2842 3182
rect 2918 3178 2922 3182
rect 3030 3178 3034 3182
rect 3174 3178 3178 3182
rect 3286 3178 3290 3182
rect 30 3168 34 3172
rect 302 3168 306 3172
rect 814 3168 818 3172
rect 2222 3168 2226 3172
rect 2310 3168 2314 3172
rect 2454 3168 2458 3172
rect 2478 3168 2482 3172
rect 2494 3168 2498 3172
rect 2662 3168 2666 3172
rect 2734 3168 2738 3172
rect 3014 3168 3018 3172
rect 3110 3168 3114 3172
rect 3158 3168 3162 3172
rect 2382 3158 2386 3162
rect 2646 3158 2650 3162
rect 2662 3158 2666 3162
rect 2758 3158 2762 3162
rect 2830 3158 2834 3162
rect 3878 3158 3882 3162
rect 4446 3158 4450 3162
rect 150 3148 154 3152
rect 726 3148 730 3152
rect 1686 3148 1690 3152
rect 1806 3148 1810 3152
rect 1990 3148 1994 3152
rect 2062 3148 2066 3152
rect 2406 3148 2410 3152
rect 2854 3148 2858 3152
rect 2862 3148 2866 3152
rect 2878 3148 2882 3152
rect 1406 3138 1410 3142
rect 1606 3138 1610 3142
rect 2078 3138 2082 3142
rect 4334 3148 4338 3152
rect 4478 3148 4482 3152
rect 4510 3148 4514 3152
rect 2494 3138 2498 3142
rect 2622 3138 2626 3142
rect 3670 3138 3674 3142
rect 4046 3138 4050 3142
rect 4118 3138 4122 3142
rect 4374 3138 4378 3142
rect 4438 3138 4442 3142
rect 4566 3138 4570 3142
rect 1566 3128 1570 3132
rect 1574 3128 1578 3132
rect 2350 3128 2354 3132
rect 2846 3128 2850 3132
rect 2870 3128 2874 3132
rect 2942 3128 2946 3132
rect 2990 3128 2994 3132
rect 3134 3128 3138 3132
rect 3246 3128 3250 3132
rect 254 3118 258 3122
rect 662 3118 666 3122
rect 1302 3118 1306 3122
rect 1678 3118 1682 3122
rect 2462 3118 2466 3122
rect 2486 3118 2490 3122
rect 2494 3118 2498 3122
rect 2622 3118 2626 3122
rect 2774 3118 2778 3122
rect 3030 3118 3034 3122
rect 3294 3118 3298 3122
rect 2310 3108 2314 3112
rect 2358 3108 2362 3112
rect 2438 3108 2442 3112
rect 3254 3108 3258 3112
rect 3646 3108 3650 3112
rect 4438 3108 4442 3112
rect 1002 3103 1006 3107
rect 1010 3103 1013 3107
rect 1013 3103 1014 3107
rect 2026 3103 2030 3107
rect 2034 3103 2037 3107
rect 2037 3103 2038 3107
rect 3050 3103 3054 3107
rect 3058 3103 3061 3107
rect 3061 3103 3062 3107
rect 4082 3103 4086 3107
rect 4090 3103 4093 3107
rect 4093 3103 4094 3107
rect 398 3098 402 3102
rect 2150 3098 2154 3102
rect 2646 3098 2650 3102
rect 2694 3098 2698 3102
rect 2862 3098 2866 3102
rect 3254 3098 3258 3102
rect 854 3088 858 3092
rect 1294 3088 1298 3092
rect 1790 3088 1794 3092
rect 1886 3088 1890 3092
rect 1998 3088 2002 3092
rect 2070 3088 2074 3092
rect 2390 3088 2394 3092
rect 2438 3088 2442 3092
rect 3030 3088 3034 3092
rect 686 3078 690 3082
rect 750 3078 754 3082
rect 1670 3078 1674 3082
rect 2214 3078 2218 3082
rect 2270 3078 2274 3082
rect 2534 3078 2538 3082
rect 2822 3078 2826 3082
rect 3150 3078 3154 3082
rect 4406 3078 4410 3082
rect 6 3068 10 3072
rect 566 3068 570 3072
rect 1382 3068 1386 3072
rect 2254 3068 2258 3072
rect 2318 3068 2322 3072
rect 2422 3068 2426 3072
rect 2486 3068 2490 3072
rect 2902 3068 2906 3072
rect 3110 3068 3114 3072
rect 3358 3068 3362 3072
rect 4534 3068 4538 3072
rect 542 3058 546 3062
rect 750 3058 754 3062
rect 1558 3058 1562 3062
rect 1854 3058 1858 3062
rect 2046 3058 2050 3062
rect 2654 3058 2658 3062
rect 2918 3058 2922 3062
rect 3006 3058 3010 3062
rect 3118 3058 3122 3062
rect 3142 3058 3146 3062
rect 3174 3058 3178 3062
rect 3206 3058 3210 3062
rect 3486 3058 3490 3062
rect 3798 3058 3802 3062
rect 6 3048 10 3052
rect 654 3048 658 3052
rect 2366 3048 2370 3052
rect 2910 3048 2914 3052
rect 3166 3048 3170 3052
rect 3318 3048 3322 3052
rect 4366 3048 4370 3052
rect 30 3038 34 3042
rect 150 3038 154 3042
rect 302 3038 306 3042
rect 2118 3038 2122 3042
rect 3126 3038 3130 3042
rect 3366 3038 3370 3042
rect 4534 3038 4538 3042
rect 782 3028 786 3032
rect 2286 3028 2290 3032
rect 2726 3028 2730 3032
rect 2766 3028 2770 3032
rect 2846 3028 2850 3032
rect 3182 3028 3186 3032
rect 4254 3028 4258 3032
rect 1582 3018 1586 3022
rect 2214 3018 2218 3022
rect 2486 3018 2490 3022
rect 3406 3018 3410 3022
rect 3486 3018 3490 3022
rect 3678 3018 3682 3022
rect 2206 3008 2210 3012
rect 2534 3008 2538 3012
rect 2774 3008 2778 3012
rect 498 3003 502 3007
rect 506 3003 509 3007
rect 509 3003 510 3007
rect 1522 3003 1526 3007
rect 1530 3003 1533 3007
rect 1533 3003 1534 3007
rect 398 2998 402 3002
rect 630 2998 634 3002
rect 1286 2998 1290 3002
rect 1862 2998 1866 3002
rect 2546 3003 2550 3007
rect 2554 3003 2557 3007
rect 2557 3003 2558 3007
rect 3570 3003 3574 3007
rect 3578 3003 3581 3007
rect 3581 3003 3582 3007
rect 2174 2998 2178 3002
rect 2390 2998 2394 3002
rect 2934 2998 2938 3002
rect 158 2988 162 2992
rect 3286 2988 3290 2992
rect 398 2978 402 2982
rect 2206 2978 2210 2982
rect 2342 2978 2346 2982
rect 3478 2978 3482 2982
rect 4118 2978 4122 2982
rect 2246 2968 2250 2972
rect 2374 2968 2378 2972
rect 3030 2968 3034 2972
rect 3694 2968 3698 2972
rect 4566 2968 4570 2972
rect 742 2958 746 2962
rect 2566 2958 2570 2962
rect 2782 2958 2786 2962
rect 2918 2958 2922 2962
rect 3246 2958 3250 2962
rect 4326 2958 4330 2962
rect 4550 2958 4554 2962
rect 566 2948 570 2952
rect 646 2948 650 2952
rect 1222 2948 1226 2952
rect 750 2938 754 2942
rect 1534 2948 1538 2952
rect 2014 2948 2018 2952
rect 2030 2948 2034 2952
rect 1062 2938 1066 2942
rect 2230 2948 2234 2952
rect 2398 2948 2402 2952
rect 2614 2948 2618 2952
rect 2110 2938 2114 2942
rect 2150 2938 2154 2942
rect 2278 2938 2282 2942
rect 2454 2938 2458 2942
rect 4318 2938 4322 2942
rect 2494 2928 2498 2932
rect 2518 2928 2522 2932
rect 2854 2928 2858 2932
rect 3078 2928 3082 2932
rect 3110 2928 3114 2932
rect 1606 2918 1610 2922
rect 1886 2918 1890 2922
rect 2454 2918 2458 2922
rect 2750 2918 2754 2922
rect 2910 2918 2914 2922
rect 3246 2918 3250 2922
rect 3534 2918 3538 2922
rect 462 2908 466 2912
rect 654 2908 658 2912
rect 2686 2908 2690 2912
rect 2894 2908 2898 2912
rect 2966 2908 2970 2912
rect 3278 2908 3282 2912
rect 1002 2903 1006 2907
rect 1010 2903 1013 2907
rect 1013 2903 1014 2907
rect 2026 2903 2030 2907
rect 2034 2903 2037 2907
rect 2037 2903 2038 2907
rect 3050 2903 3054 2907
rect 3058 2903 3061 2907
rect 3061 2903 3062 2907
rect 4082 2903 4086 2907
rect 4090 2903 4093 2907
rect 4093 2903 4094 2907
rect 366 2898 370 2902
rect 1902 2898 1906 2902
rect 2046 2898 2050 2902
rect 2646 2898 2650 2902
rect 3006 2898 3010 2902
rect 3814 2898 3818 2902
rect 438 2888 442 2892
rect 694 2888 698 2892
rect 870 2888 874 2892
rect 1382 2888 1386 2892
rect 1910 2888 1914 2892
rect 1926 2888 1930 2892
rect 2350 2888 2354 2892
rect 2518 2888 2522 2892
rect 2846 2888 2850 2892
rect 3302 2888 3306 2892
rect 3342 2888 3346 2892
rect 3494 2888 3498 2892
rect 4262 2888 4266 2892
rect 662 2878 666 2882
rect 878 2878 882 2882
rect 2158 2878 2162 2882
rect 2862 2878 2866 2882
rect 3078 2878 3082 2882
rect 3686 2878 3690 2882
rect 1646 2868 1650 2872
rect 2350 2868 2354 2872
rect 2462 2868 2466 2872
rect 2630 2868 2634 2872
rect 2878 2868 2882 2872
rect 4598 2868 4602 2872
rect 686 2858 690 2862
rect 710 2858 714 2862
rect 814 2858 818 2862
rect 1030 2858 1034 2862
rect 1582 2858 1586 2862
rect 2310 2858 2314 2862
rect 2406 2858 2410 2862
rect 2502 2858 2506 2862
rect 2590 2858 2594 2862
rect 2614 2858 2618 2862
rect 2758 2858 2762 2862
rect 3070 2858 3074 2862
rect 3662 2858 3666 2862
rect 4446 2858 4450 2862
rect 4550 2858 4554 2862
rect 2118 2848 2122 2852
rect 2886 2848 2890 2852
rect 1046 2838 1050 2842
rect 2566 2838 2570 2842
rect 2790 2838 2794 2842
rect 3662 2838 3666 2842
rect 4566 2838 4570 2842
rect 2086 2828 2090 2832
rect 2158 2828 2162 2832
rect 2350 2828 2354 2832
rect 2422 2828 2426 2832
rect 3742 2828 3746 2832
rect 814 2818 818 2822
rect 4438 2818 4442 2822
rect 2478 2808 2482 2812
rect 2574 2808 2578 2812
rect 498 2803 502 2807
rect 506 2803 509 2807
rect 509 2803 510 2807
rect 1522 2803 1526 2807
rect 1530 2803 1533 2807
rect 1533 2803 1534 2807
rect 2546 2803 2550 2807
rect 2554 2803 2557 2807
rect 2557 2803 2558 2807
rect 3570 2803 3574 2807
rect 3578 2803 3581 2807
rect 3581 2803 3582 2807
rect 1486 2798 1490 2802
rect 2294 2798 2298 2802
rect 862 2788 866 2792
rect 1406 2788 1410 2792
rect 3150 2788 3154 2792
rect 2094 2778 2098 2782
rect 2566 2778 2570 2782
rect 2934 2778 2938 2782
rect 3358 2778 3362 2782
rect 4598 2778 4602 2782
rect 1686 2768 1690 2772
rect 1902 2768 1906 2772
rect 2126 2768 2130 2772
rect 3998 2768 4002 2772
rect 694 2758 698 2762
rect 2006 2758 2010 2762
rect 2110 2758 2114 2762
rect 2526 2758 2530 2762
rect 2614 2758 2618 2762
rect 3510 2758 3514 2762
rect 638 2748 642 2752
rect 710 2748 714 2752
rect 734 2748 738 2752
rect 894 2748 898 2752
rect 1414 2748 1418 2752
rect 614 2738 618 2742
rect 2326 2748 2330 2752
rect 2902 2748 2906 2752
rect 2310 2738 2314 2742
rect 4230 2738 4234 2742
rect 2110 2728 2114 2732
rect 2494 2728 2498 2732
rect 2734 2728 2738 2732
rect 3774 2728 3778 2732
rect 4054 2728 4058 2732
rect 318 2718 322 2722
rect 694 2718 698 2722
rect 2910 2718 2914 2722
rect 2462 2708 2466 2712
rect 2998 2708 3002 2712
rect 3262 2708 3266 2712
rect 4206 2708 4210 2712
rect 1002 2703 1006 2707
rect 1010 2703 1013 2707
rect 1013 2703 1014 2707
rect 2026 2703 2030 2707
rect 2034 2703 2037 2707
rect 2037 2703 2038 2707
rect 3050 2703 3054 2707
rect 3058 2703 3061 2707
rect 3061 2703 3062 2707
rect 4082 2703 4086 2707
rect 4090 2703 4093 2707
rect 4093 2703 4094 2707
rect 1638 2698 1642 2702
rect 2406 2698 2410 2702
rect 2670 2698 2674 2702
rect 3126 2698 3130 2702
rect 3670 2698 3674 2702
rect 886 2688 890 2692
rect 1558 2688 1562 2692
rect 2070 2688 2074 2692
rect 2118 2688 2122 2692
rect 2390 2688 2394 2692
rect 2486 2688 2490 2692
rect 2494 2688 2498 2692
rect 3038 2688 3042 2692
rect 3086 2688 3090 2692
rect 3198 2688 3202 2692
rect 3390 2688 3394 2692
rect 3806 2688 3810 2692
rect 646 2678 650 2682
rect 678 2678 682 2682
rect 1726 2678 1730 2682
rect 2454 2678 2458 2682
rect 2614 2678 2618 2682
rect 2878 2678 2882 2682
rect 3142 2678 3146 2682
rect 3678 2678 3682 2682
rect 790 2668 794 2672
rect 1774 2668 1778 2672
rect 3118 2668 3122 2672
rect 3398 2668 3402 2672
rect 3438 2668 3442 2672
rect 3806 2668 3810 2672
rect 4038 2668 4042 2672
rect 318 2658 322 2662
rect 734 2658 738 2662
rect 758 2658 762 2662
rect 830 2658 834 2662
rect 1326 2658 1330 2662
rect 1726 2658 1730 2662
rect 2190 2658 2194 2662
rect 3174 2658 3178 2662
rect 3262 2658 3266 2662
rect 606 2648 610 2652
rect 718 2648 722 2652
rect 1638 2648 1642 2652
rect 2254 2648 2258 2652
rect 2846 2648 2850 2652
rect 3214 2648 3218 2652
rect 3958 2648 3962 2652
rect 4206 2648 4210 2652
rect 2046 2628 2050 2632
rect 2310 2628 2314 2632
rect 2318 2628 2322 2632
rect 2974 2628 2978 2632
rect 2990 2628 2994 2632
rect 2078 2618 2082 2622
rect 2910 2618 2914 2622
rect 3638 2618 3642 2622
rect 1022 2608 1026 2612
rect 2350 2608 2354 2612
rect 2782 2608 2786 2612
rect 498 2603 502 2607
rect 506 2603 509 2607
rect 509 2603 510 2607
rect 1522 2603 1526 2607
rect 1530 2603 1533 2607
rect 1533 2603 1534 2607
rect 2546 2603 2550 2607
rect 2554 2603 2557 2607
rect 2557 2603 2558 2607
rect 3570 2603 3574 2607
rect 3578 2603 3581 2607
rect 3581 2603 3582 2607
rect 2430 2598 2434 2602
rect 1030 2588 1034 2592
rect 1566 2588 1570 2592
rect 1662 2588 1666 2592
rect 1806 2588 1810 2592
rect 2134 2588 2138 2592
rect 2318 2588 2322 2592
rect 2462 2588 2466 2592
rect 2614 2588 2618 2592
rect 2750 2588 2754 2592
rect 3014 2588 3018 2592
rect 2190 2578 2194 2582
rect 2750 2578 2754 2582
rect 3158 2578 3162 2582
rect 3310 2578 3314 2582
rect 3374 2578 3378 2582
rect 3742 2578 3746 2582
rect 2678 2568 2682 2572
rect 2710 2568 2714 2572
rect 2814 2568 2818 2572
rect 2862 2568 2866 2572
rect 2934 2568 2938 2572
rect 3382 2568 3386 2572
rect 4230 2568 4234 2572
rect 4430 2568 4434 2572
rect 630 2558 634 2562
rect 686 2558 690 2562
rect 926 2558 930 2562
rect 1086 2558 1090 2562
rect 2902 2558 2906 2562
rect 3422 2558 3426 2562
rect 3654 2558 3658 2562
rect 3742 2558 3746 2562
rect 4302 2558 4306 2562
rect 54 2548 58 2552
rect 222 2548 226 2552
rect 726 2548 730 2552
rect 1726 2548 1730 2552
rect 1990 2548 1994 2552
rect 2126 2548 2130 2552
rect 2726 2548 2730 2552
rect 3198 2548 3202 2552
rect 3398 2548 3402 2552
rect 4550 2548 4554 2552
rect 2526 2538 2530 2542
rect 2782 2538 2786 2542
rect 2902 2538 2906 2542
rect 3246 2538 3250 2542
rect 3422 2538 3426 2542
rect 3438 2538 3442 2542
rect 3726 2538 3730 2542
rect 4182 2538 4186 2542
rect 4326 2538 4330 2542
rect 1990 2528 1994 2532
rect 2830 2528 2834 2532
rect 2838 2528 2842 2532
rect 3534 2528 3538 2532
rect 3558 2528 3562 2532
rect 3918 2528 3922 2532
rect 4342 2528 4346 2532
rect 478 2518 482 2522
rect 1294 2518 1298 2522
rect 2366 2518 2370 2522
rect 2886 2518 2890 2522
rect 2966 2518 2970 2522
rect 3206 2518 3210 2522
rect 3622 2518 3626 2522
rect 3694 2518 3698 2522
rect 446 2508 450 2512
rect 3526 2508 3530 2512
rect 3734 2508 3738 2512
rect 4190 2508 4194 2512
rect 1002 2503 1006 2507
rect 1010 2503 1013 2507
rect 1013 2503 1014 2507
rect 2026 2503 2030 2507
rect 2034 2503 2037 2507
rect 2037 2503 2038 2507
rect 3050 2503 3054 2507
rect 3058 2503 3061 2507
rect 3061 2503 3062 2507
rect 4082 2503 4086 2507
rect 4090 2503 4093 2507
rect 4093 2503 4094 2507
rect 1358 2498 1362 2502
rect 1662 2498 1666 2502
rect 2214 2498 2218 2502
rect 2390 2498 2394 2502
rect 2606 2498 2610 2502
rect 3070 2498 3074 2502
rect 3238 2498 3242 2502
rect 3350 2498 3354 2502
rect 4182 2498 4186 2502
rect 4318 2498 4322 2502
rect 774 2488 778 2492
rect 1454 2488 1458 2492
rect 1646 2488 1650 2492
rect 1982 2488 1986 2492
rect 2478 2488 2482 2492
rect 2918 2488 2922 2492
rect 3270 2488 3274 2492
rect 1038 2478 1042 2482
rect 2526 2478 2530 2482
rect 2582 2478 2586 2482
rect 2598 2478 2602 2482
rect 2774 2478 2778 2482
rect 2862 2478 2866 2482
rect 3694 2488 3698 2492
rect 4334 2488 4338 2492
rect 3166 2478 3170 2482
rect 3470 2478 3474 2482
rect 3486 2478 3490 2482
rect 3830 2478 3834 2482
rect 4038 2478 4042 2482
rect 4590 2478 4594 2482
rect 918 2468 922 2472
rect 926 2468 930 2472
rect 1006 2468 1010 2472
rect 1198 2468 1202 2472
rect 2318 2468 2322 2472
rect 2334 2468 2338 2472
rect 2758 2468 2762 2472
rect 3590 2468 3594 2472
rect 3646 2468 3650 2472
rect 4142 2468 4146 2472
rect 54 2458 58 2462
rect 694 2458 698 2462
rect 1806 2458 1810 2462
rect 1902 2458 1906 2462
rect 2230 2458 2234 2462
rect 2390 2458 2394 2462
rect 2502 2458 2506 2462
rect 2870 2458 2874 2462
rect 2990 2458 2994 2462
rect 3126 2458 3130 2462
rect 3134 2458 3138 2462
rect 3414 2458 3418 2462
rect 3814 2458 3818 2462
rect 3934 2448 3938 2452
rect 1150 2438 1154 2442
rect 1494 2428 1498 2432
rect 3814 2428 3818 2432
rect 2566 2418 2570 2422
rect 2918 2418 2922 2422
rect 4366 2418 4370 2422
rect 1558 2408 1562 2412
rect 1662 2408 1666 2412
rect 2566 2408 2570 2412
rect 2942 2408 2946 2412
rect 3238 2408 3242 2412
rect 3590 2408 3594 2412
rect 4014 2408 4018 2412
rect 4070 2408 4074 2412
rect 498 2403 502 2407
rect 506 2403 509 2407
rect 509 2403 510 2407
rect 1522 2403 1526 2407
rect 1530 2403 1533 2407
rect 1533 2403 1534 2407
rect 2546 2403 2550 2407
rect 2554 2403 2557 2407
rect 2557 2403 2558 2407
rect 3570 2403 3574 2407
rect 3578 2403 3581 2407
rect 3581 2403 3582 2407
rect 982 2398 986 2402
rect 2198 2398 2202 2402
rect 3262 2398 3266 2402
rect 1206 2388 1210 2392
rect 1358 2388 1362 2392
rect 2414 2388 2418 2392
rect 2806 2388 2810 2392
rect 3750 2388 3754 2392
rect 4214 2388 4218 2392
rect 4478 2388 4482 2392
rect 230 2378 234 2382
rect 1614 2378 1618 2382
rect 3366 2378 3370 2382
rect 1374 2368 1378 2372
rect 3374 2368 3378 2372
rect 4206 2368 4210 2372
rect 4350 2368 4354 2372
rect 4406 2368 4410 2372
rect 4510 2368 4514 2372
rect 4534 2368 4538 2372
rect 1414 2358 1418 2362
rect 2702 2358 2706 2362
rect 2814 2358 2818 2362
rect 3542 2358 3546 2362
rect 3950 2358 3954 2362
rect 3998 2358 4002 2362
rect 4142 2358 4146 2362
rect 2262 2348 2266 2352
rect 2582 2348 2586 2352
rect 2830 2348 2834 2352
rect 2974 2348 2978 2352
rect 2982 2348 2986 2352
rect 3398 2348 3402 2352
rect 3590 2348 3594 2352
rect 3862 2348 3866 2352
rect 4014 2348 4018 2352
rect 4270 2348 4274 2352
rect 4326 2348 4330 2352
rect 4574 2348 4578 2352
rect 926 2338 930 2342
rect 1278 2338 1282 2342
rect 2126 2338 2130 2342
rect 2206 2338 2210 2342
rect 2718 2338 2722 2342
rect 2758 2338 2762 2342
rect 3414 2338 3418 2342
rect 3430 2338 3434 2342
rect 3598 2338 3602 2342
rect 3974 2338 3978 2342
rect 4158 2338 4162 2342
rect 894 2328 898 2332
rect 950 2328 954 2332
rect 1726 2328 1730 2332
rect 2174 2328 2178 2332
rect 2294 2328 2298 2332
rect 2358 2328 2362 2332
rect 2462 2328 2466 2332
rect 2902 2328 2906 2332
rect 3366 2328 3370 2332
rect 3558 2328 3562 2332
rect 4310 2328 4314 2332
rect 4342 2328 4346 2332
rect 4566 2328 4570 2332
rect 1758 2318 1762 2322
rect 1918 2318 1922 2322
rect 2998 2318 3002 2322
rect 3406 2318 3410 2322
rect 214 2308 218 2312
rect 902 2308 906 2312
rect 2814 2308 2818 2312
rect 3078 2308 3082 2312
rect 3214 2308 3218 2312
rect 4310 2308 4314 2312
rect 4382 2308 4386 2312
rect 1002 2303 1006 2307
rect 1010 2303 1013 2307
rect 1013 2303 1014 2307
rect 2026 2303 2030 2307
rect 2034 2303 2037 2307
rect 2037 2303 2038 2307
rect 3050 2303 3054 2307
rect 3058 2303 3061 2307
rect 3061 2303 3062 2307
rect 4082 2303 4086 2307
rect 4090 2303 4093 2307
rect 4093 2303 4094 2307
rect 302 2298 306 2302
rect 1366 2298 1370 2302
rect 2630 2298 2634 2302
rect 2678 2298 2682 2302
rect 2734 2298 2738 2302
rect 3118 2298 3122 2302
rect 3838 2298 3842 2302
rect 4254 2298 4258 2302
rect 4518 2298 4522 2302
rect 1078 2288 1082 2292
rect 1646 2288 1650 2292
rect 2238 2288 2242 2292
rect 2270 2288 2274 2292
rect 2686 2288 2690 2292
rect 4126 2288 4130 2292
rect 4486 2288 4490 2292
rect 230 2278 234 2282
rect 1038 2278 1042 2282
rect 1086 2278 1090 2282
rect 1102 2278 1106 2282
rect 2574 2278 2578 2282
rect 2750 2278 2754 2282
rect 2774 2278 2778 2282
rect 2926 2278 2930 2282
rect 3438 2278 3442 2282
rect 3670 2278 3674 2282
rect 470 2268 474 2272
rect 774 2268 778 2272
rect 1078 2268 1082 2272
rect 1582 2268 1586 2272
rect 1926 2268 1930 2272
rect 2182 2268 2186 2272
rect 3862 2278 3866 2282
rect 2262 2268 2266 2272
rect 2390 2268 2394 2272
rect 2662 2268 2666 2272
rect 2694 2268 2698 2272
rect 2710 2268 2714 2272
rect 3166 2268 3170 2272
rect 3494 2268 3498 2272
rect 3758 2268 3762 2272
rect 4086 2268 4090 2272
rect 4326 2268 4330 2272
rect 1598 2258 1602 2262
rect 2326 2258 2330 2262
rect 2566 2258 2570 2262
rect 2942 2258 2946 2262
rect 3222 2258 3226 2262
rect 3470 2258 3474 2262
rect 4086 2258 4090 2262
rect 4134 2258 4138 2262
rect 4198 2258 4202 2262
rect 4374 2258 4378 2262
rect 4526 2258 4530 2262
rect 774 2248 778 2252
rect 2022 2248 2026 2252
rect 2566 2248 2570 2252
rect 2894 2248 2898 2252
rect 2902 2248 2906 2252
rect 3118 2248 3122 2252
rect 3374 2248 3378 2252
rect 4350 2248 4354 2252
rect 2262 2238 2266 2242
rect 2326 2238 2330 2242
rect 3222 2238 3226 2242
rect 3430 2238 3434 2242
rect 3478 2238 3482 2242
rect 4494 2238 4498 2242
rect 1862 2228 1866 2232
rect 2414 2228 2418 2232
rect 2806 2228 2810 2232
rect 3286 2228 3290 2232
rect 3838 2228 3842 2232
rect 4022 2228 4026 2232
rect 934 2218 938 2222
rect 2350 2218 2354 2222
rect 3390 2218 3394 2222
rect 1302 2208 1306 2212
rect 1606 2208 1610 2212
rect 2654 2208 2658 2212
rect 4086 2208 4090 2212
rect 498 2203 502 2207
rect 506 2203 509 2207
rect 509 2203 510 2207
rect 1522 2203 1526 2207
rect 1530 2203 1533 2207
rect 1533 2203 1534 2207
rect 2546 2203 2550 2207
rect 2554 2203 2557 2207
rect 2557 2203 2558 2207
rect 3570 2203 3574 2207
rect 3578 2203 3581 2207
rect 3581 2203 3582 2207
rect 1702 2198 1706 2202
rect 2310 2198 2314 2202
rect 2566 2198 2570 2202
rect 3710 2198 3714 2202
rect 4022 2198 4026 2202
rect 334 2188 338 2192
rect 1078 2188 1082 2192
rect 1134 2188 1138 2192
rect 1622 2188 1626 2192
rect 2430 2188 2434 2192
rect 2542 2188 2546 2192
rect 2678 2188 2682 2192
rect 3270 2188 3274 2192
rect 4134 2188 4138 2192
rect 4326 2188 4330 2192
rect 854 2178 858 2182
rect 1326 2178 1330 2182
rect 2102 2178 2106 2182
rect 3494 2178 3498 2182
rect 3782 2178 3786 2182
rect 4286 2178 4290 2182
rect 1430 2168 1434 2172
rect 3438 2168 3442 2172
rect 3750 2168 3754 2172
rect 1134 2158 1138 2162
rect 1406 2158 1410 2162
rect 2214 2158 2218 2162
rect 2582 2158 2586 2162
rect 2662 2158 2666 2162
rect 3038 2158 3042 2162
rect 3358 2158 3362 2162
rect 3510 2158 3514 2162
rect 3686 2158 3690 2162
rect 3766 2158 3770 2162
rect 4046 2158 4050 2162
rect 4206 2158 4210 2162
rect 454 2148 458 2152
rect 806 2148 810 2152
rect 1326 2148 1330 2152
rect 1334 2148 1338 2152
rect 2342 2148 2346 2152
rect 2398 2148 2402 2152
rect 2606 2148 2610 2152
rect 2678 2148 2682 2152
rect 2942 2148 2946 2152
rect 3030 2148 3034 2152
rect 3182 2148 3186 2152
rect 3230 2148 3234 2152
rect 3406 2148 3410 2152
rect 3790 2148 3794 2152
rect 3830 2148 3834 2152
rect 4126 2148 4130 2152
rect 4302 2148 4306 2152
rect 4430 2148 4434 2152
rect 846 2138 850 2142
rect 1510 2138 1514 2142
rect 1694 2138 1698 2142
rect 1734 2138 1738 2142
rect 1774 2138 1778 2142
rect 2206 2138 2210 2142
rect 2270 2138 2274 2142
rect 2454 2138 2458 2142
rect 2462 2138 2466 2142
rect 3166 2138 3170 2142
rect 3222 2138 3226 2142
rect 3246 2138 3250 2142
rect 3270 2138 3274 2142
rect 3550 2138 3554 2142
rect 3782 2138 3786 2142
rect 4502 2138 4506 2142
rect 1982 2128 1986 2132
rect 2238 2128 2242 2132
rect 2542 2128 2546 2132
rect 2974 2128 2978 2132
rect 3094 2128 3098 2132
rect 3102 2128 3106 2132
rect 3166 2128 3170 2132
rect 3646 2128 3650 2132
rect 3670 2128 3674 2132
rect 3862 2128 3866 2132
rect 1694 2118 1698 2122
rect 2046 2118 2050 2122
rect 2302 2118 2306 2122
rect 3086 2118 3090 2122
rect 3550 2118 3554 2122
rect 3838 2118 3842 2122
rect 3854 2118 3858 2122
rect 4254 2118 4258 2122
rect 4350 2118 4354 2122
rect 4398 2118 4402 2122
rect 4406 2118 4410 2122
rect 4454 2118 4458 2122
rect 974 2108 978 2112
rect 2014 2108 2018 2112
rect 3254 2108 3258 2112
rect 3326 2108 3330 2112
rect 3630 2108 3634 2112
rect 3870 2108 3874 2112
rect 1002 2103 1006 2107
rect 1010 2103 1013 2107
rect 1013 2103 1014 2107
rect 2026 2103 2030 2107
rect 2034 2103 2037 2107
rect 2037 2103 2038 2107
rect 3050 2103 3054 2107
rect 3058 2103 3061 2107
rect 3061 2103 3062 2107
rect 4082 2103 4086 2107
rect 4090 2103 4093 2107
rect 4093 2103 4094 2107
rect 990 2098 994 2102
rect 1542 2098 1546 2102
rect 2406 2098 2410 2102
rect 310 2088 314 2092
rect 966 2088 970 2092
rect 1070 2088 1074 2092
rect 2270 2088 2274 2092
rect 2662 2088 2666 2092
rect 3270 2088 3274 2092
rect 3382 2088 3386 2092
rect 4534 2088 4538 2092
rect 782 2078 786 2082
rect 1006 2078 1010 2082
rect 1078 2078 1082 2082
rect 1102 2078 1106 2082
rect 1598 2078 1602 2082
rect 1790 2078 1794 2082
rect 2710 2078 2714 2082
rect 2934 2078 2938 2082
rect 2950 2078 2954 2082
rect 4190 2078 4194 2082
rect 4262 2078 4266 2082
rect 4350 2078 4354 2082
rect 4486 2078 4490 2082
rect 278 2068 282 2072
rect 326 2068 330 2072
rect 862 2068 866 2072
rect 894 2068 898 2072
rect 1246 2068 1250 2072
rect 1566 2068 1570 2072
rect 1710 2068 1714 2072
rect 1926 2068 1930 2072
rect 2406 2068 2410 2072
rect 2582 2068 2586 2072
rect 2726 2068 2730 2072
rect 3750 2068 3754 2072
rect 3814 2068 3818 2072
rect 4246 2068 4250 2072
rect 4270 2068 4274 2072
rect 4574 2068 4578 2072
rect 766 2058 770 2062
rect 862 2058 866 2062
rect 870 2058 874 2062
rect 1262 2058 1266 2062
rect 1662 2058 1666 2062
rect 1782 2058 1786 2062
rect 2126 2058 2130 2062
rect 2134 2058 2138 2062
rect 2294 2058 2298 2062
rect 2406 2058 2410 2062
rect 2446 2058 2450 2062
rect 3070 2058 3074 2062
rect 3702 2058 3706 2062
rect 3774 2058 3778 2062
rect 4302 2058 4306 2062
rect 4318 2058 4322 2062
rect 4430 2058 4434 2062
rect 4478 2058 4482 2062
rect 4550 2058 4554 2062
rect 454 2048 458 2052
rect 470 2048 474 2052
rect 646 2048 650 2052
rect 806 2048 810 2052
rect 878 2048 882 2052
rect 1566 2048 1570 2052
rect 2158 2048 2162 2052
rect 2302 2048 2306 2052
rect 3374 2048 3378 2052
rect 3582 2048 3586 2052
rect 3758 2048 3762 2052
rect 3782 2048 3786 2052
rect 3806 2048 3810 2052
rect 3878 2048 3882 2052
rect 246 2038 250 2042
rect 1694 2038 1698 2042
rect 3814 2038 3818 2042
rect 1430 2028 1434 2032
rect 2006 2028 2010 2032
rect 2254 2028 2258 2032
rect 766 2018 770 2022
rect 1726 2018 1730 2022
rect 3358 2018 3362 2022
rect 3798 2018 3802 2022
rect 4046 2018 4050 2022
rect 478 2008 482 2012
rect 1510 2008 1514 2012
rect 1902 2008 1906 2012
rect 1918 2008 1922 2012
rect 2494 2008 2498 2012
rect 3150 2008 3154 2012
rect 3190 2008 3194 2012
rect 3750 2008 3754 2012
rect 3974 2008 3978 2012
rect 498 2003 502 2007
rect 506 2003 509 2007
rect 509 2003 510 2007
rect 1522 2003 1526 2007
rect 1530 2003 1533 2007
rect 1533 2003 1534 2007
rect 2546 2003 2550 2007
rect 2554 2003 2557 2007
rect 2557 2003 2558 2007
rect 3570 2003 3574 2007
rect 3578 2003 3581 2007
rect 3581 2003 3582 2007
rect 1438 1998 1442 2002
rect 1542 1998 1546 2002
rect 2254 1998 2258 2002
rect 2566 1998 2570 2002
rect 3686 1998 3690 2002
rect 4054 1998 4058 2002
rect 4398 1998 4402 2002
rect 1718 1988 1722 1992
rect 3182 1988 3186 1992
rect 3518 1988 3522 1992
rect 4246 1988 4250 1992
rect 478 1978 482 1982
rect 1542 1978 1546 1982
rect 1782 1978 1786 1982
rect 1974 1978 1978 1982
rect 2302 1978 2306 1982
rect 2350 1978 2354 1982
rect 2566 1978 2570 1982
rect 2670 1978 2674 1982
rect 4406 1978 4410 1982
rect 382 1968 386 1972
rect 926 1968 930 1972
rect 3022 1968 3026 1972
rect 3158 1968 3162 1972
rect 3358 1968 3362 1972
rect 3510 1968 3514 1972
rect 3678 1968 3682 1972
rect 3702 1968 3706 1972
rect 3726 1968 3730 1972
rect 318 1958 322 1962
rect 334 1958 338 1962
rect 550 1958 554 1962
rect 1718 1958 1722 1962
rect 1774 1958 1778 1962
rect 2430 1958 2434 1962
rect 2678 1958 2682 1962
rect 3038 1958 3042 1962
rect 3070 1958 3074 1962
rect 3822 1958 3826 1962
rect 3838 1958 3842 1962
rect 3958 1958 3962 1962
rect 3982 1958 3986 1962
rect 4166 1958 4170 1962
rect 4398 1958 4402 1962
rect 310 1948 314 1952
rect 1142 1948 1146 1952
rect 1270 1948 1274 1952
rect 1630 1948 1634 1952
rect 1742 1948 1746 1952
rect 2374 1948 2378 1952
rect 2526 1948 2530 1952
rect 2702 1948 2706 1952
rect 2942 1948 2946 1952
rect 3198 1948 3202 1952
rect 3710 1948 3714 1952
rect 3830 1948 3834 1952
rect 3894 1948 3898 1952
rect 4142 1948 4146 1952
rect 4198 1948 4202 1952
rect 4294 1948 4298 1952
rect 902 1938 906 1942
rect 926 1938 930 1942
rect 1910 1938 1914 1942
rect 2110 1938 2114 1942
rect 2646 1938 2650 1942
rect 2958 1938 2962 1942
rect 3158 1938 3162 1942
rect 3246 1938 3250 1942
rect 3430 1938 3434 1942
rect 3838 1938 3842 1942
rect 1126 1928 1130 1932
rect 1142 1928 1146 1932
rect 1294 1928 1298 1932
rect 1830 1928 1834 1932
rect 1838 1928 1842 1932
rect 2006 1928 2010 1932
rect 2190 1928 2194 1932
rect 2254 1928 2258 1932
rect 2726 1928 2730 1932
rect 2942 1928 2946 1932
rect 3846 1928 3850 1932
rect 4030 1928 4034 1932
rect 4038 1928 4042 1932
rect 4454 1928 4458 1932
rect 230 1918 234 1922
rect 1934 1918 1938 1922
rect 2150 1918 2154 1922
rect 4062 1918 4066 1922
rect 4262 1918 4266 1922
rect 4302 1918 4306 1922
rect 4566 1918 4570 1922
rect 550 1908 554 1912
rect 1246 1908 1250 1912
rect 1990 1908 1994 1912
rect 2238 1908 2242 1912
rect 2646 1908 2650 1912
rect 3630 1908 3634 1912
rect 3942 1908 3946 1912
rect 3966 1908 3970 1912
rect 4070 1908 4074 1912
rect 4518 1908 4522 1912
rect 1002 1903 1006 1907
rect 1010 1903 1013 1907
rect 1013 1903 1014 1907
rect 2026 1903 2030 1907
rect 2034 1903 2037 1907
rect 2037 1903 2038 1907
rect 3050 1903 3054 1907
rect 3058 1903 3061 1907
rect 3061 1903 3062 1907
rect 4082 1903 4086 1907
rect 4090 1903 4093 1907
rect 4093 1903 4094 1907
rect 1742 1898 1746 1902
rect 1798 1898 1802 1902
rect 4054 1898 4058 1902
rect 4342 1898 4346 1902
rect 1126 1888 1130 1892
rect 2246 1888 2250 1892
rect 3750 1888 3754 1892
rect 1382 1878 1386 1882
rect 1566 1878 1570 1882
rect 1774 1878 1778 1882
rect 1902 1878 1906 1882
rect 2334 1878 2338 1882
rect 2702 1878 2706 1882
rect 2750 1878 2754 1882
rect 2950 1878 2954 1882
rect 3046 1878 3050 1882
rect 3694 1878 3698 1882
rect 3958 1878 3962 1882
rect 4126 1878 4130 1882
rect 4254 1878 4258 1882
rect 214 1868 218 1872
rect 350 1868 354 1872
rect 1638 1868 1642 1872
rect 1990 1868 1994 1872
rect 2374 1868 2378 1872
rect 2622 1868 2626 1872
rect 2654 1868 2658 1872
rect 246 1858 250 1862
rect 1694 1858 1698 1862
rect 1742 1858 1746 1862
rect 1766 1858 1770 1862
rect 2838 1858 2842 1862
rect 2990 1858 2994 1862
rect 430 1848 434 1852
rect 1662 1848 1666 1852
rect 902 1838 906 1842
rect 2190 1848 2194 1852
rect 3158 1848 3162 1852
rect 3198 1848 3202 1852
rect 4286 1848 4290 1852
rect 2174 1838 2178 1842
rect 3030 1838 3034 1842
rect 3862 1838 3866 1842
rect 1734 1828 1738 1832
rect 1838 1828 1842 1832
rect 2270 1828 2274 1832
rect 2630 1828 2634 1832
rect 3494 1828 3498 1832
rect 4022 1828 4026 1832
rect 486 1818 490 1822
rect 2206 1818 2210 1822
rect 1502 1808 1506 1812
rect 3558 1808 3562 1812
rect 4518 1808 4522 1812
rect 498 1803 502 1807
rect 506 1803 509 1807
rect 509 1803 510 1807
rect 1522 1803 1526 1807
rect 1530 1803 1533 1807
rect 1533 1803 1534 1807
rect 550 1798 554 1802
rect 1190 1798 1194 1802
rect 1902 1798 1906 1802
rect 2546 1803 2550 1807
rect 2554 1803 2557 1807
rect 2557 1803 2558 1807
rect 3570 1803 3574 1807
rect 3578 1803 3581 1807
rect 3581 1803 3582 1807
rect 3150 1798 3154 1802
rect 3366 1798 3370 1802
rect 3390 1798 3394 1802
rect 4430 1798 4434 1802
rect 1206 1788 1210 1792
rect 1486 1788 1490 1792
rect 1766 1788 1770 1792
rect 2214 1788 2218 1792
rect 2518 1788 2522 1792
rect 3134 1788 3138 1792
rect 3974 1788 3978 1792
rect 574 1778 578 1782
rect 782 1778 786 1782
rect 1686 1778 1690 1782
rect 2694 1778 2698 1782
rect 2806 1778 2810 1782
rect 3814 1778 3818 1782
rect 4070 1778 4074 1782
rect 4478 1778 4482 1782
rect 310 1768 314 1772
rect 326 1768 330 1772
rect 1198 1768 1202 1772
rect 1694 1768 1698 1772
rect 1734 1768 1738 1772
rect 3350 1768 3354 1772
rect 1510 1758 1514 1762
rect 2222 1758 2226 1762
rect 2510 1758 2514 1762
rect 2694 1758 2698 1762
rect 2814 1758 2818 1762
rect 3166 1758 3170 1762
rect 3686 1758 3690 1762
rect 3774 1758 3778 1762
rect 4318 1758 4322 1762
rect 4374 1758 4378 1762
rect 1390 1748 1394 1752
rect 1542 1748 1546 1752
rect 2966 1748 2970 1752
rect 2990 1748 2994 1752
rect 3038 1748 3042 1752
rect 3190 1748 3194 1752
rect 3278 1748 3282 1752
rect 3566 1748 3570 1752
rect 3630 1748 3634 1752
rect 3982 1748 3986 1752
rect 3990 1748 3994 1752
rect 4182 1748 4186 1752
rect 4230 1748 4234 1752
rect 4350 1748 4354 1752
rect 4406 1748 4410 1752
rect 798 1738 802 1742
rect 1198 1738 1202 1742
rect 1262 1738 1266 1742
rect 2262 1738 2266 1742
rect 2462 1738 2466 1742
rect 2494 1738 2498 1742
rect 3198 1738 3202 1742
rect 3238 1738 3242 1742
rect 3294 1738 3298 1742
rect 3542 1738 3546 1742
rect 3918 1738 3922 1742
rect 4142 1738 4146 1742
rect 4254 1738 4258 1742
rect 4286 1738 4290 1742
rect 318 1728 322 1732
rect 350 1728 354 1732
rect 1102 1728 1106 1732
rect 1230 1728 1234 1732
rect 2278 1728 2282 1732
rect 2622 1728 2626 1732
rect 2646 1728 2650 1732
rect 2814 1728 2818 1732
rect 3510 1728 3514 1732
rect 3566 1728 3570 1732
rect 3958 1728 3962 1732
rect 4510 1728 4514 1732
rect 2326 1718 2330 1722
rect 2358 1718 2362 1722
rect 2830 1718 2834 1722
rect 3502 1718 3506 1722
rect 3838 1718 3842 1722
rect 4310 1718 4314 1722
rect 462 1708 466 1712
rect 1214 1708 1218 1712
rect 1974 1708 1978 1712
rect 2910 1708 2914 1712
rect 3022 1708 3026 1712
rect 3766 1708 3770 1712
rect 3974 1708 3978 1712
rect 1002 1703 1006 1707
rect 1010 1703 1013 1707
rect 1013 1703 1014 1707
rect 2026 1703 2030 1707
rect 2034 1703 2037 1707
rect 2037 1703 2038 1707
rect 3050 1703 3054 1707
rect 3058 1703 3061 1707
rect 3061 1703 3062 1707
rect 4082 1703 4086 1707
rect 4090 1703 4093 1707
rect 4093 1703 4094 1707
rect 654 1698 658 1702
rect 790 1698 794 1702
rect 1662 1698 1666 1702
rect 2054 1698 2058 1702
rect 2486 1698 2490 1702
rect 2982 1698 2986 1702
rect 3038 1698 3042 1702
rect 3166 1698 3170 1702
rect 3550 1698 3554 1702
rect 4182 1698 4186 1702
rect 4238 1698 4242 1702
rect 766 1688 770 1692
rect 1158 1688 1162 1692
rect 1230 1688 1234 1692
rect 1342 1688 1346 1692
rect 2438 1688 2442 1692
rect 2526 1688 2530 1692
rect 2630 1688 2634 1692
rect 2694 1688 2698 1692
rect 2726 1688 2730 1692
rect 2838 1688 2842 1692
rect 190 1678 194 1682
rect 1206 1678 1210 1682
rect 1302 1678 1306 1682
rect 1318 1678 1322 1682
rect 1446 1678 1450 1682
rect 1606 1678 1610 1682
rect 1974 1678 1978 1682
rect 2102 1678 2106 1682
rect 2782 1678 2786 1682
rect 2926 1678 2930 1682
rect 2934 1678 2938 1682
rect 3030 1678 3034 1682
rect 3110 1678 3114 1682
rect 3270 1678 3274 1682
rect 3414 1678 3418 1682
rect 3478 1678 3482 1682
rect 3494 1678 3498 1682
rect 3550 1678 3554 1682
rect 3710 1678 3714 1682
rect 4110 1678 4114 1682
rect 4366 1678 4370 1682
rect 4598 1678 4602 1682
rect 1238 1668 1242 1672
rect 1702 1668 1706 1672
rect 1902 1668 1906 1672
rect 2486 1668 2490 1672
rect 2670 1668 2674 1672
rect 2918 1668 2922 1672
rect 3182 1668 3186 1672
rect 3206 1668 3210 1672
rect 3358 1668 3362 1672
rect 3678 1668 3682 1672
rect 3702 1668 3706 1672
rect 3958 1668 3962 1672
rect 3966 1668 3970 1672
rect 4454 1668 4458 1672
rect 326 1658 330 1662
rect 934 1658 938 1662
rect 1158 1658 1162 1662
rect 1190 1658 1194 1662
rect 1630 1658 1634 1662
rect 1662 1658 1666 1662
rect 2246 1658 2250 1662
rect 2358 1658 2362 1662
rect 2822 1658 2826 1662
rect 2982 1658 2986 1662
rect 3102 1658 3106 1662
rect 3118 1658 3122 1662
rect 3390 1658 3394 1662
rect 3542 1658 3546 1662
rect 3766 1658 3770 1662
rect 4190 1658 4194 1662
rect 598 1648 602 1652
rect 1750 1648 1754 1652
rect 1950 1648 1954 1652
rect 2670 1648 2674 1652
rect 2966 1648 2970 1652
rect 3198 1648 3202 1652
rect 3838 1648 3842 1652
rect 4006 1648 4010 1652
rect 4182 1648 4186 1652
rect 4398 1648 4402 1652
rect 4526 1648 4530 1652
rect 3694 1638 3698 1642
rect 4246 1638 4250 1642
rect 4310 1638 4314 1642
rect 654 1628 658 1632
rect 2854 1628 2858 1632
rect 2862 1628 2866 1632
rect 3030 1628 3034 1632
rect 4254 1628 4258 1632
rect 198 1618 202 1622
rect 2070 1618 2074 1622
rect 2398 1618 2402 1622
rect 2630 1618 2634 1622
rect 3222 1618 3226 1622
rect 3454 1618 3458 1622
rect 1742 1608 1746 1612
rect 1886 1608 1890 1612
rect 2710 1608 2714 1612
rect 4142 1608 4146 1612
rect 4238 1608 4242 1612
rect 498 1603 502 1607
rect 506 1603 509 1607
rect 509 1603 510 1607
rect 1522 1603 1526 1607
rect 1530 1603 1533 1607
rect 1533 1603 1534 1607
rect 2546 1603 2550 1607
rect 2554 1603 2557 1607
rect 2557 1603 2558 1607
rect 3570 1603 3574 1607
rect 3578 1603 3581 1607
rect 3581 1603 3582 1607
rect 846 1598 850 1602
rect 2278 1598 2282 1602
rect 2502 1598 2506 1602
rect 2518 1598 2522 1602
rect 2766 1598 2770 1602
rect 2894 1598 2898 1602
rect 3030 1598 3034 1602
rect 4006 1598 4010 1602
rect 4238 1598 4242 1602
rect 430 1588 434 1592
rect 1750 1588 1754 1592
rect 1926 1588 1930 1592
rect 1990 1588 1994 1592
rect 3190 1588 3194 1592
rect 3510 1588 3514 1592
rect 4078 1588 4082 1592
rect 598 1578 602 1582
rect 774 1578 778 1582
rect 2710 1578 2714 1582
rect 3630 1578 3634 1582
rect 3718 1578 3722 1582
rect 4150 1578 4154 1582
rect 4278 1578 4282 1582
rect 1790 1568 1794 1572
rect 2662 1568 2666 1572
rect 2846 1568 2850 1572
rect 3070 1568 3074 1572
rect 3350 1568 3354 1572
rect 3686 1568 3690 1572
rect 4022 1568 4026 1572
rect 4230 1568 4234 1572
rect 4390 1568 4394 1572
rect 222 1558 226 1562
rect 1022 1558 1026 1562
rect 1054 1558 1058 1562
rect 1198 1558 1202 1562
rect 1870 1558 1874 1562
rect 2366 1558 2370 1562
rect 2734 1558 2738 1562
rect 2854 1558 2858 1562
rect 3286 1558 3290 1562
rect 4254 1558 4258 1562
rect 4262 1558 4266 1562
rect 158 1548 162 1552
rect 294 1548 298 1552
rect 518 1548 522 1552
rect 1038 1548 1042 1552
rect 1446 1548 1450 1552
rect 1454 1548 1458 1552
rect 2350 1548 2354 1552
rect 2550 1548 2554 1552
rect 2670 1548 2674 1552
rect 2742 1548 2746 1552
rect 2790 1548 2794 1552
rect 2870 1548 2874 1552
rect 2886 1548 2890 1552
rect 3190 1548 3194 1552
rect 3278 1548 3282 1552
rect 3302 1548 3306 1552
rect 3374 1548 3378 1552
rect 3398 1548 3402 1552
rect 3526 1548 3530 1552
rect 3614 1548 3618 1552
rect 3950 1548 3954 1552
rect 4062 1548 4066 1552
rect 4166 1548 4170 1552
rect 4342 1548 4346 1552
rect 4398 1548 4402 1552
rect 4510 1548 4514 1552
rect 1046 1538 1050 1542
rect 1726 1538 1730 1542
rect 1766 1538 1770 1542
rect 1846 1538 1850 1542
rect 1878 1538 1882 1542
rect 2270 1538 2274 1542
rect 2390 1538 2394 1542
rect 2622 1538 2626 1542
rect 2894 1538 2898 1542
rect 2910 1538 2914 1542
rect 2998 1538 3002 1542
rect 4102 1538 4106 1542
rect 4182 1538 4186 1542
rect 4230 1538 4234 1542
rect 4254 1538 4258 1542
rect 4302 1538 4306 1542
rect 1598 1528 1602 1532
rect 1894 1528 1898 1532
rect 2726 1528 2730 1532
rect 2902 1528 2906 1532
rect 3086 1528 3090 1532
rect 3134 1528 3138 1532
rect 3502 1528 3506 1532
rect 3998 1528 4002 1532
rect 4054 1528 4058 1532
rect 4302 1528 4306 1532
rect 4574 1528 4578 1532
rect 1246 1518 1250 1522
rect 2270 1518 2274 1522
rect 2694 1518 2698 1522
rect 3198 1518 3202 1522
rect 3942 1518 3946 1522
rect 4038 1518 4042 1522
rect 4166 1518 4170 1522
rect 4174 1518 4178 1522
rect 4278 1518 4282 1522
rect 326 1508 330 1512
rect 558 1508 562 1512
rect 1022 1508 1026 1512
rect 1694 1508 1698 1512
rect 1902 1508 1906 1512
rect 2046 1508 2050 1512
rect 2198 1508 2202 1512
rect 2214 1508 2218 1512
rect 2334 1508 2338 1512
rect 2502 1508 2506 1512
rect 3110 1508 3114 1512
rect 3334 1508 3338 1512
rect 3366 1508 3370 1512
rect 3414 1508 3418 1512
rect 4198 1508 4202 1512
rect 1002 1503 1006 1507
rect 1010 1503 1013 1507
rect 1013 1503 1014 1507
rect 2026 1503 2030 1507
rect 2034 1503 2037 1507
rect 2037 1503 2038 1507
rect 3050 1503 3054 1507
rect 3058 1503 3061 1507
rect 3061 1503 3062 1507
rect 4082 1503 4086 1507
rect 4090 1503 4093 1507
rect 4093 1503 4094 1507
rect 1350 1498 1354 1502
rect 1614 1498 1618 1502
rect 1918 1498 1922 1502
rect 2102 1498 2106 1502
rect 2398 1498 2402 1502
rect 2878 1498 2882 1502
rect 3734 1498 3738 1502
rect 4214 1498 4218 1502
rect 430 1488 434 1492
rect 566 1488 570 1492
rect 1622 1488 1626 1492
rect 1710 1488 1714 1492
rect 1774 1488 1778 1492
rect 2862 1488 2866 1492
rect 2870 1488 2874 1492
rect 4550 1488 4554 1492
rect 1166 1478 1170 1482
rect 1662 1478 1666 1482
rect 1702 1478 1706 1482
rect 1790 1478 1794 1482
rect 2390 1478 2394 1482
rect 2494 1478 2498 1482
rect 2742 1478 2746 1482
rect 2830 1478 2834 1482
rect 2846 1478 2850 1482
rect 2854 1478 2858 1482
rect 3870 1478 3874 1482
rect 4118 1478 4122 1482
rect 214 1468 218 1472
rect 438 1468 442 1472
rect 1310 1468 1314 1472
rect 1446 1468 1450 1472
rect 158 1458 162 1462
rect 574 1458 578 1462
rect 598 1458 602 1462
rect 790 1458 794 1462
rect 1262 1458 1266 1462
rect 1350 1458 1354 1462
rect 1622 1458 1626 1462
rect 1814 1458 1818 1462
rect 2342 1468 2346 1472
rect 2470 1468 2474 1472
rect 2590 1468 2594 1472
rect 3054 1468 3058 1472
rect 3086 1468 3090 1472
rect 3110 1468 3114 1472
rect 3206 1468 3210 1472
rect 3230 1468 3234 1472
rect 3646 1468 3650 1472
rect 3982 1468 3986 1472
rect 3990 1468 3994 1472
rect 4230 1468 4234 1472
rect 4382 1468 4386 1472
rect 4558 1468 4562 1472
rect 4574 1468 4578 1472
rect 2150 1458 2154 1462
rect 2390 1458 2394 1462
rect 2694 1458 2698 1462
rect 2710 1458 2714 1462
rect 2886 1458 2890 1462
rect 3118 1458 3122 1462
rect 3126 1458 3130 1462
rect 3278 1458 3282 1462
rect 3302 1458 3306 1462
rect 3350 1458 3354 1462
rect 3390 1458 3394 1462
rect 3606 1458 3610 1462
rect 3694 1458 3698 1462
rect 3742 1458 3746 1462
rect 3878 1458 3882 1462
rect 3974 1458 3978 1462
rect 4014 1458 4018 1462
rect 4030 1458 4034 1462
rect 4150 1458 4154 1462
rect 4238 1458 4242 1462
rect 4270 1458 4274 1462
rect 4318 1458 4322 1462
rect 4334 1458 4338 1462
rect 1990 1448 1994 1452
rect 2262 1448 2266 1452
rect 2486 1448 2490 1452
rect 2662 1448 2666 1452
rect 3078 1448 3082 1452
rect 3614 1448 3618 1452
rect 4134 1448 4138 1452
rect 4166 1448 4170 1452
rect 4406 1448 4410 1452
rect 550 1438 554 1442
rect 2190 1438 2194 1442
rect 2878 1438 2882 1442
rect 2966 1438 2970 1442
rect 3086 1438 3090 1442
rect 3998 1438 4002 1442
rect 4558 1438 4562 1442
rect 334 1428 338 1432
rect 942 1428 946 1432
rect 1286 1428 1290 1432
rect 1646 1428 1650 1432
rect 1878 1428 1882 1432
rect 3214 1428 3218 1432
rect 4062 1428 4066 1432
rect 4494 1428 4498 1432
rect 1318 1418 1322 1422
rect 1414 1418 1418 1422
rect 2358 1418 2362 1422
rect 3166 1418 3170 1422
rect 3782 1418 3786 1422
rect 4326 1418 4330 1422
rect 1414 1408 1418 1412
rect 1958 1408 1962 1412
rect 2438 1408 2442 1412
rect 2534 1408 2538 1412
rect 2846 1408 2850 1412
rect 3158 1408 3162 1412
rect 3206 1408 3210 1412
rect 3238 1408 3242 1412
rect 3518 1408 3522 1412
rect 4230 1408 4234 1412
rect 4478 1408 4482 1412
rect 498 1403 502 1407
rect 506 1403 509 1407
rect 509 1403 510 1407
rect 1522 1403 1526 1407
rect 1530 1403 1533 1407
rect 1533 1403 1534 1407
rect 2546 1403 2550 1407
rect 2554 1403 2557 1407
rect 2557 1403 2558 1407
rect 3570 1403 3574 1407
rect 3578 1403 3581 1407
rect 3581 1403 3582 1407
rect 2934 1398 2938 1402
rect 4158 1398 4162 1402
rect 4190 1398 4194 1402
rect 4254 1398 4258 1402
rect 262 1388 266 1392
rect 1510 1388 1514 1392
rect 2206 1388 2210 1392
rect 2638 1388 2642 1392
rect 2646 1388 2650 1392
rect 3166 1388 3170 1392
rect 3214 1388 3218 1392
rect 3486 1388 3490 1392
rect 4054 1388 4058 1392
rect 4174 1388 4178 1392
rect 4246 1388 4250 1392
rect 4302 1388 4306 1392
rect 1142 1378 1146 1382
rect 2478 1378 2482 1382
rect 2526 1378 2530 1382
rect 2726 1378 2730 1382
rect 2766 1378 2770 1382
rect 2862 1378 2866 1382
rect 2870 1378 2874 1382
rect 3086 1378 3090 1382
rect 3134 1378 3138 1382
rect 3278 1378 3282 1382
rect 3670 1378 3674 1382
rect 3910 1378 3914 1382
rect 4574 1378 4578 1382
rect 350 1368 354 1372
rect 902 1368 906 1372
rect 1462 1368 1466 1372
rect 1502 1368 1506 1372
rect 1726 1368 1730 1372
rect 1870 1368 1874 1372
rect 2630 1368 2634 1372
rect 2966 1368 2970 1372
rect 2974 1368 2978 1372
rect 3374 1368 3378 1372
rect 3614 1368 3618 1372
rect 3766 1368 3770 1372
rect 3870 1368 3874 1372
rect 4182 1368 4186 1372
rect 4294 1368 4298 1372
rect 4526 1368 4530 1372
rect 846 1358 850 1362
rect 1054 1358 1058 1362
rect 1366 1358 1370 1362
rect 1478 1358 1482 1362
rect 2286 1358 2290 1362
rect 2366 1358 2370 1362
rect 2382 1358 2386 1362
rect 2734 1358 2738 1362
rect 2742 1358 2746 1362
rect 2894 1358 2898 1362
rect 2942 1358 2946 1362
rect 3582 1358 3586 1362
rect 3894 1358 3898 1362
rect 4006 1358 4010 1362
rect 4014 1358 4018 1362
rect 766 1348 770 1352
rect 2358 1348 2362 1352
rect 2454 1348 2458 1352
rect 2510 1348 2514 1352
rect 2646 1348 2650 1352
rect 2902 1348 2906 1352
rect 3070 1348 3074 1352
rect 3190 1348 3194 1352
rect 3206 1348 3210 1352
rect 3462 1348 3466 1352
rect 3526 1348 3530 1352
rect 3598 1348 3602 1352
rect 4022 1348 4026 1352
rect 4238 1348 4242 1352
rect 4318 1348 4322 1352
rect 4502 1348 4506 1352
rect 4566 1348 4570 1352
rect 558 1338 562 1342
rect 1558 1338 1562 1342
rect 2134 1338 2138 1342
rect 2262 1338 2266 1342
rect 2934 1338 2938 1342
rect 2950 1338 2954 1342
rect 3038 1338 3042 1342
rect 3278 1338 3282 1342
rect 3334 1338 3338 1342
rect 3734 1338 3738 1342
rect 4030 1338 4034 1342
rect 4214 1338 4218 1342
rect 158 1328 162 1332
rect 566 1328 570 1332
rect 1230 1328 1234 1332
rect 1566 1328 1570 1332
rect 1582 1328 1586 1332
rect 1694 1328 1698 1332
rect 1966 1328 1970 1332
rect 2214 1328 2218 1332
rect 2454 1328 2458 1332
rect 2662 1328 2666 1332
rect 2838 1328 2842 1332
rect 2926 1328 2930 1332
rect 3006 1328 3010 1332
rect 3110 1328 3114 1332
rect 3126 1328 3130 1332
rect 3206 1328 3210 1332
rect 3222 1328 3226 1332
rect 3526 1328 3530 1332
rect 3598 1328 3602 1332
rect 3966 1328 3970 1332
rect 4342 1328 4346 1332
rect 750 1318 754 1322
rect 1886 1318 1890 1322
rect 2646 1318 2650 1322
rect 3174 1318 3178 1322
rect 3222 1318 3226 1322
rect 3278 1318 3282 1322
rect 3590 1318 3594 1322
rect 3966 1318 3970 1322
rect 4214 1318 4218 1322
rect 4230 1318 4234 1322
rect 262 1308 266 1312
rect 1086 1308 1090 1312
rect 1406 1308 1410 1312
rect 1702 1308 1706 1312
rect 2766 1308 2770 1312
rect 2830 1308 2834 1312
rect 2854 1308 2858 1312
rect 3078 1308 3082 1312
rect 3294 1308 3298 1312
rect 3502 1308 3506 1312
rect 3694 1308 3698 1312
rect 4142 1308 4146 1312
rect 4358 1308 4362 1312
rect 1002 1303 1006 1307
rect 1010 1303 1013 1307
rect 1013 1303 1014 1307
rect 2026 1303 2030 1307
rect 2034 1303 2037 1307
rect 2037 1303 2038 1307
rect 1222 1298 1226 1302
rect 3050 1303 3054 1307
rect 3058 1303 3061 1307
rect 3061 1303 3062 1307
rect 4082 1303 4086 1307
rect 4090 1303 4093 1307
rect 4093 1303 4094 1307
rect 2926 1298 2930 1302
rect 3094 1298 3098 1302
rect 3142 1298 3146 1302
rect 3246 1298 3250 1302
rect 3486 1298 3490 1302
rect 3518 1298 3522 1302
rect 3670 1298 3674 1302
rect 3686 1298 3690 1302
rect 3798 1298 3802 1302
rect 3910 1298 3914 1302
rect 4278 1298 4282 1302
rect 1678 1288 1682 1292
rect 2662 1288 2666 1292
rect 2678 1288 2682 1292
rect 2718 1288 2722 1292
rect 2750 1288 2754 1292
rect 2966 1288 2970 1292
rect 3478 1288 3482 1292
rect 3654 1288 3658 1292
rect 430 1278 434 1282
rect 1382 1278 1386 1282
rect 1414 1278 1418 1282
rect 1878 1278 1882 1282
rect 2246 1278 2250 1282
rect 2518 1278 2522 1282
rect 2838 1278 2842 1282
rect 3030 1278 3034 1282
rect 3590 1278 3594 1282
rect 3750 1278 3754 1282
rect 3878 1278 3882 1282
rect 3958 1278 3962 1282
rect 4014 1278 4018 1282
rect 4030 1278 4034 1282
rect 4590 1278 4594 1282
rect 230 1268 234 1272
rect 302 1268 306 1272
rect 902 1268 906 1272
rect 1174 1268 1178 1272
rect 1206 1268 1210 1272
rect 1454 1268 1458 1272
rect 2102 1268 2106 1272
rect 2390 1268 2394 1272
rect 2542 1268 2546 1272
rect 2614 1268 2618 1272
rect 2734 1268 2738 1272
rect 3230 1268 3234 1272
rect 3270 1268 3274 1272
rect 3310 1268 3314 1272
rect 3318 1268 3322 1272
rect 3622 1268 3626 1272
rect 4094 1268 4098 1272
rect 4174 1268 4178 1272
rect 446 1258 450 1262
rect 486 1258 490 1262
rect 542 1258 546 1262
rect 1158 1258 1162 1262
rect 1542 1258 1546 1262
rect 1662 1258 1666 1262
rect 1734 1258 1738 1262
rect 2094 1258 2098 1262
rect 2150 1258 2154 1262
rect 2318 1258 2322 1262
rect 2494 1258 2498 1262
rect 2510 1258 2514 1262
rect 2654 1258 2658 1262
rect 2798 1258 2802 1262
rect 2886 1258 2890 1262
rect 2902 1258 2906 1262
rect 2918 1258 2922 1262
rect 2974 1258 2978 1262
rect 3142 1258 3146 1262
rect 3398 1258 3402 1262
rect 3470 1258 3474 1262
rect 3478 1258 3482 1262
rect 3550 1258 3554 1262
rect 3678 1258 3682 1262
rect 3702 1258 3706 1262
rect 3886 1258 3890 1262
rect 3982 1258 3986 1262
rect 4254 1258 4258 1262
rect 4318 1258 4322 1262
rect 4358 1258 4362 1262
rect 4550 1258 4554 1262
rect 750 1248 754 1252
rect 1222 1248 1226 1252
rect 1366 1248 1370 1252
rect 1382 1248 1386 1252
rect 1646 1248 1650 1252
rect 2238 1248 2242 1252
rect 2310 1248 2314 1252
rect 2574 1248 2578 1252
rect 2582 1248 2586 1252
rect 2710 1248 2714 1252
rect 2774 1248 2778 1252
rect 2846 1248 2850 1252
rect 2862 1248 2866 1252
rect 2886 1248 2890 1252
rect 2926 1248 2930 1252
rect 3054 1248 3058 1252
rect 3070 1248 3074 1252
rect 3078 1248 3082 1252
rect 3110 1248 3114 1252
rect 3478 1248 3482 1252
rect 3502 1248 3506 1252
rect 3598 1248 3602 1252
rect 4062 1248 4066 1252
rect 4302 1248 4306 1252
rect 4510 1248 4514 1252
rect 1606 1238 1610 1242
rect 1910 1238 1914 1242
rect 2654 1238 2658 1242
rect 2838 1238 2842 1242
rect 3038 1238 3042 1242
rect 3958 1238 3962 1242
rect 4462 1238 4466 1242
rect 1246 1228 1250 1232
rect 1438 1228 1442 1232
rect 1838 1228 1842 1232
rect 2734 1228 2738 1232
rect 2886 1228 2890 1232
rect 3054 1228 3058 1232
rect 3254 1228 3258 1232
rect 3414 1228 3418 1232
rect 3422 1228 3426 1232
rect 3542 1228 3546 1232
rect 3646 1228 3650 1232
rect 4046 1228 4050 1232
rect 4206 1228 4210 1232
rect 4238 1228 4242 1232
rect 4374 1228 4378 1232
rect 1286 1218 1290 1222
rect 1798 1218 1802 1222
rect 2910 1218 2914 1222
rect 3510 1218 3514 1222
rect 3630 1218 3634 1222
rect 4022 1218 4026 1222
rect 1142 1208 1146 1212
rect 1294 1208 1298 1212
rect 1694 1208 1698 1212
rect 2110 1208 2114 1212
rect 2318 1208 2322 1212
rect 2710 1208 2714 1212
rect 3366 1208 3370 1212
rect 3646 1208 3650 1212
rect 3966 1208 3970 1212
rect 4062 1208 4066 1212
rect 4326 1208 4330 1212
rect 498 1203 502 1207
rect 506 1203 509 1207
rect 509 1203 510 1207
rect 1522 1203 1526 1207
rect 1530 1203 1533 1207
rect 1533 1203 1534 1207
rect 2546 1203 2550 1207
rect 2554 1203 2557 1207
rect 2557 1203 2558 1207
rect 3570 1203 3574 1207
rect 3578 1203 3581 1207
rect 3581 1203 3582 1207
rect 542 1198 546 1202
rect 2046 1198 2050 1202
rect 2262 1198 2266 1202
rect 2742 1198 2746 1202
rect 3014 1198 3018 1202
rect 3166 1198 3170 1202
rect 3214 1198 3218 1202
rect 3342 1198 3346 1202
rect 3358 1198 3362 1202
rect 3542 1198 3546 1202
rect 3614 1198 3618 1202
rect 3670 1198 3674 1202
rect 4142 1198 4146 1202
rect 406 1188 410 1192
rect 1198 1188 1202 1192
rect 1598 1188 1602 1192
rect 1990 1188 1994 1192
rect 2414 1188 2418 1192
rect 2798 1188 2802 1192
rect 2878 1188 2882 1192
rect 3206 1188 3210 1192
rect 3486 1188 3490 1192
rect 3654 1188 3658 1192
rect 3726 1188 3730 1192
rect 3742 1188 3746 1192
rect 4182 1188 4186 1192
rect 526 1178 530 1182
rect 2350 1178 2354 1182
rect 2622 1178 2626 1182
rect 3774 1178 3778 1182
rect 3998 1178 4002 1182
rect 4022 1178 4026 1182
rect 4158 1178 4162 1182
rect 4278 1178 4282 1182
rect 1182 1168 1186 1172
rect 1246 1168 1250 1172
rect 1606 1168 1610 1172
rect 1702 1168 1706 1172
rect 1902 1168 1906 1172
rect 1958 1168 1962 1172
rect 2742 1168 2746 1172
rect 2854 1168 2858 1172
rect 2878 1168 2882 1172
rect 2998 1168 3002 1172
rect 3014 1168 3018 1172
rect 3262 1168 3266 1172
rect 3926 1168 3930 1172
rect 4422 1168 4426 1172
rect 398 1158 402 1162
rect 454 1158 458 1162
rect 494 1158 498 1162
rect 654 1158 658 1162
rect 1262 1158 1266 1162
rect 1406 1158 1410 1162
rect 2126 1158 2130 1162
rect 2246 1158 2250 1162
rect 2422 1158 2426 1162
rect 2470 1158 2474 1162
rect 2934 1158 2938 1162
rect 3094 1158 3098 1162
rect 3110 1158 3114 1162
rect 3142 1158 3146 1162
rect 3182 1158 3186 1162
rect 3358 1158 3362 1162
rect 3438 1158 3442 1162
rect 3446 1158 3450 1162
rect 3486 1158 3490 1162
rect 3830 1158 3834 1162
rect 4014 1158 4018 1162
rect 4134 1158 4138 1162
rect 4206 1158 4210 1162
rect 4438 1158 4442 1162
rect 4486 1158 4490 1162
rect 4598 1158 4602 1162
rect 406 1148 410 1152
rect 790 1148 794 1152
rect 806 1148 810 1152
rect 1054 1148 1058 1152
rect 1222 1148 1226 1152
rect 1286 1148 1290 1152
rect 1486 1148 1490 1152
rect 1686 1148 1690 1152
rect 1742 1148 1746 1152
rect 1814 1148 1818 1152
rect 2350 1148 2354 1152
rect 2398 1148 2402 1152
rect 2430 1148 2434 1152
rect 2478 1148 2482 1152
rect 2606 1148 2610 1152
rect 2758 1148 2762 1152
rect 2766 1148 2770 1152
rect 2798 1148 2802 1152
rect 3006 1148 3010 1152
rect 3038 1148 3042 1152
rect 3110 1148 3114 1152
rect 3734 1148 3738 1152
rect 3966 1148 3970 1152
rect 4198 1148 4202 1152
rect 4262 1148 4266 1152
rect 4438 1148 4442 1152
rect 1942 1138 1946 1142
rect 2398 1138 2402 1142
rect 2430 1138 2434 1142
rect 2630 1138 2634 1142
rect 2662 1138 2666 1142
rect 3102 1138 3106 1142
rect 3134 1138 3138 1142
rect 3270 1138 3274 1142
rect 3286 1138 3290 1142
rect 3302 1138 3306 1142
rect 3326 1138 3330 1142
rect 3414 1138 3418 1142
rect 3790 1138 3794 1142
rect 3870 1138 3874 1142
rect 4126 1138 4130 1142
rect 326 1128 330 1132
rect 526 1128 530 1132
rect 942 1128 946 1132
rect 1086 1128 1090 1132
rect 1286 1128 1290 1132
rect 1406 1128 1410 1132
rect 1454 1128 1458 1132
rect 1990 1128 1994 1132
rect 2046 1128 2050 1132
rect 2238 1128 2242 1132
rect 2574 1128 2578 1132
rect 2590 1128 2594 1132
rect 2926 1128 2930 1132
rect 3318 1128 3322 1132
rect 3550 1128 3554 1132
rect 3558 1128 3562 1132
rect 3606 1128 3610 1132
rect 3630 1128 3634 1132
rect 3766 1128 3770 1132
rect 4070 1128 4074 1132
rect 4158 1128 4162 1132
rect 4238 1128 4242 1132
rect 4318 1128 4322 1132
rect 4478 1128 4482 1132
rect 1870 1118 1874 1122
rect 2110 1118 2114 1122
rect 2702 1118 2706 1122
rect 2934 1118 2938 1122
rect 2982 1118 2986 1122
rect 2998 1118 3002 1122
rect 3166 1118 3170 1122
rect 3206 1118 3210 1122
rect 3278 1118 3282 1122
rect 3526 1118 3530 1122
rect 3758 1118 3762 1122
rect 4342 1118 4346 1122
rect 310 1108 314 1112
rect 1190 1108 1194 1112
rect 1614 1108 1618 1112
rect 1814 1108 1818 1112
rect 2006 1108 2010 1112
rect 2446 1108 2450 1112
rect 2718 1108 2722 1112
rect 3038 1108 3042 1112
rect 3110 1108 3114 1112
rect 3270 1108 3274 1112
rect 3454 1108 3458 1112
rect 3774 1108 3778 1112
rect 4030 1108 4034 1112
rect 4126 1108 4130 1112
rect 4214 1108 4218 1112
rect 4422 1108 4426 1112
rect 1002 1103 1006 1107
rect 1010 1103 1013 1107
rect 1013 1103 1014 1107
rect 678 1098 682 1102
rect 1198 1098 1202 1102
rect 1358 1098 1362 1102
rect 1366 1098 1370 1102
rect 2026 1103 2030 1107
rect 2034 1103 2037 1107
rect 2037 1103 2038 1107
rect 3050 1103 3054 1107
rect 3058 1103 3061 1107
rect 3061 1103 3062 1107
rect 4082 1103 4086 1107
rect 4090 1103 4093 1107
rect 4093 1103 4094 1107
rect 1486 1098 1490 1102
rect 1998 1098 2002 1102
rect 2326 1098 2330 1102
rect 2358 1098 2362 1102
rect 2470 1098 2474 1102
rect 2622 1098 2626 1102
rect 2830 1098 2834 1102
rect 3070 1098 3074 1102
rect 3542 1098 3546 1102
rect 3846 1098 3850 1102
rect 3854 1098 3858 1102
rect 4414 1098 4418 1102
rect 1238 1088 1242 1092
rect 1510 1088 1514 1092
rect 2150 1088 2154 1092
rect 2678 1088 2682 1092
rect 2902 1088 2906 1092
rect 2942 1088 2946 1092
rect 3630 1088 3634 1092
rect 3766 1088 3770 1092
rect 3782 1088 3786 1092
rect 4150 1088 4154 1092
rect 4190 1088 4194 1092
rect 4358 1088 4362 1092
rect 918 1078 922 1082
rect 1446 1078 1450 1082
rect 2174 1078 2178 1082
rect 2206 1078 2210 1082
rect 2270 1078 2274 1082
rect 2494 1078 2498 1082
rect 2830 1078 2834 1082
rect 3262 1078 3266 1082
rect 3310 1078 3314 1082
rect 3518 1078 3522 1082
rect 3806 1078 3810 1082
rect 3982 1078 3986 1082
rect 4214 1078 4218 1082
rect 4294 1078 4298 1082
rect 4342 1078 4346 1082
rect 4478 1078 4482 1082
rect 4486 1078 4490 1082
rect 302 1068 306 1072
rect 1230 1068 1234 1072
rect 1454 1068 1458 1072
rect 1718 1068 1722 1072
rect 1854 1068 1858 1072
rect 2046 1068 2050 1072
rect 2070 1068 2074 1072
rect 2102 1068 2106 1072
rect 2302 1068 2306 1072
rect 2446 1068 2450 1072
rect 2590 1068 2594 1072
rect 2654 1068 2658 1072
rect 2718 1068 2722 1072
rect 2750 1068 2754 1072
rect 2814 1068 2818 1072
rect 2958 1068 2962 1072
rect 2998 1068 3002 1072
rect 3014 1068 3018 1072
rect 3030 1068 3034 1072
rect 3294 1068 3298 1072
rect 3326 1068 3330 1072
rect 3350 1068 3354 1072
rect 3430 1068 3434 1072
rect 3470 1068 3474 1072
rect 3502 1068 3506 1072
rect 3534 1068 3538 1072
rect 3574 1068 3578 1072
rect 3606 1068 3610 1072
rect 3638 1068 3642 1072
rect 3670 1068 3674 1072
rect 3734 1068 3738 1072
rect 3782 1068 3786 1072
rect 4038 1068 4042 1072
rect 4198 1068 4202 1072
rect 4238 1068 4242 1072
rect 4454 1068 4458 1072
rect 230 1058 234 1062
rect 366 1058 370 1062
rect 430 1058 434 1062
rect 934 1058 938 1062
rect 1302 1058 1306 1062
rect 1486 1058 1490 1062
rect 1950 1058 1954 1062
rect 1966 1058 1970 1062
rect 1990 1058 1994 1062
rect 2094 1058 2098 1062
rect 2110 1058 2114 1062
rect 2334 1058 2338 1062
rect 2438 1058 2442 1062
rect 2454 1058 2458 1062
rect 2614 1058 2618 1062
rect 2726 1058 2730 1062
rect 2798 1058 2802 1062
rect 3006 1058 3010 1062
rect 3038 1058 3042 1062
rect 3118 1058 3122 1062
rect 3190 1058 3194 1062
rect 3238 1058 3242 1062
rect 3590 1058 3594 1062
rect 3966 1058 3970 1062
rect 4046 1058 4050 1062
rect 4454 1058 4458 1062
rect 350 1048 354 1052
rect 1774 1048 1778 1052
rect 1998 1048 2002 1052
rect 2086 1048 2090 1052
rect 2654 1048 2658 1052
rect 2694 1048 2698 1052
rect 2766 1048 2770 1052
rect 3118 1048 3122 1052
rect 3158 1048 3162 1052
rect 3358 1048 3362 1052
rect 3390 1048 3394 1052
rect 3454 1048 3458 1052
rect 3502 1048 3506 1052
rect 3662 1048 3666 1052
rect 3702 1048 3706 1052
rect 3774 1048 3778 1052
rect 3822 1048 3826 1052
rect 3846 1048 3850 1052
rect 4118 1048 4122 1052
rect 4334 1048 4338 1052
rect 4398 1048 4402 1052
rect 966 1038 970 1042
rect 2166 1038 2170 1042
rect 2942 1038 2946 1042
rect 2998 1038 3002 1042
rect 3190 1038 3194 1042
rect 3222 1038 3226 1042
rect 3238 1038 3242 1042
rect 3486 1038 3490 1042
rect 3694 1038 3698 1042
rect 3742 1038 3746 1042
rect 3918 1038 3922 1042
rect 4094 1038 4098 1042
rect 4438 1038 4442 1042
rect 4558 1038 4562 1042
rect 1054 1028 1058 1032
rect 1694 1028 1698 1032
rect 2086 1028 2090 1032
rect 2206 1028 2210 1032
rect 3134 1028 3138 1032
rect 4006 1028 4010 1032
rect 4014 1028 4018 1032
rect 4438 1028 4442 1032
rect 2646 1018 2650 1022
rect 2878 1018 2882 1022
rect 3278 1018 3282 1022
rect 3478 1018 3482 1022
rect 3766 1018 3770 1022
rect 4022 1018 4026 1022
rect 4326 1018 4330 1022
rect 4382 1018 4386 1022
rect 4566 1018 4570 1022
rect 2318 1008 2322 1012
rect 3126 1008 3130 1012
rect 3838 1008 3842 1012
rect 3862 1008 3866 1012
rect 4190 1008 4194 1012
rect 4390 1008 4394 1012
rect 498 1003 502 1007
rect 506 1003 509 1007
rect 509 1003 510 1007
rect 1522 1003 1526 1007
rect 1530 1003 1533 1007
rect 1533 1003 1534 1007
rect 2546 1003 2550 1007
rect 2554 1003 2557 1007
rect 2557 1003 2558 1007
rect 3570 1003 3574 1007
rect 3578 1003 3581 1007
rect 3581 1003 3582 1007
rect 222 998 226 1002
rect 1134 998 1138 1002
rect 1166 998 1170 1002
rect 1862 998 1866 1002
rect 1894 998 1898 1002
rect 2006 998 2010 1002
rect 2638 998 2642 1002
rect 2742 998 2746 1002
rect 2942 998 2946 1002
rect 2974 998 2978 1002
rect 2998 998 3002 1002
rect 3230 998 3234 1002
rect 3382 998 3386 1002
rect 4166 998 4170 1002
rect 4598 998 4602 1002
rect 2054 988 2058 992
rect 2174 988 2178 992
rect 3334 988 3338 992
rect 3390 988 3394 992
rect 4390 988 4394 992
rect 4406 988 4410 992
rect 1366 978 1370 982
rect 1742 978 1746 982
rect 2030 978 2034 982
rect 2478 978 2482 982
rect 2502 978 2506 982
rect 2782 978 2786 982
rect 3254 978 3258 982
rect 3334 978 3338 982
rect 3550 978 3554 982
rect 1758 968 1762 972
rect 1878 968 1882 972
rect 1934 968 1938 972
rect 2142 968 2146 972
rect 2974 968 2978 972
rect 3182 968 3186 972
rect 3262 968 3266 972
rect 3390 968 3394 972
rect 3430 968 3434 972
rect 3574 968 3578 972
rect 3686 968 3690 972
rect 310 958 314 962
rect 1014 958 1018 962
rect 1070 958 1074 962
rect 1198 958 1202 962
rect 1878 958 1882 962
rect 1894 958 1898 962
rect 2014 958 2018 962
rect 2366 958 2370 962
rect 2406 958 2410 962
rect 2606 958 2610 962
rect 2622 958 2626 962
rect 4110 968 4114 972
rect 4414 968 4418 972
rect 3078 958 3082 962
rect 3086 958 3090 962
rect 3358 958 3362 962
rect 3406 958 3410 962
rect 3670 958 3674 962
rect 3798 958 3802 962
rect 3806 958 3810 962
rect 3870 958 3874 962
rect 3886 958 3890 962
rect 4270 958 4274 962
rect 4366 958 4370 962
rect 4486 958 4490 962
rect 366 948 370 952
rect 1190 948 1194 952
rect 1222 948 1226 952
rect 1486 948 1490 952
rect 1686 948 1690 952
rect 2198 948 2202 952
rect 2414 948 2418 952
rect 2518 948 2522 952
rect 2542 948 2546 952
rect 2598 948 2602 952
rect 2790 948 2794 952
rect 2806 948 2810 952
rect 2894 948 2898 952
rect 2974 948 2978 952
rect 3006 948 3010 952
rect 3206 948 3210 952
rect 3222 948 3226 952
rect 3358 948 3362 952
rect 3566 948 3570 952
rect 3726 948 3730 952
rect 3766 948 3770 952
rect 3782 948 3786 952
rect 3830 948 3834 952
rect 3982 948 3986 952
rect 3990 948 3994 952
rect 4086 948 4090 952
rect 4174 948 4178 952
rect 4198 948 4202 952
rect 4230 948 4234 952
rect 4318 948 4322 952
rect 4454 948 4458 952
rect 4550 948 4554 952
rect 318 938 322 942
rect 982 938 986 942
rect 1078 938 1082 942
rect 1606 938 1610 942
rect 1782 938 1786 942
rect 1982 938 1986 942
rect 2158 938 2162 942
rect 2270 938 2274 942
rect 2398 938 2402 942
rect 2806 938 2810 942
rect 2862 938 2866 942
rect 2910 938 2914 942
rect 2926 938 2930 942
rect 2958 938 2962 942
rect 3046 938 3050 942
rect 3166 938 3170 942
rect 3238 938 3242 942
rect 3318 938 3322 942
rect 3350 938 3354 942
rect 3502 938 3506 942
rect 3550 938 3554 942
rect 3694 938 3698 942
rect 4030 938 4034 942
rect 4102 938 4106 942
rect 4110 938 4114 942
rect 4558 938 4562 942
rect 1158 928 1162 932
rect 1174 928 1178 932
rect 1374 928 1378 932
rect 1566 928 1570 932
rect 1814 928 1818 932
rect 1854 928 1858 932
rect 1926 928 1930 932
rect 2070 928 2074 932
rect 2086 928 2090 932
rect 2158 928 2162 932
rect 2446 928 2450 932
rect 2518 928 2522 932
rect 2590 928 2594 932
rect 2670 928 2674 932
rect 2702 928 2706 932
rect 2718 928 2722 932
rect 2854 928 2858 932
rect 3094 928 3098 932
rect 3262 928 3266 932
rect 3398 928 3402 932
rect 3430 928 3434 932
rect 3438 928 3442 932
rect 3470 928 3474 932
rect 3614 928 3618 932
rect 3630 928 3634 932
rect 3670 928 3674 932
rect 3710 928 3714 932
rect 3854 928 3858 932
rect 3886 928 3890 932
rect 4054 928 4058 932
rect 4414 928 4418 932
rect 4542 928 4546 932
rect 1294 918 1298 922
rect 1478 918 1482 922
rect 1678 918 1682 922
rect 1726 918 1730 922
rect 1958 918 1962 922
rect 2486 918 2490 922
rect 2630 918 2634 922
rect 2774 918 2778 922
rect 2830 918 2834 922
rect 2990 918 2994 922
rect 3006 918 3010 922
rect 3094 918 3098 922
rect 3110 918 3114 922
rect 3374 918 3378 922
rect 3622 918 3626 922
rect 3742 918 3746 922
rect 3766 918 3770 922
rect 4030 918 4034 922
rect 4038 918 4042 922
rect 4310 918 4314 922
rect 4534 918 4538 922
rect 1174 908 1178 912
rect 1590 908 1594 912
rect 1638 908 1642 912
rect 1686 908 1690 912
rect 1942 908 1946 912
rect 2766 908 2770 912
rect 3966 908 3970 912
rect 4182 908 4186 912
rect 1002 903 1006 907
rect 1010 903 1013 907
rect 1013 903 1014 907
rect 2026 903 2030 907
rect 2034 903 2037 907
rect 2037 903 2038 907
rect 1630 898 1634 902
rect 3050 903 3054 907
rect 3058 903 3061 907
rect 3061 903 3062 907
rect 4082 903 4086 907
rect 4090 903 4093 907
rect 4093 903 4094 907
rect 2406 898 2410 902
rect 1158 888 1162 892
rect 1190 888 1194 892
rect 1462 888 1466 892
rect 1478 888 1482 892
rect 1638 888 1642 892
rect 3222 898 3226 902
rect 3638 898 3642 902
rect 3790 898 3794 902
rect 4238 898 4242 902
rect 4526 898 4530 902
rect 2118 888 2122 892
rect 2302 888 2306 892
rect 2694 888 2698 892
rect 2758 888 2762 892
rect 3070 888 3074 892
rect 3134 888 3138 892
rect 3270 888 3274 892
rect 3446 888 3450 892
rect 3518 888 3522 892
rect 3542 888 3546 892
rect 3662 888 3666 892
rect 1614 878 1618 882
rect 1678 878 1682 882
rect 1758 878 1762 882
rect 1862 878 1866 882
rect 2126 878 2130 882
rect 2230 878 2234 882
rect 3350 878 3354 882
rect 3382 878 3386 882
rect 4278 888 4282 892
rect 3526 878 3530 882
rect 3726 878 3730 882
rect 3926 878 3930 882
rect 3934 878 3938 882
rect 4206 878 4210 882
rect 934 868 938 872
rect 1126 868 1130 872
rect 1198 868 1202 872
rect 1214 868 1218 872
rect 4486 878 4490 882
rect 1374 868 1378 872
rect 1478 868 1482 872
rect 1614 868 1618 872
rect 1694 868 1698 872
rect 558 858 562 862
rect 2150 868 2154 872
rect 2318 868 2322 872
rect 2342 868 2346 872
rect 2382 868 2386 872
rect 2454 868 2458 872
rect 2470 868 2474 872
rect 2502 868 2506 872
rect 2726 868 2730 872
rect 2958 868 2962 872
rect 2974 868 2978 872
rect 3014 868 3018 872
rect 3030 868 3034 872
rect 3046 868 3050 872
rect 3110 868 3114 872
rect 3142 868 3146 872
rect 3166 868 3170 872
rect 3206 868 3210 872
rect 3254 868 3258 872
rect 3302 868 3306 872
rect 3790 868 3794 872
rect 3870 868 3874 872
rect 4438 868 4442 872
rect 974 858 978 862
rect 1326 858 1330 862
rect 1742 858 1746 862
rect 1790 858 1794 862
rect 1886 858 1890 862
rect 2110 858 2114 862
rect 2126 858 2130 862
rect 2166 858 2170 862
rect 2726 858 2730 862
rect 2742 858 2746 862
rect 2766 858 2770 862
rect 2846 858 2850 862
rect 2854 858 2858 862
rect 2878 858 2882 862
rect 3150 858 3154 862
rect 3214 858 3218 862
rect 3582 858 3586 862
rect 3782 858 3786 862
rect 4070 858 4074 862
rect 4198 858 4202 862
rect 4262 858 4266 862
rect 4286 858 4290 862
rect 4294 858 4298 862
rect 4318 858 4322 862
rect 4422 858 4426 862
rect 4510 858 4514 862
rect 1182 848 1186 852
rect 1278 848 1282 852
rect 1334 848 1338 852
rect 1414 848 1418 852
rect 2014 848 2018 852
rect 2230 848 2234 852
rect 2694 848 2698 852
rect 2862 848 2866 852
rect 3062 848 3066 852
rect 3110 848 3114 852
rect 3350 848 3354 852
rect 3390 848 3394 852
rect 3398 848 3402 852
rect 3646 848 3650 852
rect 3846 848 3850 852
rect 3910 848 3914 852
rect 3942 848 3946 852
rect 3966 848 3970 852
rect 4158 848 4162 852
rect 4230 848 4234 852
rect 4286 848 4290 852
rect 4334 848 4338 852
rect 4590 848 4594 852
rect 222 838 226 842
rect 558 838 562 842
rect 1214 838 1218 842
rect 1590 838 1594 842
rect 1814 838 1818 842
rect 2142 838 2146 842
rect 2334 838 2338 842
rect 2478 838 2482 842
rect 3198 838 3202 842
rect 3310 838 3314 842
rect 3422 838 3426 842
rect 3702 838 3706 842
rect 3814 838 3818 842
rect 3830 838 3834 842
rect 4006 838 4010 842
rect 4030 838 4034 842
rect 4142 838 4146 842
rect 4454 838 4458 842
rect 1982 828 1986 832
rect 2062 828 2066 832
rect 2510 828 2514 832
rect 2958 828 2962 832
rect 3406 828 3410 832
rect 3454 828 3458 832
rect 3542 828 3546 832
rect 4214 828 4218 832
rect 4366 828 4370 832
rect 3422 818 3426 822
rect 3510 818 3514 822
rect 3694 818 3698 822
rect 4182 818 4186 822
rect 4350 818 4354 822
rect 2510 808 2514 812
rect 2710 808 2714 812
rect 2934 808 2938 812
rect 3158 808 3162 812
rect 3478 808 3482 812
rect 3518 808 3522 812
rect 3630 808 3634 812
rect 3702 808 3706 812
rect 3822 808 3826 812
rect 3830 808 3834 812
rect 498 803 502 807
rect 506 803 509 807
rect 509 803 510 807
rect 1522 803 1526 807
rect 1530 803 1533 807
rect 1533 803 1534 807
rect 2546 803 2550 807
rect 2554 803 2557 807
rect 2557 803 2558 807
rect 3570 803 3574 807
rect 3578 803 3581 807
rect 3581 803 3582 807
rect 582 798 586 802
rect 1878 798 1882 802
rect 2054 798 2058 802
rect 2566 798 2570 802
rect 3166 798 3170 802
rect 3230 798 3234 802
rect 3638 798 3642 802
rect 3830 798 3834 802
rect 3838 798 3842 802
rect 2294 788 2298 792
rect 2766 788 2770 792
rect 2822 788 2826 792
rect 2934 788 2938 792
rect 2982 788 2986 792
rect 3822 788 3826 792
rect 3950 788 3954 792
rect 3982 788 3986 792
rect 4118 788 4122 792
rect 4126 788 4130 792
rect 4302 788 4306 792
rect 310 778 314 782
rect 678 778 682 782
rect 2166 778 2170 782
rect 2534 778 2538 782
rect 2654 778 2658 782
rect 4206 778 4210 782
rect 1550 768 1554 772
rect 1630 768 1634 772
rect 2566 768 2570 772
rect 2590 768 2594 772
rect 2846 768 2850 772
rect 2926 768 2930 772
rect 3246 768 3250 772
rect 3502 768 3506 772
rect 4206 768 4210 772
rect 310 758 314 762
rect 366 758 370 762
rect 766 758 770 762
rect 1822 758 1826 762
rect 2358 758 2362 762
rect 2614 758 2618 762
rect 2638 758 2642 762
rect 2726 758 2730 762
rect 2966 758 2970 762
rect 2974 758 2978 762
rect 3214 758 3218 762
rect 3254 758 3258 762
rect 3398 758 3402 762
rect 3414 758 3418 762
rect 3438 758 3442 762
rect 3502 758 3506 762
rect 3718 758 3722 762
rect 3774 758 3778 762
rect 3830 758 3834 762
rect 4006 758 4010 762
rect 582 748 586 752
rect 1566 748 1570 752
rect 1598 748 1602 752
rect 1846 748 1850 752
rect 1878 748 1882 752
rect 2126 748 2130 752
rect 2198 748 2202 752
rect 2270 748 2274 752
rect 2438 748 2442 752
rect 2486 748 2490 752
rect 2526 748 2530 752
rect 2734 748 2738 752
rect 2790 748 2794 752
rect 2934 748 2938 752
rect 3198 748 3202 752
rect 3278 748 3282 752
rect 3294 748 3298 752
rect 3366 748 3370 752
rect 3374 748 3378 752
rect 3438 748 3442 752
rect 3462 748 3466 752
rect 3606 748 3610 752
rect 3614 748 3618 752
rect 3702 748 3706 752
rect 4014 748 4018 752
rect 4110 748 4114 752
rect 4158 748 4162 752
rect 4438 748 4442 752
rect 158 738 162 742
rect 198 738 202 742
rect 766 738 770 742
rect 1150 738 1154 742
rect 1254 738 1258 742
rect 1606 738 1610 742
rect 1774 738 1778 742
rect 2334 738 2338 742
rect 2414 738 2418 742
rect 2662 738 2666 742
rect 2798 738 2802 742
rect 2862 738 2866 742
rect 2886 738 2890 742
rect 2942 738 2946 742
rect 3430 738 3434 742
rect 3558 738 3562 742
rect 3574 738 3578 742
rect 3782 738 3786 742
rect 4022 738 4026 742
rect 4030 738 4034 742
rect 4070 738 4074 742
rect 4214 738 4218 742
rect 4262 738 4266 742
rect 4406 738 4410 742
rect 1622 728 1626 732
rect 2398 728 2402 732
rect 2694 728 2698 732
rect 2998 728 3002 732
rect 3038 728 3042 732
rect 3118 728 3122 732
rect 3462 728 3466 732
rect 3918 728 3922 732
rect 4054 728 4058 732
rect 4134 728 4138 732
rect 4358 728 4362 732
rect 4374 728 4378 732
rect 414 718 418 722
rect 430 718 434 722
rect 1294 718 1298 722
rect 1398 718 1402 722
rect 2182 718 2186 722
rect 2606 718 2610 722
rect 2622 718 2626 722
rect 2806 718 2810 722
rect 2934 718 2938 722
rect 3334 718 3338 722
rect 3478 718 3482 722
rect 3822 718 3826 722
rect 3854 718 3858 722
rect 3894 718 3898 722
rect 4342 718 4346 722
rect 2006 708 2010 712
rect 2414 708 2418 712
rect 3038 708 3042 712
rect 3134 708 3138 712
rect 3238 708 3242 712
rect 3262 708 3266 712
rect 3502 708 3506 712
rect 3606 708 3610 712
rect 3878 708 3882 712
rect 4502 708 4506 712
rect 1002 703 1006 707
rect 1010 703 1013 707
rect 1013 703 1014 707
rect 2026 703 2030 707
rect 2034 703 2037 707
rect 2037 703 2038 707
rect 3050 703 3054 707
rect 3058 703 3061 707
rect 3061 703 3062 707
rect 4082 703 4086 707
rect 4090 703 4093 707
rect 4093 703 4094 707
rect 1334 698 1338 702
rect 2574 698 2578 702
rect 2606 698 2610 702
rect 2838 698 2842 702
rect 3134 698 3138 702
rect 3294 698 3298 702
rect 3806 698 3810 702
rect 4422 698 4426 702
rect 1822 688 1826 692
rect 2030 688 2034 692
rect 2038 688 2042 692
rect 2622 688 2626 692
rect 2702 688 2706 692
rect 2774 688 2778 692
rect 2918 688 2922 692
rect 3750 688 3754 692
rect 3758 688 3762 692
rect 3894 688 3898 692
rect 3902 688 3906 692
rect 446 678 450 682
rect 526 678 530 682
rect 558 678 562 682
rect 278 668 282 672
rect 790 668 794 672
rect 1302 678 1306 682
rect 1646 678 1650 682
rect 2678 678 2682 682
rect 2718 678 2722 682
rect 2998 678 3002 682
rect 3070 678 3074 682
rect 3174 678 3178 682
rect 3598 678 3602 682
rect 3654 678 3658 682
rect 3726 678 3730 682
rect 4558 678 4562 682
rect 1462 668 1466 672
rect 1606 668 1610 672
rect 1614 668 1618 672
rect 1630 668 1634 672
rect 1734 668 1738 672
rect 2198 668 2202 672
rect 2222 668 2226 672
rect 2278 668 2282 672
rect 2286 668 2290 672
rect 3358 668 3362 672
rect 3430 668 3434 672
rect 3854 668 3858 672
rect 4150 668 4154 672
rect 4238 668 4242 672
rect 4246 668 4250 672
rect 302 658 306 662
rect 366 658 370 662
rect 1206 658 1210 662
rect 1598 658 1602 662
rect 1622 658 1626 662
rect 1638 658 1642 662
rect 1846 658 1850 662
rect 2030 658 2034 662
rect 2102 658 2106 662
rect 2126 658 2130 662
rect 2158 658 2162 662
rect 2486 658 2490 662
rect 2630 658 2634 662
rect 2726 658 2730 662
rect 2790 658 2794 662
rect 2814 658 2818 662
rect 3678 658 3682 662
rect 4182 658 4186 662
rect 4590 658 4594 662
rect 238 648 242 652
rect 1302 648 1306 652
rect 1430 648 1434 652
rect 1926 648 1930 652
rect 2006 648 2010 652
rect 2606 648 2610 652
rect 2766 648 2770 652
rect 3006 648 3010 652
rect 3126 648 3130 652
rect 3182 648 3186 652
rect 3270 648 3274 652
rect 3406 648 3410 652
rect 3470 648 3474 652
rect 3662 648 3666 652
rect 4118 648 4122 652
rect 406 638 410 642
rect 1270 638 1274 642
rect 1870 638 1874 642
rect 2414 638 2418 642
rect 3022 638 3026 642
rect 3286 638 3290 642
rect 3622 638 3626 642
rect 254 628 258 632
rect 646 628 650 632
rect 1862 628 1866 632
rect 4070 628 4074 632
rect 4350 628 4354 632
rect 1094 618 1098 622
rect 1286 618 1290 622
rect 1558 618 1562 622
rect 1798 618 1802 622
rect 2790 618 2794 622
rect 2830 618 2834 622
rect 2958 618 2962 622
rect 3182 618 3186 622
rect 3662 618 3666 622
rect 4214 618 4218 622
rect 4518 618 4522 622
rect 1934 608 1938 612
rect 2238 608 2242 612
rect 2422 608 2426 612
rect 2478 608 2482 612
rect 2518 608 2522 612
rect 3678 608 3682 612
rect 498 603 502 607
rect 506 603 509 607
rect 509 603 510 607
rect 1522 603 1526 607
rect 1530 603 1533 607
rect 1533 603 1534 607
rect 2546 603 2550 607
rect 2554 603 2557 607
rect 2557 603 2558 607
rect 3570 603 3574 607
rect 3578 603 3581 607
rect 3581 603 3582 607
rect 646 598 650 602
rect 2534 598 2538 602
rect 2654 598 2658 602
rect 3102 598 3106 602
rect 3862 598 3866 602
rect 3974 598 3978 602
rect 4206 598 4210 602
rect 4486 598 4490 602
rect 1126 588 1130 592
rect 1494 588 1498 592
rect 2126 588 2130 592
rect 2774 588 2778 592
rect 2990 588 2994 592
rect 3238 588 3242 592
rect 3702 588 3706 592
rect 4030 588 4034 592
rect 4070 588 4074 592
rect 2142 578 2146 582
rect 2606 578 2610 582
rect 2902 578 2906 582
rect 3086 578 3090 582
rect 3134 578 3138 582
rect 3598 578 3602 582
rect 790 568 794 572
rect 1334 568 1338 572
rect 2150 568 2154 572
rect 2254 568 2258 572
rect 2590 568 2594 572
rect 2870 568 2874 572
rect 3390 568 3394 572
rect 3694 568 3698 572
rect 3710 568 3714 572
rect 4310 568 4314 572
rect 1126 558 1130 562
rect 1694 558 1698 562
rect 1750 558 1754 562
rect 2014 558 2018 562
rect 2262 558 2266 562
rect 2374 558 2378 562
rect 2742 558 2746 562
rect 3014 558 3018 562
rect 3198 558 3202 562
rect 3262 558 3266 562
rect 3598 558 3602 562
rect 3622 558 3626 562
rect 3782 558 3786 562
rect 4390 558 4394 562
rect 4574 558 4578 562
rect 526 548 530 552
rect 942 548 946 552
rect 1134 548 1138 552
rect 1870 548 1874 552
rect 1982 548 1986 552
rect 2014 548 2018 552
rect 2118 548 2122 552
rect 2806 548 2810 552
rect 2886 548 2890 552
rect 2950 548 2954 552
rect 3070 548 3074 552
rect 3158 548 3162 552
rect 3422 548 3426 552
rect 3734 548 3738 552
rect 3822 548 3826 552
rect 4078 548 4082 552
rect 4454 548 4458 552
rect 4510 548 4514 552
rect 1422 538 1426 542
rect 1718 538 1722 542
rect 2110 538 2114 542
rect 2262 538 2266 542
rect 2638 538 2642 542
rect 3110 538 3114 542
rect 3118 538 3122 542
rect 3238 538 3242 542
rect 3406 538 3410 542
rect 3502 538 3506 542
rect 3942 538 3946 542
rect 4038 538 4042 542
rect 4134 538 4138 542
rect 4158 538 4162 542
rect 4214 538 4218 542
rect 4294 538 4298 542
rect 4566 538 4570 542
rect 1318 528 1322 532
rect 1654 528 1658 532
rect 1782 528 1786 532
rect 1838 528 1842 532
rect 1894 528 1898 532
rect 1942 528 1946 532
rect 2062 528 2066 532
rect 2190 528 2194 532
rect 2230 528 2234 532
rect 2798 528 2802 532
rect 3430 528 3434 532
rect 4054 528 4058 532
rect 326 518 330 522
rect 1142 518 1146 522
rect 1214 518 1218 522
rect 1854 518 1858 522
rect 2574 518 2578 522
rect 2790 518 2794 522
rect 2934 518 2938 522
rect 3174 518 3178 522
rect 3182 518 3186 522
rect 3206 518 3210 522
rect 3942 518 3946 522
rect 4270 518 4274 522
rect 1422 508 1426 512
rect 1430 508 1434 512
rect 1934 508 1938 512
rect 2222 508 2226 512
rect 2598 508 2602 512
rect 2822 508 2826 512
rect 3358 508 3362 512
rect 3422 508 3426 512
rect 1002 503 1006 507
rect 1010 503 1013 507
rect 1013 503 1014 507
rect 2026 503 2030 507
rect 2034 503 2037 507
rect 2037 503 2038 507
rect 3050 503 3054 507
rect 3058 503 3061 507
rect 3061 503 3062 507
rect 4082 503 4086 507
rect 4090 503 4093 507
rect 4093 503 4094 507
rect 310 498 314 502
rect 598 498 602 502
rect 1486 498 1490 502
rect 1910 498 1914 502
rect 2238 498 2242 502
rect 2486 498 2490 502
rect 2718 498 2722 502
rect 3086 498 3090 502
rect 3470 498 3474 502
rect 4014 498 4018 502
rect 4454 498 4458 502
rect 942 488 946 492
rect 2006 488 2010 492
rect 2046 488 2050 492
rect 2670 488 2674 492
rect 270 478 274 482
rect 1638 478 1642 482
rect 1790 478 1794 482
rect 3310 488 3314 492
rect 3494 488 3498 492
rect 3814 488 3818 492
rect 2582 478 2586 482
rect 3174 478 3178 482
rect 3510 478 3514 482
rect 3742 478 3746 482
rect 4054 478 4058 482
rect 4422 478 4426 482
rect 246 468 250 472
rect 390 468 394 472
rect 950 468 954 472
rect 1334 468 1338 472
rect 1614 468 1618 472
rect 1630 468 1634 472
rect 2054 468 2058 472
rect 2214 468 2218 472
rect 2398 468 2402 472
rect 2454 468 2458 472
rect 2502 468 2506 472
rect 2606 468 2610 472
rect 2822 468 2826 472
rect 2854 468 2858 472
rect 2894 468 2898 472
rect 2958 468 2962 472
rect 3350 468 3354 472
rect 4030 468 4034 472
rect 4342 468 4346 472
rect 4574 468 4578 472
rect 206 458 210 462
rect 262 458 266 462
rect 366 458 370 462
rect 694 458 698 462
rect 1206 458 1210 462
rect 1606 458 1610 462
rect 1678 458 1682 462
rect 1766 458 1770 462
rect 1814 458 1818 462
rect 1982 458 1986 462
rect 2238 458 2242 462
rect 2582 458 2586 462
rect 2646 458 2650 462
rect 2782 458 2786 462
rect 2878 458 2882 462
rect 3358 458 3362 462
rect 3854 458 3858 462
rect 4294 458 4298 462
rect 4358 458 4362 462
rect 4462 458 4466 462
rect 702 448 706 452
rect 1422 448 1426 452
rect 2070 448 2074 452
rect 2118 448 2122 452
rect 2238 448 2242 452
rect 2270 448 2274 452
rect 2622 448 2626 452
rect 2710 448 2714 452
rect 2806 448 2810 452
rect 2942 448 2946 452
rect 3070 448 3074 452
rect 3126 448 3130 452
rect 3230 448 3234 452
rect 3294 448 3298 452
rect 3662 448 3666 452
rect 3678 448 3682 452
rect 3694 448 3698 452
rect 3822 448 3826 452
rect 3830 448 3834 452
rect 3966 448 3970 452
rect 4462 448 4466 452
rect 4510 448 4514 452
rect 286 438 290 442
rect 294 438 298 442
rect 1246 438 1250 442
rect 2598 438 2602 442
rect 2702 438 2706 442
rect 3022 438 3026 442
rect 3406 438 3410 442
rect 3518 438 3522 442
rect 3702 438 3706 442
rect 4038 438 4042 442
rect 4182 438 4186 442
rect 4238 438 4242 442
rect 4310 438 4314 442
rect 4550 438 4554 442
rect 1438 428 1442 432
rect 1454 428 1458 432
rect 1854 428 1858 432
rect 1878 428 1882 432
rect 2014 428 2018 432
rect 2414 428 2418 432
rect 2430 428 2434 432
rect 2502 428 2506 432
rect 2750 428 2754 432
rect 3038 428 3042 432
rect 3902 428 3906 432
rect 1686 418 1690 422
rect 1798 418 1802 422
rect 2230 418 2234 422
rect 3102 418 3106 422
rect 3502 418 3506 422
rect 3758 418 3762 422
rect 1822 408 1826 412
rect 2734 408 2738 412
rect 3742 408 3746 412
rect 3846 408 3850 412
rect 498 403 502 407
rect 506 403 509 407
rect 509 403 510 407
rect 1522 403 1526 407
rect 1530 403 1533 407
rect 1533 403 1534 407
rect 2546 403 2550 407
rect 2554 403 2557 407
rect 2557 403 2558 407
rect 3570 403 3574 407
rect 3578 403 3581 407
rect 3581 403 3582 407
rect 198 398 202 402
rect 1134 398 1138 402
rect 2318 398 2322 402
rect 2502 398 2506 402
rect 2574 398 2578 402
rect 2678 398 2682 402
rect 3086 398 3090 402
rect 3206 398 3210 402
rect 3606 398 3610 402
rect 3966 398 3970 402
rect 4174 398 4178 402
rect 4334 398 4338 402
rect 2774 388 2778 392
rect 3662 388 3666 392
rect 1294 378 1298 382
rect 1934 378 1938 382
rect 2110 378 2114 382
rect 2654 378 2658 382
rect 2966 378 2970 382
rect 3806 378 3810 382
rect 3958 378 3962 382
rect 1710 368 1714 372
rect 1942 368 1946 372
rect 2142 368 2146 372
rect 222 358 226 362
rect 414 358 418 362
rect 1726 358 1730 362
rect 1750 358 1754 362
rect 1814 358 1818 362
rect 2462 368 2466 372
rect 2678 368 2682 372
rect 2726 368 2730 372
rect 2822 368 2826 372
rect 3446 368 3450 372
rect 3718 368 3722 372
rect 3814 368 3818 372
rect 4246 368 4250 372
rect 4254 368 4258 372
rect 4270 368 4274 372
rect 2126 358 2130 362
rect 2150 358 2154 362
rect 2390 358 2394 362
rect 2750 358 2754 362
rect 2846 358 2850 362
rect 3022 358 3026 362
rect 3158 358 3162 362
rect 3974 358 3978 362
rect 4246 358 4250 362
rect 4438 358 4442 362
rect 310 348 314 352
rect 1174 348 1178 352
rect 1438 348 1442 352
rect 1846 348 1850 352
rect 2350 348 2354 352
rect 2446 348 2450 352
rect 2462 348 2466 352
rect 2486 348 2490 352
rect 2694 348 2698 352
rect 2830 348 2834 352
rect 3150 348 3154 352
rect 3174 348 3178 352
rect 3646 348 3650 352
rect 3718 348 3722 352
rect 3998 348 4002 352
rect 4150 348 4154 352
rect 4230 348 4234 352
rect 4286 348 4290 352
rect 4582 348 4586 352
rect 350 338 354 342
rect 430 338 434 342
rect 766 338 770 342
rect 1574 338 1578 342
rect 1726 338 1730 342
rect 1838 338 1842 342
rect 2102 338 2106 342
rect 2478 338 2482 342
rect 2630 338 2634 342
rect 2678 338 2682 342
rect 2734 338 2738 342
rect 2766 338 2770 342
rect 2822 338 2826 342
rect 2982 338 2986 342
rect 3222 338 3226 342
rect 3286 338 3290 342
rect 3302 338 3306 342
rect 3758 338 3762 342
rect 3918 338 3922 342
rect 3974 338 3978 342
rect 3990 338 3994 342
rect 4054 338 4058 342
rect 4542 338 4546 342
rect 1678 328 1682 332
rect 1854 328 1858 332
rect 1982 328 1986 332
rect 2006 328 2010 332
rect 3022 328 3026 332
rect 3398 328 3402 332
rect 3406 328 3410 332
rect 3422 328 3426 332
rect 3670 328 3674 332
rect 3990 328 3994 332
rect 4014 328 4018 332
rect 4238 328 4242 332
rect 4254 328 4258 332
rect 4278 328 4282 332
rect 4494 328 4498 332
rect 254 318 258 322
rect 1070 318 1074 322
rect 1390 318 1394 322
rect 1606 318 1610 322
rect 1918 318 1922 322
rect 2150 318 2154 322
rect 2166 318 2170 322
rect 2766 318 2770 322
rect 2782 318 2786 322
rect 2814 318 2818 322
rect 2846 318 2850 322
rect 3094 318 3098 322
rect 3462 318 3466 322
rect 3486 318 3490 322
rect 3694 318 3698 322
rect 3734 318 3738 322
rect 2262 308 2266 312
rect 2606 308 2610 312
rect 2694 308 2698 312
rect 3174 308 3178 312
rect 3262 308 3266 312
rect 3590 308 3594 312
rect 3614 308 3618 312
rect 4070 308 4074 312
rect 4222 308 4226 312
rect 4446 308 4450 312
rect 1002 303 1006 307
rect 1010 303 1013 307
rect 1013 303 1014 307
rect 2026 303 2030 307
rect 2034 303 2037 307
rect 2037 303 2038 307
rect 3050 303 3054 307
rect 3058 303 3061 307
rect 3061 303 3062 307
rect 4082 303 4086 307
rect 4090 303 4093 307
rect 4093 303 4094 307
rect 310 298 314 302
rect 1134 298 1138 302
rect 1646 298 1650 302
rect 2014 298 2018 302
rect 2142 298 2146 302
rect 2710 298 2714 302
rect 3302 298 3306 302
rect 3510 298 3514 302
rect 4038 298 4042 302
rect 2590 288 2594 292
rect 3542 288 3546 292
rect 3550 288 3554 292
rect 4206 288 4210 292
rect 4486 288 4490 292
rect 278 278 282 282
rect 1030 278 1034 282
rect 2286 278 2290 282
rect 2294 278 2298 282
rect 2494 278 2498 282
rect 2614 278 2618 282
rect 2758 278 2762 282
rect 2766 278 2770 282
rect 3382 278 3386 282
rect 3454 278 3458 282
rect 3502 278 3506 282
rect 3670 278 3674 282
rect 3742 278 3746 282
rect 3974 278 3978 282
rect 4214 278 4218 282
rect 414 268 418 272
rect 1670 268 1674 272
rect 1830 268 1834 272
rect 1934 268 1938 272
rect 2590 268 2594 272
rect 2702 268 2706 272
rect 2958 268 2962 272
rect 3438 268 3442 272
rect 3678 268 3682 272
rect 3710 268 3714 272
rect 3814 268 3818 272
rect 3894 268 3898 272
rect 4150 268 4154 272
rect 262 258 266 262
rect 270 258 274 262
rect 606 258 610 262
rect 614 258 618 262
rect 1606 258 1610 262
rect 1910 258 1914 262
rect 2166 258 2170 262
rect 2670 258 2674 262
rect 2798 258 2802 262
rect 3190 258 3194 262
rect 3206 258 3210 262
rect 3350 258 3354 262
rect 3782 258 3786 262
rect 3934 258 3938 262
rect 4086 258 4090 262
rect 4214 258 4218 262
rect 4310 258 4314 262
rect 182 248 186 252
rect 246 248 250 252
rect 358 248 362 252
rect 1438 248 1442 252
rect 2190 248 2194 252
rect 2230 248 2234 252
rect 2438 248 2442 252
rect 2510 248 2514 252
rect 2542 248 2546 252
rect 2750 248 2754 252
rect 2934 248 2938 252
rect 2966 248 2970 252
rect 3078 248 3082 252
rect 3262 248 3266 252
rect 4294 248 4298 252
rect 4390 248 4394 252
rect 238 238 242 242
rect 294 238 298 242
rect 350 238 354 242
rect 1806 238 1810 242
rect 2238 238 2242 242
rect 2950 238 2954 242
rect 3310 238 3314 242
rect 3758 238 3762 242
rect 3942 238 3946 242
rect 4054 238 4058 242
rect 4078 238 4082 242
rect 4286 238 4290 242
rect 1454 228 1458 232
rect 2518 228 2522 232
rect 2622 228 2626 232
rect 2942 228 2946 232
rect 2982 228 2986 232
rect 3686 228 3690 232
rect 1398 218 1402 222
rect 3078 218 3082 222
rect 3478 218 3482 222
rect 3502 218 3506 222
rect 3718 218 3722 222
rect 3782 218 3786 222
rect 3918 218 3922 222
rect 4078 218 4082 222
rect 4094 218 4098 222
rect 1094 208 1098 212
rect 1894 208 1898 212
rect 2278 208 2282 212
rect 2494 208 2498 212
rect 3782 208 3786 212
rect 3982 208 3986 212
rect 4038 208 4042 212
rect 498 203 502 207
rect 506 203 509 207
rect 509 203 510 207
rect 1522 203 1526 207
rect 1530 203 1533 207
rect 1533 203 1534 207
rect 2546 203 2550 207
rect 2554 203 2557 207
rect 2557 203 2558 207
rect 3570 203 3574 207
rect 3578 203 3581 207
rect 3581 203 3582 207
rect 2790 198 2794 202
rect 3470 198 3474 202
rect 3558 198 3562 202
rect 3774 198 3778 202
rect 4262 198 4266 202
rect 4486 198 4490 202
rect 246 188 250 192
rect 1870 188 1874 192
rect 2862 188 2866 192
rect 2870 188 2874 192
rect 2974 188 2978 192
rect 3150 188 3154 192
rect 3886 188 3890 192
rect 326 178 330 182
rect 702 178 706 182
rect 1046 178 1050 182
rect 1142 178 1146 182
rect 1286 178 1290 182
rect 2350 178 2354 182
rect 2398 178 2402 182
rect 3918 178 3922 182
rect 3958 178 3962 182
rect 4318 178 4322 182
rect 2742 168 2746 172
rect 2950 168 2954 172
rect 2982 168 2986 172
rect 3126 168 3130 172
rect 3238 168 3242 172
rect 3806 168 3810 172
rect 4062 168 4066 172
rect 4150 168 4154 172
rect 4230 168 4234 172
rect 270 158 274 162
rect 430 158 434 162
rect 926 158 930 162
rect 1198 158 1202 162
rect 2134 158 2138 162
rect 3030 158 3034 162
rect 3038 158 3042 162
rect 3110 158 3114 162
rect 3254 158 3258 162
rect 3278 158 3282 162
rect 3318 158 3322 162
rect 3678 158 3682 162
rect 3702 158 3706 162
rect 3782 158 3786 162
rect 3942 158 3946 162
rect 4038 158 4042 162
rect 4158 158 4162 162
rect 4246 158 4250 162
rect 254 148 258 152
rect 950 148 954 152
rect 1694 148 1698 152
rect 2118 148 2122 152
rect 2374 148 2378 152
rect 2606 148 2610 152
rect 2742 148 2746 152
rect 2750 148 2754 152
rect 2774 148 2778 152
rect 3518 148 3522 152
rect 3606 148 3610 152
rect 4158 148 4162 152
rect 4166 148 4170 152
rect 4198 148 4202 152
rect 4214 148 4218 152
rect 4342 148 4346 152
rect 4374 148 4378 152
rect 4502 148 4506 152
rect 4542 148 4546 152
rect 2302 138 2306 142
rect 2366 138 2370 142
rect 2414 138 2418 142
rect 2430 138 2434 142
rect 2462 138 2466 142
rect 2798 138 2802 142
rect 2942 138 2946 142
rect 3014 138 3018 142
rect 3214 138 3218 142
rect 3222 138 3226 142
rect 3438 138 3442 142
rect 3534 138 3538 142
rect 3566 138 3570 142
rect 3590 138 3594 142
rect 3654 138 3658 142
rect 3742 138 3746 142
rect 3830 138 3834 142
rect 3854 138 3858 142
rect 3918 138 3922 142
rect 3934 138 3938 142
rect 3974 138 3978 142
rect 4038 138 4042 142
rect 4150 138 4154 142
rect 4206 138 4210 142
rect 4358 138 4362 142
rect 4534 138 4538 142
rect 2374 128 2378 132
rect 2382 128 2386 132
rect 2598 128 2602 132
rect 2646 128 2650 132
rect 3542 128 3546 132
rect 3598 128 3602 132
rect 3606 128 3610 132
rect 3766 128 3770 132
rect 3886 128 3890 132
rect 3902 128 3906 132
rect 3942 128 3946 132
rect 4054 128 4058 132
rect 4110 128 4114 132
rect 4166 128 4170 132
rect 4174 128 4178 132
rect 4334 128 4338 132
rect 4350 128 4354 132
rect 4438 128 4442 132
rect 1070 118 1074 122
rect 1518 118 1522 122
rect 1982 118 1986 122
rect 2150 118 2154 122
rect 2606 118 2610 122
rect 2630 118 2634 122
rect 3278 118 3282 122
rect 3366 118 3370 122
rect 3462 118 3466 122
rect 3590 118 3594 122
rect 4598 118 4602 122
rect 1390 108 1394 112
rect 2006 108 2010 112
rect 2278 108 2282 112
rect 2374 108 2378 112
rect 2774 108 2778 112
rect 2790 108 2794 112
rect 3174 108 3178 112
rect 3262 108 3266 112
rect 3366 108 3370 112
rect 3446 108 3450 112
rect 3558 108 3562 112
rect 3574 108 3578 112
rect 3774 108 3778 112
rect 3806 108 3810 112
rect 3870 108 3874 112
rect 3910 108 3914 112
rect 4070 108 4074 112
rect 4118 108 4122 112
rect 4126 108 4130 112
rect 4310 108 4314 112
rect 4350 108 4354 112
rect 1002 103 1006 107
rect 1010 103 1013 107
rect 1013 103 1014 107
rect 2026 103 2030 107
rect 2034 103 2037 107
rect 2037 103 2038 107
rect 3050 103 3054 107
rect 3058 103 3061 107
rect 3061 103 3062 107
rect 4082 103 4086 107
rect 4090 103 4093 107
rect 4093 103 4094 107
rect 918 98 922 102
rect 2198 98 2202 102
rect 2726 98 2730 102
rect 2814 98 2818 102
rect 2934 98 2938 102
rect 2958 98 2962 102
rect 3582 98 3586 102
rect 3662 98 3666 102
rect 4006 98 4010 102
rect 4110 98 4114 102
rect 4334 98 4338 102
rect 686 88 690 92
rect 694 88 698 92
rect 2422 88 2426 92
rect 2462 88 2466 92
rect 3846 88 3850 92
rect 3998 88 4002 92
rect 4102 88 4106 92
rect 4182 88 4186 92
rect 4190 88 4194 92
rect 4270 88 4274 92
rect 4278 88 4282 92
rect 4478 88 4482 92
rect 2286 78 2290 82
rect 2358 78 2362 82
rect 2630 78 2634 82
rect 3078 78 3082 82
rect 3158 78 3162 82
rect 3254 78 3258 82
rect 3310 78 3314 82
rect 3430 78 3434 82
rect 3718 78 3722 82
rect 3742 78 3746 82
rect 3774 78 3778 82
rect 3798 78 3802 82
rect 3838 78 3842 82
rect 3878 78 3882 82
rect 3910 78 3914 82
rect 3934 78 3938 82
rect 3974 78 3978 82
rect 4134 78 4138 82
rect 4262 78 4266 82
rect 4270 78 4274 82
rect 4342 78 4346 82
rect 4430 78 4434 82
rect 4534 78 4538 82
rect 942 68 946 72
rect 2270 68 2274 72
rect 2398 68 2402 72
rect 2510 68 2514 72
rect 2518 68 2522 72
rect 2566 68 2570 72
rect 2822 68 2826 72
rect 2838 68 2842 72
rect 2990 68 2994 72
rect 2998 68 3002 72
rect 3286 68 3290 72
rect 3526 68 3530 72
rect 3822 68 3826 72
rect 3862 68 3866 72
rect 3894 68 3898 72
rect 3950 68 3954 72
rect 4030 68 4034 72
rect 4046 68 4050 72
rect 4142 68 4146 72
rect 4174 68 4178 72
rect 4254 68 4258 72
rect 4270 68 4274 72
rect 4398 68 4402 72
rect 4526 68 4530 72
rect 574 58 578 62
rect 1046 58 1050 62
rect 1510 58 1514 62
rect 1806 58 1810 62
rect 3022 58 3026 62
rect 3046 58 3050 62
rect 3486 58 3490 62
rect 3726 58 3730 62
rect 3798 58 3802 62
rect 3854 58 3858 62
rect 3902 58 3906 62
rect 3918 58 3922 62
rect 3966 58 3970 62
rect 4022 58 4026 62
rect 4126 58 4130 62
rect 4342 58 4346 62
rect 2062 48 2066 52
rect 2238 48 2242 52
rect 2286 48 2290 52
rect 2870 48 2874 52
rect 2982 48 2986 52
rect 3022 48 3026 52
rect 3110 48 3114 52
rect 3118 48 3122 52
rect 3150 48 3154 52
rect 3246 48 3250 52
rect 3270 48 3274 52
rect 3294 48 3298 52
rect 3302 48 3306 52
rect 3598 48 3602 52
rect 3614 48 3618 52
rect 3758 48 3762 52
rect 3814 48 3818 52
rect 3846 48 3850 52
rect 3934 48 3938 52
rect 3966 48 3970 52
rect 4190 48 4194 52
rect 4230 48 4234 52
rect 4414 48 4418 52
rect 3790 38 3794 42
rect 4014 38 4018 42
rect 4198 38 4202 42
rect 4302 38 4306 42
rect 3318 28 3322 32
rect 3886 28 3890 32
rect 3950 28 3954 32
rect 4366 28 4370 32
rect 4382 28 4386 32
rect 3910 18 3914 22
rect 4078 18 4082 22
rect 4222 18 4226 22
rect 782 8 786 12
rect 1038 8 1042 12
rect 3958 8 3962 12
rect 498 3 502 7
rect 506 3 509 7
rect 509 3 510 7
rect 1522 3 1526 7
rect 1530 3 1533 7
rect 1533 3 1534 7
rect 2546 3 2550 7
rect 2554 3 2557 7
rect 2557 3 2558 7
rect 3570 3 3574 7
rect 3578 3 3581 7
rect 3581 3 3582 7
<< metal4 >>
rect 496 4403 498 4407
rect 502 4403 505 4407
rect 510 4403 512 4407
rect 1520 4403 1522 4407
rect 1526 4403 1529 4407
rect 1534 4403 1536 4407
rect 2544 4403 2546 4407
rect 2550 4403 2553 4407
rect 2558 4403 2560 4407
rect 3568 4403 3570 4407
rect 3574 4403 3577 4407
rect 3582 4403 3584 4407
rect 3826 4398 3833 4401
rect 4010 4398 4014 4401
rect 1762 4358 1769 4361
rect 790 4332 793 4358
rect 270 4152 273 4218
rect 174 3992 177 4078
rect 166 3978 174 3981
rect 166 3682 169 3978
rect 238 3792 241 4068
rect 246 4012 249 4128
rect 270 3912 273 4148
rect 302 3992 305 4268
rect 334 4142 337 4308
rect 354 4298 361 4301
rect 334 4052 337 4068
rect 358 4022 361 4298
rect 534 4252 537 4268
rect 522 4248 526 4251
rect 470 4232 473 4238
rect 496 4203 498 4207
rect 502 4203 505 4207
rect 510 4203 512 4207
rect 342 3872 345 3948
rect 358 3692 361 4018
rect 382 3862 385 4158
rect 422 3882 425 3948
rect 382 3672 385 3858
rect 406 3582 409 3738
rect 222 3458 230 3461
rect 6 3052 9 3068
rect 30 3042 33 3168
rect 150 3042 153 3148
rect 158 2992 161 3348
rect 222 2552 225 3458
rect 254 3122 257 3448
rect 298 3268 302 3271
rect 322 3268 326 3271
rect 302 3042 305 3168
rect 54 2462 57 2548
rect 214 1872 217 2308
rect 230 2282 233 2378
rect 302 2302 305 3038
rect 366 2902 369 3258
rect 398 3102 401 3548
rect 398 3002 401 3098
rect 398 2982 401 2998
rect 438 2892 441 3318
rect 318 2662 321 2718
rect 446 2512 449 3918
rect 462 3452 465 3558
rect 470 3482 473 4088
rect 486 4012 489 4048
rect 496 4003 498 4007
rect 502 4003 505 4007
rect 510 4003 512 4007
rect 478 3802 481 3928
rect 462 2912 465 3448
rect 470 3352 473 3478
rect 282 2068 286 2071
rect 194 1678 201 1681
rect 198 1622 201 1678
rect 158 1462 161 1548
rect 214 1472 217 1868
rect 230 1561 233 1918
rect 246 1862 249 2038
rect 310 1952 313 2088
rect 322 2068 326 2071
rect 334 1962 337 2188
rect 450 2148 454 2151
rect 470 2052 473 2268
rect 478 2082 481 2518
rect 458 2048 465 2051
rect 386 1968 390 1971
rect 318 1942 321 1958
rect 310 1731 313 1768
rect 310 1728 318 1731
rect 326 1662 329 1768
rect 350 1732 353 1868
rect 434 1848 441 1851
rect 226 1558 233 1561
rect 298 1548 302 1551
rect 330 1508 337 1511
rect 158 1332 161 1458
rect 334 1432 337 1508
rect 430 1492 433 1588
rect 438 1472 441 1848
rect 462 1712 465 2048
rect 478 1982 481 2008
rect 486 1822 489 3958
rect 496 3803 498 3807
rect 502 3803 505 3807
rect 510 3803 512 3807
rect 542 3662 545 4138
rect 574 3892 577 4118
rect 614 3792 617 4328
rect 678 4232 681 4318
rect 934 4312 937 4328
rect 1000 4303 1002 4307
rect 1006 4303 1009 4307
rect 1014 4303 1016 4307
rect 866 4268 870 4271
rect 810 4248 814 4251
rect 702 4162 705 4188
rect 634 4148 638 4151
rect 638 3942 641 4148
rect 496 3603 498 3607
rect 502 3603 505 3607
rect 510 3603 512 3607
rect 496 3403 498 3407
rect 502 3403 505 3407
rect 510 3403 512 3407
rect 494 3272 497 3278
rect 496 3203 498 3207
rect 502 3203 505 3207
rect 510 3203 512 3207
rect 542 3062 545 3658
rect 566 3542 569 3768
rect 566 3072 569 3538
rect 646 3332 649 3968
rect 710 3752 713 4248
rect 942 4242 945 4248
rect 958 4242 961 4288
rect 1562 4268 1566 4271
rect 1102 4262 1105 4268
rect 1202 4258 1206 4261
rect 718 4158 726 4161
rect 718 4122 721 4158
rect 798 3942 801 4148
rect 496 3003 498 3007
rect 502 3003 505 3007
rect 510 3003 512 3007
rect 566 2952 569 3068
rect 496 2803 498 2807
rect 502 2803 505 2807
rect 510 2803 512 2807
rect 614 2742 617 3318
rect 610 2648 614 2651
rect 496 2603 498 2607
rect 502 2603 505 2607
rect 510 2603 512 2607
rect 630 2562 633 2998
rect 646 2952 649 3328
rect 718 3292 721 3878
rect 766 3732 769 3938
rect 778 3738 782 3741
rect 806 3688 814 3691
rect 774 3638 782 3641
rect 726 3332 729 3518
rect 654 2912 657 3048
rect 662 2882 665 3118
rect 686 2862 689 3078
rect 694 2762 697 2888
rect 710 2752 713 2858
rect 642 2748 646 2751
rect 650 2678 654 2681
rect 682 2678 689 2681
rect 686 2562 689 2678
rect 694 2462 697 2718
rect 714 2648 718 2651
rect 726 2552 729 3148
rect 742 2962 745 3298
rect 750 3062 753 3078
rect 750 2942 753 3058
rect 734 2662 737 2748
rect 754 2658 758 2661
rect 496 2403 498 2407
rect 502 2403 505 2407
rect 510 2403 512 2407
rect 496 2203 498 2207
rect 502 2203 505 2207
rect 510 2203 512 2207
rect 646 2052 649 2128
rect 766 2062 769 3208
rect 774 2492 777 3638
rect 798 3562 801 3648
rect 798 3322 801 3558
rect 806 3222 809 3688
rect 830 3482 833 4068
rect 838 3972 841 4198
rect 1126 4192 1129 4258
rect 1246 4252 1249 4258
rect 1046 4142 1049 4148
rect 854 4042 857 4138
rect 1254 4132 1257 4168
rect 1306 4158 1310 4161
rect 838 3862 841 3958
rect 934 3892 937 3948
rect 774 2252 777 2268
rect 782 2082 785 3028
rect 814 2862 817 3168
rect 790 2672 793 2678
rect 802 2148 806 2151
rect 496 2003 498 2007
rect 502 2003 505 2007
rect 510 2003 512 2007
rect 550 1912 553 1958
rect 158 742 161 1328
rect 262 1312 265 1388
rect 230 1062 233 1268
rect 302 1072 305 1268
rect 318 1128 326 1131
rect 222 842 225 998
rect 310 962 313 1108
rect 318 942 321 1128
rect 350 1052 353 1368
rect 398 1162 401 1168
rect 406 1152 409 1188
rect 430 1062 433 1278
rect 486 1262 489 1818
rect 496 1803 498 1807
rect 502 1803 505 1807
rect 510 1803 512 1807
rect 550 1802 553 1908
rect 496 1603 498 1607
rect 502 1603 505 1607
rect 510 1603 512 1607
rect 514 1548 518 1551
rect 550 1442 553 1688
rect 496 1403 498 1407
rect 502 1403 505 1407
rect 510 1403 512 1407
rect 558 1342 561 1508
rect 566 1332 569 1488
rect 574 1462 577 1778
rect 598 1652 601 1678
rect 654 1632 657 1698
rect 766 1692 769 2018
rect 782 1782 785 2078
rect 814 2051 817 2818
rect 826 2658 830 2661
rect 854 2182 857 3088
rect 910 3082 913 3658
rect 926 3338 934 3341
rect 926 3282 929 3338
rect 966 3272 969 3818
rect 990 3662 993 4128
rect 1000 4103 1002 4107
rect 1006 4103 1009 4107
rect 1014 4103 1016 4107
rect 1102 4022 1105 4038
rect 1000 3903 1002 3907
rect 1006 3903 1009 3907
rect 1014 3903 1016 3907
rect 1034 3838 1041 3841
rect 1000 3703 1002 3707
rect 1006 3703 1009 3707
rect 1014 3703 1016 3707
rect 1000 3503 1002 3507
rect 1006 3503 1009 3507
rect 1014 3503 1016 3507
rect 1022 3492 1025 3708
rect 1038 3692 1041 3838
rect 1000 3303 1002 3307
rect 1006 3303 1009 3307
rect 1014 3303 1016 3307
rect 1000 3103 1002 3107
rect 1006 3103 1009 3107
rect 1014 3103 1016 3107
rect 850 2138 854 2141
rect 862 2072 865 2788
rect 870 2062 873 2888
rect 810 2048 817 2051
rect 806 1741 809 2048
rect 862 1762 865 2058
rect 870 1992 873 2058
rect 878 2052 881 2878
rect 890 2748 894 2751
rect 890 2688 894 2691
rect 898 2328 902 2331
rect 878 1772 881 2048
rect 894 2032 897 2068
rect 902 1942 905 2308
rect 902 1842 905 1938
rect 802 1738 809 1741
rect 602 1578 606 1581
rect 366 952 369 1058
rect 198 402 201 738
rect 206 462 209 468
rect 222 362 225 838
rect 310 762 313 778
rect 366 762 369 948
rect 406 718 414 721
rect 242 648 246 651
rect 182 252 185 268
rect 238 242 241 258
rect 246 252 249 468
rect 254 322 257 628
rect 278 481 281 668
rect 306 658 310 661
rect 274 478 281 481
rect 262 262 265 458
rect 278 282 281 478
rect 286 442 289 458
rect 246 192 249 248
rect 270 162 273 258
rect 294 242 297 438
rect 310 352 313 498
rect 310 302 313 348
rect 326 182 329 518
rect 366 462 369 658
rect 406 642 409 718
rect 430 652 433 718
rect 446 682 449 1258
rect 496 1203 498 1207
rect 502 1203 505 1207
rect 510 1203 512 1207
rect 542 1202 545 1258
rect 458 1158 462 1161
rect 490 1158 494 1161
rect 526 1132 529 1178
rect 496 1003 498 1007
rect 502 1003 505 1007
rect 510 1003 512 1007
rect 558 842 561 858
rect 496 803 498 807
rect 502 803 505 807
rect 510 803 512 807
rect 582 752 585 798
rect 574 748 582 751
rect 496 603 498 607
rect 502 603 505 607
rect 510 603 512 607
rect 526 552 529 678
rect 558 662 561 678
rect 386 468 390 471
rect 496 403 498 407
rect 502 403 505 407
rect 510 403 512 407
rect 350 242 353 338
rect 414 272 417 358
rect 362 248 366 251
rect 430 162 433 338
rect 496 203 498 207
rect 502 203 505 207
rect 510 203 512 207
rect 258 148 262 151
rect 574 62 577 748
rect 598 502 601 1458
rect 654 1162 657 1628
rect 766 1352 769 1688
rect 778 1578 782 1581
rect 790 1462 793 1698
rect 750 1252 753 1318
rect 678 782 681 1098
rect 766 762 769 1348
rect 806 1152 809 1738
rect 846 1362 849 1598
rect 910 1431 913 3078
rect 1000 2903 1002 2907
rect 1006 2903 1009 2907
rect 1014 2903 1016 2907
rect 1034 2858 1038 2861
rect 1000 2703 1002 2707
rect 1006 2703 1009 2707
rect 1014 2703 1016 2707
rect 1022 2612 1025 2618
rect 1030 2592 1033 2858
rect 918 2472 921 2478
rect 926 2472 929 2558
rect 1000 2503 1002 2507
rect 1006 2503 1009 2507
rect 1014 2503 1016 2507
rect 1038 2482 1041 2488
rect 1006 2472 1009 2478
rect 930 2338 934 2341
rect 946 2328 950 2331
rect 922 1968 926 1971
rect 922 1938 926 1941
rect 934 1662 937 2218
rect 966 1882 969 2088
rect 974 1792 977 2108
rect 910 1428 921 1431
rect 902 1272 905 1368
rect 646 602 649 628
rect 614 262 617 268
rect 606 252 609 258
rect 686 92 689 118
rect 694 92 697 458
rect 702 182 705 448
rect 766 342 769 738
rect 790 672 793 1148
rect 918 1082 921 1428
rect 934 1062 937 1658
rect 942 1132 945 1428
rect 970 1038 977 1041
rect 938 868 942 871
rect 974 862 977 1038
rect 982 942 985 2398
rect 1000 2303 1002 2307
rect 1006 2303 1009 2307
rect 1014 2303 1016 2307
rect 990 2102 993 2118
rect 1000 2103 1002 2107
rect 1006 2103 1009 2107
rect 1014 2103 1016 2107
rect 1006 2072 1009 2078
rect 1000 1903 1002 1907
rect 1006 1903 1009 1907
rect 1014 1903 1016 1907
rect 1000 1703 1002 1707
rect 1006 1703 1009 1707
rect 1014 1703 1016 1707
rect 1022 1512 1025 1558
rect 1038 1552 1041 2278
rect 1046 1542 1049 2838
rect 1054 2692 1057 3658
rect 1062 2942 1065 3748
rect 1078 2482 1081 3548
rect 1102 3212 1105 3828
rect 1110 3692 1113 3898
rect 1230 3392 1233 3428
rect 1078 2272 1081 2288
rect 1086 2282 1089 2558
rect 1102 2282 1105 2688
rect 1134 2192 1137 3348
rect 1070 2062 1073 2088
rect 1078 2082 1081 2188
rect 1102 2072 1105 2078
rect 1126 1892 1129 1928
rect 1134 1872 1137 2158
rect 1142 1932 1145 1948
rect 1106 1728 1110 1731
rect 1000 1503 1002 1507
rect 1006 1503 1009 1507
rect 1014 1503 1016 1507
rect 1054 1362 1057 1558
rect 1000 1303 1002 1307
rect 1006 1303 1009 1307
rect 1014 1303 1016 1307
rect 1000 1103 1002 1107
rect 1006 1103 1009 1107
rect 1014 1103 1016 1107
rect 1054 1032 1057 1148
rect 1086 1132 1089 1308
rect 1142 1212 1145 1378
rect 1014 942 1017 958
rect 1070 952 1073 958
rect 1078 942 1081 958
rect 1000 903 1002 907
rect 1006 903 1009 907
rect 1014 903 1016 907
rect 1122 868 1126 871
rect 1000 703 1002 707
rect 1006 703 1009 707
rect 1014 703 1016 707
rect 790 11 793 568
rect 942 492 945 548
rect 1000 503 1002 507
rect 1006 503 1009 507
rect 1014 503 1016 507
rect 930 158 934 161
rect 918 62 921 98
rect 942 72 945 488
rect 950 152 953 468
rect 1000 303 1002 307
rect 1006 303 1009 307
rect 1014 303 1016 307
rect 1000 103 1002 107
rect 1006 103 1009 107
rect 1014 103 1016 107
rect 786 8 793 11
rect 1030 11 1033 278
rect 1046 62 1049 178
rect 1070 122 1073 318
rect 1094 212 1097 618
rect 1126 562 1129 588
rect 1134 552 1137 998
rect 1150 742 1153 2438
rect 1158 1692 1161 1748
rect 1158 1262 1161 1658
rect 1166 1482 1169 3278
rect 1222 2922 1225 2948
rect 1194 2468 1198 2471
rect 1206 2392 1209 2468
rect 1246 1912 1249 2068
rect 1190 1662 1193 1798
rect 1198 1742 1201 1768
rect 1206 1682 1209 1788
rect 1226 1728 1230 1731
rect 1218 1708 1225 1711
rect 1222 1692 1225 1708
rect 1230 1682 1233 1688
rect 1202 1558 1206 1561
rect 1178 1268 1182 1271
rect 1178 1168 1182 1171
rect 1166 931 1169 998
rect 1190 952 1193 1108
rect 1198 1102 1201 1188
rect 1166 928 1174 931
rect 1158 892 1161 928
rect 1134 402 1137 548
rect 1134 302 1137 398
rect 1142 182 1145 518
rect 1174 352 1177 908
rect 1190 892 1193 948
rect 1198 872 1201 958
rect 1186 848 1190 851
rect 1206 662 1209 1268
rect 1222 1252 1225 1298
rect 1222 1152 1225 1248
rect 1230 1072 1233 1328
rect 1238 1092 1241 1668
rect 1246 1232 1249 1518
rect 1218 948 1222 951
rect 1214 842 1217 868
rect 1214 522 1217 838
rect 1202 458 1206 461
rect 1246 442 1249 1168
rect 1254 742 1257 2918
rect 1270 2622 1273 3948
rect 1278 3001 1281 3798
rect 1302 3122 1305 3928
rect 1298 3088 1302 3091
rect 1278 2998 1286 3001
rect 1274 2338 1278 2341
rect 1262 1742 1265 2058
rect 1274 1948 1278 1951
rect 1294 1932 1297 2518
rect 1302 1682 1305 2208
rect 1318 1682 1321 3388
rect 1350 3252 1353 3838
rect 1330 2658 1334 2661
rect 1326 2152 1329 2178
rect 1334 2132 1337 2148
rect 1342 1692 1345 3228
rect 1358 2502 1361 4258
rect 1366 2442 1369 4258
rect 1466 4238 1470 4241
rect 1442 4158 1446 4161
rect 1398 4002 1401 4088
rect 1398 3792 1401 3998
rect 1406 3862 1409 4148
rect 1486 4022 1489 4258
rect 1494 4062 1497 4218
rect 1520 4203 1522 4207
rect 1526 4203 1529 4207
rect 1534 4203 1536 4207
rect 1694 4152 1697 4188
rect 1502 3892 1505 4058
rect 1520 4003 1522 4007
rect 1526 4003 1529 4007
rect 1534 4003 1536 4007
rect 1522 3958 1526 3961
rect 1494 3872 1497 3888
rect 1382 3252 1385 3778
rect 1398 3552 1401 3738
rect 1406 3232 1409 3858
rect 1478 3352 1481 3838
rect 1520 3803 1522 3807
rect 1526 3803 1529 3807
rect 1534 3803 1536 3807
rect 1520 3603 1522 3607
rect 1526 3603 1529 3607
rect 1534 3603 1536 3607
rect 1498 3548 1502 3551
rect 1518 3542 1521 3548
rect 1590 3442 1593 3658
rect 1520 3403 1522 3407
rect 1526 3403 1529 3407
rect 1534 3403 1536 3407
rect 1478 3212 1481 3348
rect 1406 3142 1409 3208
rect 1382 2892 1385 3068
rect 1306 1678 1310 1681
rect 1262 1162 1265 1458
rect 1286 1222 1289 1428
rect 1310 1421 1313 1468
rect 1350 1462 1353 1498
rect 1310 1418 1318 1421
rect 1286 1132 1289 1148
rect 1294 1061 1297 1208
rect 1358 1102 1361 2388
rect 1366 2302 1369 2438
rect 1366 1252 1369 1358
rect 1294 1058 1302 1061
rect 1366 982 1369 1098
rect 1374 932 1377 2368
rect 1382 1882 1385 2618
rect 1406 2162 1409 2788
rect 1414 2752 1417 3198
rect 1486 2802 1489 3238
rect 1520 3203 1522 3207
rect 1526 3203 1529 3207
rect 1534 3203 1536 3207
rect 1520 3003 1522 3007
rect 1526 3003 1529 3007
rect 1534 3003 1536 3007
rect 1538 2948 1542 2951
rect 1520 2803 1522 2807
rect 1526 2803 1529 2807
rect 1534 2803 1536 2807
rect 1418 2748 1422 2751
rect 1454 2492 1457 2518
rect 1414 2362 1417 2368
rect 1386 1748 1390 1751
rect 1414 1412 1417 1418
rect 1382 1252 1385 1278
rect 1406 1162 1409 1308
rect 1414 1282 1417 1408
rect 1406 1132 1409 1158
rect 1286 918 1294 921
rect 1270 848 1278 851
rect 1270 642 1273 848
rect 1286 622 1289 918
rect 1374 872 1377 928
rect 1286 182 1289 618
rect 1294 382 1297 718
rect 1302 652 1305 678
rect 1326 531 1329 858
rect 1410 848 1414 851
rect 1334 702 1337 848
rect 1322 528 1329 531
rect 1334 472 1337 568
rect 1194 158 1198 161
rect 1390 112 1393 318
rect 1398 222 1401 718
rect 1422 542 1425 2468
rect 1430 2032 1433 2168
rect 1430 2001 1433 2028
rect 1430 1998 1438 2001
rect 1446 1552 1449 1678
rect 1454 1552 1457 1558
rect 1446 1472 1449 1548
rect 1430 512 1433 648
rect 1422 452 1425 508
rect 1438 432 1441 1228
rect 1446 1082 1449 1468
rect 1462 1372 1465 1418
rect 1454 1132 1457 1268
rect 1454 962 1457 1068
rect 1462 672 1465 888
rect 1470 871 1473 2658
rect 1486 1792 1489 2798
rect 1558 2692 1561 3058
rect 1520 2603 1522 2607
rect 1526 2603 1529 2607
rect 1534 2603 1536 2607
rect 1566 2592 1569 3128
rect 1574 3092 1577 3128
rect 1582 2862 1585 3018
rect 1494 1371 1497 2428
rect 1520 2403 1522 2407
rect 1526 2403 1529 2407
rect 1534 2403 1536 2407
rect 1520 2203 1522 2207
rect 1526 2203 1529 2207
rect 1534 2203 1536 2207
rect 1542 2142 1545 2428
rect 1562 2408 1566 2411
rect 1510 2122 1513 2138
rect 1542 2102 1545 2138
rect 1502 1812 1505 1828
rect 1510 1762 1513 2008
rect 1520 2003 1522 2007
rect 1526 2003 1529 2007
rect 1534 2003 1536 2007
rect 1542 1982 1545 1998
rect 1520 1803 1522 1807
rect 1526 1803 1529 1807
rect 1534 1803 1536 1807
rect 1542 1752 1545 1758
rect 1520 1603 1522 1607
rect 1526 1603 1529 1607
rect 1534 1603 1536 1607
rect 1520 1403 1522 1407
rect 1526 1403 1529 1407
rect 1534 1403 1536 1407
rect 1494 1368 1502 1371
rect 1478 1061 1481 1358
rect 1486 1102 1489 1148
rect 1510 1092 1513 1388
rect 1542 1262 1545 1268
rect 1520 1203 1522 1207
rect 1526 1203 1529 1207
rect 1534 1203 1536 1207
rect 1478 1058 1486 1061
rect 1520 1003 1522 1007
rect 1526 1003 1529 1007
rect 1534 1003 1536 1007
rect 1486 942 1489 948
rect 1478 892 1481 918
rect 1470 868 1478 871
rect 1520 803 1522 807
rect 1526 803 1529 807
rect 1534 803 1536 807
rect 1550 772 1553 2358
rect 1558 1342 1561 2408
rect 1566 2052 1569 2068
rect 1566 1882 1569 1888
rect 1558 1328 1566 1331
rect 1558 622 1561 1328
rect 1566 782 1569 928
rect 1566 752 1569 778
rect 1520 603 1522 607
rect 1526 603 1529 607
rect 1534 603 1536 607
rect 1486 588 1494 591
rect 1486 502 1489 588
rect 1438 252 1441 348
rect 1454 232 1457 428
rect 1520 403 1522 407
rect 1526 403 1529 407
rect 1534 403 1536 407
rect 1574 342 1577 2858
rect 1590 2272 1593 3438
rect 1610 3138 1614 3141
rect 1586 2268 1590 2271
rect 1598 2242 1601 2258
rect 1598 2082 1601 2238
rect 1606 2212 1609 2918
rect 1638 2652 1641 2698
rect 1646 2492 1649 2868
rect 1662 2592 1665 3948
rect 1686 3152 1689 3308
rect 1670 3082 1673 3088
rect 1678 2771 1681 3118
rect 1678 2768 1686 2771
rect 1606 1682 1609 2208
rect 1602 1528 1609 1531
rect 1586 1328 1590 1331
rect 1606 1242 1609 1528
rect 1614 1502 1617 2378
rect 1590 842 1593 908
rect 1598 752 1601 1188
rect 1606 942 1609 1168
rect 1614 1112 1617 1498
rect 1622 1492 1625 2188
rect 1630 1662 1633 1948
rect 1638 1872 1641 2438
rect 1662 2412 1665 2498
rect 1646 1741 1649 2288
rect 1662 1852 1665 2058
rect 1638 1738 1649 1741
rect 1622 1462 1625 1488
rect 1598 662 1601 748
rect 1606 742 1609 938
rect 1638 912 1641 1738
rect 1662 1662 1665 1698
rect 1658 1478 1662 1481
rect 1646 1422 1649 1428
rect 1658 1258 1662 1261
rect 1650 1248 1654 1251
rect 1642 908 1649 911
rect 1618 878 1622 881
rect 1606 672 1609 738
rect 1614 672 1617 868
rect 1630 772 1633 898
rect 1614 472 1617 668
rect 1622 662 1625 728
rect 1630 622 1633 668
rect 1638 662 1641 888
rect 1646 682 1649 908
rect 1630 472 1633 528
rect 1638 482 1641 658
rect 1646 528 1654 531
rect 1606 422 1609 458
rect 1606 322 1609 418
rect 1646 302 1649 528
rect 1670 272 1673 2748
rect 1726 2662 1729 2678
rect 1726 2332 1729 2548
rect 1758 2322 1761 4338
rect 1766 4322 1769 4358
rect 1818 4268 1822 4271
rect 1986 4238 1990 4241
rect 1934 4182 1937 4228
rect 1794 4158 1798 4161
rect 1766 4142 1769 4148
rect 1766 3991 1769 4088
rect 1838 4072 1841 4078
rect 1766 3988 1774 3991
rect 1782 3492 1785 4058
rect 1846 4032 1849 4148
rect 1910 4141 1913 4148
rect 1910 4138 1918 4141
rect 1918 3982 1921 4058
rect 1810 3958 1814 3961
rect 1770 3348 1774 3351
rect 1778 3248 1782 3251
rect 1790 3092 1793 3638
rect 1798 3602 1801 3698
rect 1846 3662 1849 3708
rect 1814 3552 1817 3558
rect 1806 3152 1809 3408
rect 1770 2668 1774 2671
rect 1806 2592 1809 3148
rect 1850 3058 1854 3061
rect 1806 2462 1809 2468
rect 1694 2142 1697 2188
rect 1694 2042 1697 2118
rect 1702 2071 1705 2198
rect 1774 2142 1777 2168
rect 1734 2132 1737 2138
rect 1702 2068 1710 2071
rect 1778 2058 1782 2061
rect 1694 2012 1697 2038
rect 1678 1292 1681 1998
rect 1718 1962 1721 1988
rect 1690 1858 1694 1861
rect 1686 1152 1689 1778
rect 1694 1512 1697 1768
rect 1694 1332 1697 1508
rect 1702 1482 1705 1668
rect 1726 1551 1729 2018
rect 1734 1948 1742 1951
rect 1734 1832 1737 1948
rect 1742 1882 1745 1898
rect 1766 1881 1769 1978
rect 1774 1962 1777 1968
rect 1782 1942 1785 1978
rect 1766 1878 1774 1881
rect 1742 1862 1745 1878
rect 1790 1862 1793 2078
rect 1846 2002 1849 3058
rect 1862 3002 1865 3258
rect 1882 3088 1886 3091
rect 1838 1932 1841 1948
rect 1826 1928 1830 1931
rect 1762 1858 1766 1861
rect 1738 1768 1742 1771
rect 1754 1648 1758 1651
rect 1718 1548 1729 1551
rect 1710 1482 1713 1488
rect 1694 1212 1697 1328
rect 1702 1312 1705 1478
rect 1702 1172 1705 1308
rect 1678 922 1681 1008
rect 1686 952 1689 1148
rect 1718 1072 1721 1548
rect 1726 1372 1729 1538
rect 1730 1258 1734 1261
rect 1742 1152 1745 1608
rect 1678 882 1681 918
rect 1686 912 1689 948
rect 1694 872 1697 1028
rect 1694 562 1697 868
rect 1718 792 1721 1068
rect 1730 918 1734 921
rect 1742 862 1745 978
rect 1738 668 1742 671
rect 1750 562 1753 1588
rect 1766 1542 1769 1788
rect 1790 1572 1793 1858
rect 1758 882 1761 968
rect 1722 538 1726 541
rect 1766 462 1769 1458
rect 1774 1052 1777 1488
rect 1790 1482 1793 1568
rect 1798 1222 1801 1898
rect 1842 1828 1846 1831
rect 1842 1538 1846 1541
rect 1802 1218 1809 1221
rect 1774 742 1777 748
rect 1782 532 1785 938
rect 1790 482 1793 858
rect 1678 332 1681 458
rect 1686 422 1689 428
rect 1798 422 1801 618
rect 1710 362 1713 368
rect 1746 358 1750 361
rect 1726 342 1729 358
rect 1602 258 1606 261
rect 1806 242 1809 1218
rect 1814 1152 1817 1458
rect 1838 1232 1841 1538
rect 1814 932 1817 1108
rect 1854 1072 1857 1768
rect 1862 1012 1865 2228
rect 1886 1612 1889 2918
rect 1902 2902 1905 3748
rect 1910 3292 1913 3958
rect 1918 3912 1921 3978
rect 1918 3492 1921 3798
rect 1918 3362 1921 3488
rect 1926 2892 1929 4038
rect 1958 3992 1961 4228
rect 1966 3932 1969 4128
rect 1974 4112 1977 4118
rect 1986 3988 1993 3991
rect 1950 3838 1958 3841
rect 1950 3522 1953 3838
rect 1958 3662 1961 3698
rect 1966 3492 1969 3848
rect 1990 3652 1993 3988
rect 1998 3952 2001 4388
rect 2024 4303 2026 4307
rect 2030 4303 2033 4307
rect 2038 4303 2040 4307
rect 2082 4288 2086 4291
rect 2266 4288 2270 4291
rect 2006 4252 2009 4258
rect 2024 4103 2026 4107
rect 2030 4103 2033 4107
rect 2038 4103 2040 4107
rect 2006 3842 2009 4038
rect 2086 3922 2089 4128
rect 2110 4082 2113 4268
rect 2170 4258 2174 4261
rect 2154 4248 2158 4251
rect 2274 4248 2278 4251
rect 2286 4192 2289 4268
rect 2238 4182 2241 4188
rect 2206 4131 2209 4158
rect 2206 4128 2217 4131
rect 2024 3903 2026 3907
rect 2030 3903 2033 3907
rect 2038 3903 2040 3907
rect 2090 3868 2094 3871
rect 2024 3703 2026 3707
rect 2030 3703 2033 3707
rect 2038 3703 2040 3707
rect 1978 3548 1982 3551
rect 2006 3532 2009 3538
rect 1946 3468 1950 3471
rect 1934 3272 1937 3288
rect 1914 2888 1918 2891
rect 1902 2772 1905 2778
rect 1902 2362 1905 2458
rect 1918 2271 1921 2318
rect 1918 2268 1926 2271
rect 1894 2011 1897 2028
rect 1894 2008 1902 2011
rect 1910 1942 1913 1988
rect 1902 1802 1905 1878
rect 1902 1672 1905 1798
rect 1870 1541 1873 1558
rect 1870 1538 1878 1541
rect 1870 1372 1873 1378
rect 1878 1282 1881 1428
rect 1886 1312 1889 1318
rect 1894 1232 1897 1528
rect 1902 1172 1905 1508
rect 1918 1502 1921 2008
rect 1926 1592 1929 2068
rect 1938 1918 1942 1921
rect 1946 1648 1950 1651
rect 1966 1611 1969 3488
rect 1982 2492 1985 3508
rect 1990 3152 1993 3358
rect 1990 3091 1993 3148
rect 1990 3088 1998 3091
rect 1990 2532 1993 2548
rect 1974 1982 1977 2038
rect 1974 1712 1977 1978
rect 1974 1682 1977 1708
rect 1958 1608 1969 1611
rect 1958 1412 1961 1608
rect 1970 1328 1977 1331
rect 1974 1322 1977 1328
rect 1910 1242 1913 1248
rect 1814 761 1817 838
rect 1814 758 1822 761
rect 1846 742 1849 748
rect 1814 362 1817 458
rect 1822 412 1825 688
rect 1846 662 1849 738
rect 1838 362 1841 528
rect 1854 522 1857 928
rect 1862 882 1865 998
rect 1870 642 1873 1118
rect 1886 1001 1889 1148
rect 1886 998 1894 1001
rect 1934 972 1937 1058
rect 1882 968 1886 971
rect 1878 952 1881 958
rect 1878 772 1881 798
rect 1878 752 1881 758
rect 1866 628 1870 631
rect 1886 551 1889 858
rect 1874 548 1889 551
rect 1878 432 1881 548
rect 1894 532 1897 958
rect 1910 502 1913 748
rect 1926 652 1929 928
rect 1942 912 1945 1138
rect 1958 1061 1961 1168
rect 1958 1058 1966 1061
rect 1950 692 1953 1058
rect 1982 942 1985 2128
rect 1990 1872 1993 1908
rect 1990 1452 1993 1588
rect 1998 1321 2001 2958
rect 2006 2762 2009 3518
rect 2014 3292 2017 3638
rect 2024 3503 2026 3507
rect 2030 3503 2033 3507
rect 2038 3503 2040 3507
rect 2026 3468 2030 3471
rect 2024 3303 2026 3307
rect 2030 3303 2033 3307
rect 2038 3303 2040 3307
rect 2024 3103 2026 3107
rect 2030 3103 2033 3107
rect 2038 3103 2040 3107
rect 2046 3042 2049 3058
rect 2026 2948 2030 2951
rect 2014 2942 2017 2948
rect 2024 2903 2026 2907
rect 2030 2903 2033 2907
rect 2038 2903 2040 2907
rect 2046 2892 2049 2898
rect 2024 2703 2026 2707
rect 2030 2703 2033 2707
rect 2038 2703 2040 2707
rect 2024 2503 2026 2507
rect 2030 2503 2033 2507
rect 2038 2503 2040 2507
rect 2014 2251 2017 2318
rect 2024 2303 2026 2307
rect 2030 2303 2033 2307
rect 2038 2303 2040 2307
rect 2014 2248 2022 2251
rect 2006 2032 2009 2248
rect 2046 2122 2049 2628
rect 2014 2112 2017 2118
rect 2024 2103 2026 2107
rect 2030 2103 2033 2107
rect 2038 2103 2040 2107
rect 2054 2032 2057 3748
rect 2066 3738 2070 3741
rect 2102 3632 2105 3878
rect 2110 3822 2113 3968
rect 2118 3792 2121 3988
rect 2174 3872 2177 3958
rect 2182 3952 2185 3958
rect 2130 3658 2134 3661
rect 2094 3342 2097 3478
rect 2110 3352 2113 3358
rect 2098 3258 2102 3261
rect 2006 1932 2009 2028
rect 2024 1903 2026 1907
rect 2030 1903 2033 1907
rect 2038 1903 2040 1907
rect 2024 1703 2026 1707
rect 2030 1703 2033 1707
rect 2038 1703 2040 1707
rect 2054 1702 2057 1958
rect 2024 1503 2026 1507
rect 2030 1503 2033 1507
rect 2038 1503 2040 1507
rect 1990 1318 2001 1321
rect 1990 1192 1993 1318
rect 2024 1303 2026 1307
rect 2030 1303 2033 1307
rect 2038 1303 2040 1307
rect 2046 1202 2049 1508
rect 1994 1128 1998 1131
rect 2050 1128 2054 1131
rect 1998 1092 2001 1098
rect 1958 852 1961 918
rect 1934 512 1937 608
rect 1982 552 1985 828
rect 1838 342 1841 358
rect 1846 342 1849 348
rect 1854 332 1857 428
rect 1830 272 1833 278
rect 1910 262 1913 498
rect 1918 322 1921 348
rect 1934 272 1937 378
rect 1942 372 1945 528
rect 1990 482 1993 1058
rect 1998 1052 2001 1088
rect 2006 1022 2009 1108
rect 2024 1103 2026 1107
rect 2030 1103 2033 1107
rect 2038 1103 2040 1107
rect 2006 712 2009 998
rect 2034 978 2038 981
rect 2018 958 2022 961
rect 2024 903 2026 907
rect 2030 903 2033 907
rect 2038 903 2040 907
rect 2014 852 2017 858
rect 2024 703 2026 707
rect 2030 703 2033 707
rect 2038 703 2040 707
rect 2030 662 2033 688
rect 2038 682 2041 688
rect 2006 492 2009 648
rect 2014 562 2017 568
rect 1974 461 1977 478
rect 1974 458 1982 461
rect 2014 432 2017 548
rect 2046 542 2049 1068
rect 2054 992 2057 998
rect 2062 941 2065 3148
rect 2082 3138 2086 3141
rect 2070 2692 2073 3088
rect 2078 2422 2081 2618
rect 2070 1072 2073 1618
rect 2086 1052 2089 2828
rect 2094 2772 2097 2778
rect 2110 2762 2113 2938
rect 2118 2852 2121 3038
rect 2110 2732 2113 2758
rect 2118 2692 2121 2848
rect 2126 2772 2129 3318
rect 2134 2592 2137 3618
rect 2150 3102 2153 3668
rect 2162 3558 2166 3561
rect 2158 3192 2161 3208
rect 2166 3192 2169 3558
rect 2146 2938 2150 2941
rect 2158 2832 2161 2878
rect 2130 2548 2134 2551
rect 2102 1682 2105 2178
rect 2126 2062 2129 2338
rect 2174 2332 2177 2998
rect 2182 2272 2185 3278
rect 2198 3182 2201 3958
rect 2214 3592 2217 4128
rect 2222 4022 2225 4158
rect 2238 3842 2241 4108
rect 2246 3872 2249 3878
rect 2254 3762 2257 4148
rect 2302 4042 2305 4338
rect 2270 3702 2273 3908
rect 2270 3652 2273 3688
rect 2214 3282 2217 3398
rect 2214 3082 2217 3268
rect 2222 3162 2225 3168
rect 2206 2982 2209 3008
rect 2190 2662 2193 2678
rect 2114 1938 2121 1941
rect 2118 1832 2121 1938
rect 2094 1262 2097 1308
rect 2102 1272 2105 1498
rect 2094 1062 2097 1258
rect 2102 1072 2105 1268
rect 2110 1212 2113 1818
rect 2134 1342 2137 2058
rect 2158 2032 2161 2048
rect 2150 1922 2153 1938
rect 2190 1932 2193 2578
rect 2214 2502 2217 3018
rect 2190 1852 2193 1878
rect 2174 1842 2177 1848
rect 2110 1092 2113 1118
rect 2054 938 2065 941
rect 2054 802 2057 938
rect 2086 932 2089 1028
rect 2062 928 2070 931
rect 2062 832 2065 928
rect 2110 862 2113 1058
rect 2126 902 2129 1158
rect 2024 503 2026 507
rect 2030 503 2033 507
rect 2038 503 2040 507
rect 2046 492 2049 538
rect 2054 472 2057 578
rect 2066 528 2073 531
rect 2070 452 2073 528
rect 2102 342 2105 658
rect 2110 542 2113 858
rect 2118 552 2121 888
rect 2126 872 2129 878
rect 2126 852 2129 858
rect 2126 662 2129 748
rect 2126 592 2129 598
rect 2110 382 2113 538
rect 1982 322 1985 328
rect 1886 208 1894 211
rect 1520 203 1522 207
rect 1526 203 1529 207
rect 1534 203 1536 207
rect 1870 182 1873 188
rect 1886 162 1889 208
rect 1690 148 1694 151
rect 1514 118 1518 121
rect 1986 118 1990 121
rect 2006 112 2009 328
rect 2024 303 2026 307
rect 2030 303 2033 307
rect 2038 303 2040 307
rect 2014 292 2017 298
rect 2118 152 2121 448
rect 2126 362 2129 368
rect 2134 162 2137 1338
rect 2150 1262 2153 1458
rect 2142 1091 2145 1158
rect 2142 1088 2150 1091
rect 2142 842 2145 968
rect 2158 942 2161 1838
rect 2198 1512 2201 2398
rect 2206 2142 2209 2338
rect 2214 2152 2217 2158
rect 2206 1822 2209 2138
rect 2210 1788 2214 1791
rect 2222 1762 2225 3068
rect 2230 2962 2233 3488
rect 2246 2972 2249 3368
rect 2254 3272 2257 3388
rect 2262 3362 2265 3618
rect 2278 3572 2281 3828
rect 2254 3072 2257 3268
rect 2262 3252 2265 3258
rect 2270 3182 2273 3518
rect 2302 3402 2305 3798
rect 2302 3351 2305 3358
rect 2298 3348 2305 3351
rect 2278 3318 2286 3321
rect 2278 3312 2281 3318
rect 2282 3288 2286 3291
rect 2266 3078 2270 3081
rect 2286 3032 2289 3198
rect 2234 2948 2238 2951
rect 2282 2938 2286 2941
rect 2294 2802 2297 3338
rect 2258 2648 2262 2651
rect 2166 1042 2169 1478
rect 2190 1422 2193 1438
rect 2206 1392 2209 1618
rect 2214 1332 2217 1508
rect 2174 992 2177 1078
rect 2206 1032 2209 1078
rect 2194 948 2198 951
rect 2142 582 2145 678
rect 2150 572 2153 868
rect 2158 781 2161 928
rect 2230 912 2233 2458
rect 2238 2282 2241 2288
rect 2238 2102 2241 2128
rect 2238 1912 2241 1918
rect 2246 1892 2249 2388
rect 2262 2272 2265 2348
rect 2270 2292 2273 2448
rect 2302 2412 2305 3258
rect 2310 3172 2313 3538
rect 2318 3372 2321 4208
rect 2334 4152 2337 4268
rect 2410 4258 2417 4261
rect 2334 4062 2337 4148
rect 2342 3771 2345 4148
rect 2350 4122 2353 4138
rect 2358 4102 2361 4118
rect 2390 4042 2393 4058
rect 2366 3772 2369 3788
rect 2342 3768 2350 3771
rect 2338 3718 2342 3721
rect 2326 3662 2329 3678
rect 2326 3542 2329 3588
rect 2334 3442 2337 3708
rect 2350 3422 2353 3508
rect 2358 3402 2361 3728
rect 2366 3432 2369 3678
rect 2314 3108 2318 3111
rect 2318 3062 2321 3068
rect 2310 2862 2313 2878
rect 2326 2752 2329 3208
rect 2310 2632 2313 2738
rect 2318 2592 2321 2628
rect 2318 2472 2321 2588
rect 2334 2492 2337 3388
rect 2342 3302 2345 3368
rect 2342 3202 2345 3268
rect 2350 3252 2353 3378
rect 2374 3352 2377 3818
rect 2350 3202 2353 3218
rect 2342 2982 2345 3038
rect 2350 2892 2353 3128
rect 2358 3112 2361 3298
rect 2366 3052 2369 3318
rect 2374 2972 2377 3328
rect 2382 3322 2385 3928
rect 2390 3562 2393 3878
rect 2390 3442 2393 3518
rect 2398 3332 2401 4258
rect 2414 4232 2417 4258
rect 2414 4172 2417 4188
rect 2422 3982 2425 4328
rect 2478 4242 2481 4268
rect 2506 4248 2510 4251
rect 2430 4162 2433 4178
rect 2442 4078 2446 4081
rect 2470 4062 2473 4078
rect 2510 4052 2513 4168
rect 2526 4162 2529 4348
rect 2534 4212 2537 4268
rect 2650 4248 2654 4251
rect 2662 4242 2665 4318
rect 2678 4212 2681 4358
rect 2544 4203 2546 4207
rect 2550 4203 2553 4207
rect 2558 4203 2560 4207
rect 2762 4188 2766 4191
rect 2654 4082 2657 4118
rect 2662 4092 2665 4118
rect 2634 4078 2638 4081
rect 2626 4068 2630 4071
rect 2590 4062 2593 4068
rect 2498 4048 2502 4051
rect 2618 4048 2622 4051
rect 2406 3892 2409 3938
rect 2406 3342 2409 3888
rect 2414 3512 2417 3538
rect 2422 3522 2425 3528
rect 2430 3432 2433 3628
rect 2414 3372 2417 3388
rect 2394 3308 2398 3311
rect 2382 3162 2385 3168
rect 2390 3092 2393 3238
rect 2406 3152 2409 3318
rect 2350 2872 2353 2888
rect 2350 2612 2353 2828
rect 2390 2692 2393 2998
rect 2390 2672 2393 2688
rect 2334 2472 2337 2488
rect 2294 2332 2297 2378
rect 2254 2032 2257 2048
rect 2254 2002 2257 2008
rect 2246 1662 2249 1738
rect 2254 1332 2257 1928
rect 2262 1742 2265 2238
rect 2270 2142 2273 2288
rect 2270 1832 2273 2088
rect 2294 2062 2297 2328
rect 2302 2122 2305 2408
rect 2366 2371 2369 2518
rect 2390 2462 2393 2498
rect 2366 2368 2374 2371
rect 2362 2328 2366 2331
rect 2382 2268 2390 2271
rect 2382 2262 2385 2268
rect 2326 2242 2329 2258
rect 2310 2182 2313 2198
rect 2302 2052 2305 2058
rect 2302 1982 2305 1988
rect 2282 1728 2286 1731
rect 2270 1522 2273 1538
rect 2278 1472 2281 1598
rect 2262 1342 2265 1448
rect 2278 1361 2281 1468
rect 2278 1358 2286 1361
rect 2246 1272 2249 1278
rect 2242 1248 2246 1251
rect 2246 1131 2249 1158
rect 2242 1128 2249 1131
rect 2222 878 2230 881
rect 2170 858 2174 861
rect 2158 778 2166 781
rect 2174 718 2182 721
rect 2158 582 2161 658
rect 2142 302 2145 368
rect 2150 362 2153 568
rect 2174 492 2177 718
rect 2198 672 2201 748
rect 2194 668 2198 671
rect 2214 671 2217 878
rect 2222 872 2225 878
rect 2230 852 2233 858
rect 2214 668 2222 671
rect 2162 318 2166 321
rect 2150 312 2153 318
rect 2162 258 2166 261
rect 2190 252 2193 528
rect 2222 512 2225 668
rect 2218 468 2222 471
rect 2230 422 2233 528
rect 2238 502 2241 608
rect 2254 572 2257 1328
rect 2262 1202 2265 1338
rect 2318 1262 2321 1918
rect 2334 1892 2337 2078
rect 2334 1882 2337 1888
rect 2330 1718 2334 1721
rect 2342 1682 2345 2148
rect 2350 1982 2353 2218
rect 2398 2152 2401 2948
rect 2406 2862 2409 2888
rect 2406 2102 2409 2698
rect 2414 2392 2417 3368
rect 2422 2832 2425 3068
rect 2430 2602 2433 3388
rect 2438 3112 2441 3598
rect 2446 3382 2449 4008
rect 2544 4003 2546 4007
rect 2550 4003 2553 4007
rect 2558 4003 2560 4007
rect 2566 3952 2569 3998
rect 2490 3878 2494 3881
rect 2494 3862 2497 3868
rect 2502 3852 2505 3868
rect 2566 3852 2569 3858
rect 2546 3848 2550 3851
rect 2544 3803 2546 3807
rect 2550 3803 2553 3807
rect 2558 3803 2560 3807
rect 2534 3772 2537 3798
rect 2530 3758 2534 3761
rect 2454 3572 2457 3688
rect 2470 3652 2473 3658
rect 2482 3568 2486 3571
rect 2462 3171 2465 3178
rect 2458 3168 2465 3171
rect 2478 3172 2481 3528
rect 2486 3322 2489 3468
rect 2494 3172 2497 3598
rect 2502 3592 2505 3598
rect 2506 3568 2510 3571
rect 2518 3522 2521 3648
rect 2502 3202 2505 3418
rect 2526 3392 2529 3398
rect 2518 3362 2521 3368
rect 2522 3328 2526 3331
rect 2534 3292 2537 3738
rect 2558 3652 2561 3658
rect 2574 3642 2577 3898
rect 2544 3603 2546 3607
rect 2550 3603 2553 3607
rect 2558 3603 2560 3607
rect 2590 3602 2593 3628
rect 2544 3403 2546 3407
rect 2550 3403 2553 3407
rect 2558 3403 2560 3407
rect 2554 3318 2558 3321
rect 2494 3122 2497 3138
rect 2478 3118 2486 3121
rect 2438 3102 2441 3108
rect 2418 2228 2422 2231
rect 2406 2072 2409 2078
rect 2406 2052 2409 2058
rect 2358 1722 2361 2018
rect 2374 1952 2377 1958
rect 2370 1868 2374 1871
rect 2334 1512 2337 1538
rect 2314 1248 2318 1251
rect 2310 1208 2318 1211
rect 2270 942 2273 1078
rect 2302 892 2305 1068
rect 2310 871 2313 1208
rect 2318 972 2321 1008
rect 2310 868 2318 871
rect 2266 748 2270 751
rect 2270 712 2273 748
rect 2274 668 2278 671
rect 2294 671 2297 788
rect 2290 668 2297 671
rect 2266 558 2273 561
rect 2238 462 2241 498
rect 2230 242 2233 248
rect 2238 242 2241 448
rect 2262 312 2265 538
rect 2270 452 2273 558
rect 2318 402 2321 828
rect 2326 582 2329 1098
rect 2334 1062 2337 1508
rect 2342 1312 2345 1468
rect 2350 1182 2353 1548
rect 2358 1422 2361 1658
rect 2366 1362 2369 1558
rect 2390 1482 2393 1538
rect 2398 1502 2401 1618
rect 2358 1352 2361 1358
rect 2342 862 2345 868
rect 2338 838 2342 841
rect 2334 742 2337 788
rect 2350 352 2353 1148
rect 2358 762 2361 1098
rect 2366 952 2369 958
rect 2382 882 2385 1358
rect 2390 1272 2393 1458
rect 2414 1192 2417 2068
rect 2430 1962 2433 2188
rect 2438 2072 2441 3088
rect 2454 2922 2457 2938
rect 2462 2872 2465 3118
rect 2478 2812 2481 3118
rect 2534 3082 2537 3258
rect 2544 3203 2546 3207
rect 2550 3203 2553 3207
rect 2558 3203 2560 3207
rect 2486 3072 2489 3078
rect 2454 2142 2457 2678
rect 2462 2592 2465 2708
rect 2486 2692 2489 3018
rect 2494 2932 2497 2938
rect 2518 2932 2521 2948
rect 2502 2862 2505 2868
rect 2494 2692 2497 2728
rect 2462 2332 2465 2538
rect 2462 2142 2465 2328
rect 2442 2058 2446 2061
rect 2430 1691 2433 1958
rect 2462 1742 2465 1778
rect 2430 1688 2438 1691
rect 2466 1468 2470 1471
rect 2438 1332 2441 1408
rect 2458 1348 2462 1351
rect 2394 1148 2398 1151
rect 2402 1138 2406 1141
rect 2394 938 2398 941
rect 2406 902 2409 958
rect 2414 942 2417 948
rect 2382 852 2385 868
rect 2402 728 2406 731
rect 2414 712 2417 738
rect 2370 558 2374 561
rect 2398 472 2401 518
rect 2414 432 2417 638
rect 2422 612 2425 1158
rect 2430 1152 2433 1158
rect 2430 432 2433 1138
rect 2446 1072 2449 1108
rect 2454 1062 2457 1328
rect 2470 1162 2473 1468
rect 2478 1462 2481 2488
rect 2518 2481 2521 2888
rect 2526 2542 2529 2758
rect 2534 2722 2537 3008
rect 2544 3003 2546 3007
rect 2550 3003 2553 3007
rect 2558 3003 2560 3007
rect 2566 2962 2569 3298
rect 2574 3202 2577 3268
rect 2606 3261 2609 3708
rect 2622 3472 2625 3928
rect 2630 3572 2633 3958
rect 2602 3258 2609 3261
rect 2566 2842 2569 2958
rect 2614 2952 2617 3258
rect 2630 3242 2633 3318
rect 2638 3292 2641 3548
rect 2654 3522 2657 3538
rect 2646 3462 2649 3468
rect 2622 3122 2625 3138
rect 2544 2803 2546 2807
rect 2550 2803 2553 2807
rect 2558 2803 2560 2807
rect 2544 2603 2546 2607
rect 2550 2603 2553 2607
rect 2558 2603 2560 2607
rect 2518 2478 2526 2481
rect 2506 2458 2510 2461
rect 2566 2422 2569 2778
rect 2544 2403 2546 2407
rect 2550 2403 2553 2407
rect 2558 2403 2560 2407
rect 2566 2262 2569 2408
rect 2574 2282 2577 2808
rect 2590 2482 2593 2858
rect 2614 2762 2617 2858
rect 2614 2592 2617 2678
rect 2594 2478 2598 2481
rect 2582 2352 2585 2478
rect 2544 2203 2546 2207
rect 2550 2203 2553 2207
rect 2558 2203 2560 2207
rect 2566 2202 2569 2248
rect 2542 2132 2545 2188
rect 2586 2158 2590 2161
rect 2606 2152 2609 2498
rect 2630 2302 2633 2868
rect 2590 2071 2593 2078
rect 2586 2068 2593 2071
rect 2494 1932 2497 2008
rect 2526 1952 2529 2068
rect 2544 2003 2546 2007
rect 2550 2003 2553 2007
rect 2558 2003 2560 2007
rect 2566 1982 2569 1998
rect 2626 1868 2630 1871
rect 2544 1803 2546 1807
rect 2550 1803 2553 1807
rect 2558 1803 2560 1807
rect 2494 1732 2497 1738
rect 2486 1672 2489 1698
rect 2502 1512 2505 1598
rect 2478 1448 2486 1451
rect 2478 1442 2481 1448
rect 2478 1382 2481 1438
rect 2494 1262 2497 1478
rect 2478 1112 2481 1148
rect 2474 1098 2478 1101
rect 2494 1082 2497 1088
rect 2438 752 2441 1058
rect 2502 982 2505 1508
rect 2510 1352 2513 1758
rect 2518 1602 2521 1788
rect 2622 1732 2625 1748
rect 2630 1692 2633 1828
rect 2526 1682 2529 1688
rect 2630 1622 2633 1668
rect 2544 1603 2546 1607
rect 2550 1603 2553 1607
rect 2558 1603 2560 1607
rect 2554 1548 2558 1551
rect 2534 1412 2537 1428
rect 2544 1403 2546 1407
rect 2550 1403 2553 1407
rect 2558 1403 2560 1407
rect 2446 382 2449 928
rect 2458 868 2462 871
rect 2478 871 2481 978
rect 2502 962 2505 978
rect 2474 868 2481 871
rect 2486 882 2489 918
rect 2474 838 2478 841
rect 2486 752 2489 878
rect 2498 868 2502 871
rect 2510 862 2513 1258
rect 2518 962 2521 1278
rect 2518 952 2521 958
rect 2510 832 2513 838
rect 2510 792 2513 808
rect 2490 658 2494 661
rect 2518 612 2521 928
rect 2526 752 2529 1378
rect 2542 1272 2545 1278
rect 2544 1203 2546 1207
rect 2550 1203 2553 1207
rect 2558 1203 2560 1207
rect 2574 1132 2577 1248
rect 2544 1003 2546 1007
rect 2550 1003 2553 1007
rect 2558 1003 2560 1007
rect 2550 952 2553 968
rect 2546 948 2550 951
rect 2544 803 2546 807
rect 2550 803 2553 807
rect 2558 803 2560 807
rect 2534 782 2537 798
rect 2566 772 2569 798
rect 2574 702 2577 948
rect 2458 468 2462 471
rect 2390 362 2393 368
rect 2462 352 2465 368
rect 2294 282 2297 308
rect 2150 122 2153 148
rect 2024 103 2026 107
rect 2030 103 2033 107
rect 2038 103 2040 107
rect 2198 102 2201 138
rect 2278 112 2281 208
rect 2286 82 2289 278
rect 2446 251 2449 348
rect 2478 342 2481 608
rect 2534 602 2537 688
rect 2544 603 2546 607
rect 2550 603 2553 607
rect 2558 603 2560 607
rect 2486 352 2489 498
rect 2502 432 2505 468
rect 2502 402 2505 428
rect 2544 403 2546 407
rect 2550 403 2553 407
rect 2558 403 2560 407
rect 2574 402 2577 518
rect 2582 482 2585 1248
rect 2590 1132 2593 1468
rect 2610 1268 2614 1271
rect 2622 1182 2625 1538
rect 2638 1392 2641 3288
rect 2646 3162 2649 3168
rect 2646 2902 2649 3098
rect 2654 3062 2657 3498
rect 2662 3172 2665 3728
rect 2670 3432 2673 3558
rect 2670 3272 2673 3428
rect 2678 3411 2681 4188
rect 2686 4162 2689 4168
rect 2706 4058 2710 4061
rect 2694 3662 2697 3688
rect 2686 3442 2689 3488
rect 2702 3432 2705 4008
rect 2710 3722 2713 3878
rect 2718 3752 2721 3908
rect 2714 3688 2718 3691
rect 2710 3522 2713 3658
rect 2718 3562 2721 3678
rect 2726 3412 2729 4148
rect 2738 3708 2745 3711
rect 2742 3692 2745 3708
rect 2734 3452 2737 3668
rect 2678 3408 2686 3411
rect 2678 3392 2681 3398
rect 2666 3158 2670 3161
rect 2694 3102 2697 3318
rect 2706 3308 2713 3311
rect 2710 3302 2713 3308
rect 2734 3172 2737 3378
rect 2742 3112 2745 3688
rect 2750 3662 2753 3998
rect 2758 3162 2761 3808
rect 2766 3682 2769 3938
rect 2766 3032 2769 3588
rect 2774 3131 2777 3568
rect 2798 3492 2801 4178
rect 2814 4142 2817 4328
rect 3048 4303 3050 4307
rect 3054 4303 3057 4307
rect 3062 4303 3064 4307
rect 2842 4268 2846 4271
rect 2830 4062 2833 4068
rect 2798 3452 2801 3458
rect 2782 3372 2785 3418
rect 2774 3128 2785 3131
rect 2686 2892 2689 2908
rect 2670 2652 2673 2698
rect 2678 2492 2681 2568
rect 2654 2212 2657 2408
rect 2662 2272 2665 2398
rect 2678 2242 2681 2298
rect 2658 2158 2662 2161
rect 2678 2152 2681 2188
rect 2666 2088 2670 2091
rect 2646 1912 2649 1938
rect 2658 1868 2662 1871
rect 2650 1728 2657 1731
rect 2654 1722 2657 1728
rect 2670 1672 2673 1978
rect 2678 1952 2681 1958
rect 2670 1652 2673 1668
rect 2662 1452 2665 1568
rect 2670 1542 2673 1548
rect 2646 1372 2649 1388
rect 2590 1022 2593 1068
rect 2606 962 2609 1148
rect 2630 1142 2633 1368
rect 2642 1348 2646 1351
rect 2666 1328 2670 1331
rect 2614 1062 2617 1118
rect 2622 1062 2625 1098
rect 2590 832 2593 928
rect 2598 822 2601 948
rect 2590 762 2593 768
rect 2614 762 2617 1028
rect 2638 1002 2641 1088
rect 2646 1022 2649 1318
rect 2662 1292 2665 1318
rect 2678 1292 2681 1568
rect 2654 1242 2657 1258
rect 2654 1222 2657 1238
rect 2658 1138 2662 1141
rect 2678 1082 2681 1088
rect 2654 1052 2657 1068
rect 2622 962 2625 978
rect 2610 718 2614 721
rect 2606 652 2609 698
rect 2622 692 2625 718
rect 2630 662 2633 918
rect 2590 562 2593 568
rect 2586 458 2590 461
rect 2598 442 2601 508
rect 2606 472 2609 578
rect 2638 542 2641 758
rect 2610 468 2617 471
rect 2442 248 2449 251
rect 2302 142 2305 248
rect 2350 172 2353 178
rect 2378 148 2382 151
rect 2366 132 2369 138
rect 2382 132 2385 148
rect 2374 122 2377 128
rect 2374 112 2377 118
rect 2358 82 2361 88
rect 2398 82 2401 178
rect 2414 142 2417 228
rect 2494 212 2497 278
rect 2590 272 2593 288
rect 2542 252 2545 258
rect 2506 248 2510 251
rect 2518 232 2521 238
rect 2544 203 2546 207
rect 2550 203 2553 207
rect 2558 203 2560 207
rect 2606 152 2609 308
rect 2614 282 2617 468
rect 2646 462 2649 958
rect 2654 782 2657 1048
rect 2674 928 2678 931
rect 2662 702 2665 738
rect 2626 448 2630 451
rect 2654 382 2657 598
rect 2630 342 2633 348
rect 2670 262 2673 488
rect 2678 402 2681 678
rect 2678 352 2681 368
rect 2678 332 2681 338
rect 2686 282 2689 2288
rect 2694 1782 2697 2268
rect 2702 2132 2705 2358
rect 2710 2272 2713 2568
rect 2726 2552 2729 3028
rect 2774 3012 2777 3118
rect 2782 2962 2785 3128
rect 2722 2338 2726 2341
rect 2734 2302 2737 2728
rect 2750 2592 2753 2918
rect 2750 2562 2753 2578
rect 2758 2472 2761 2858
rect 2790 2842 2793 3318
rect 2798 3232 2801 3328
rect 2806 3182 2809 4018
rect 2830 3972 2833 3998
rect 2814 3872 2817 3898
rect 2814 3372 2817 3438
rect 2830 3402 2833 3798
rect 2838 3642 2841 3658
rect 2838 3442 2841 3578
rect 2846 3552 2849 3658
rect 2854 3392 2857 4098
rect 2894 4062 2897 4128
rect 3070 4112 3073 4348
rect 3234 4338 3238 4341
rect 3358 4338 3366 4341
rect 2874 3868 2878 3871
rect 2902 3862 2905 3878
rect 2870 3702 2873 3838
rect 2890 3678 2894 3681
rect 2862 3652 2865 3658
rect 2870 3522 2873 3658
rect 2874 3468 2881 3471
rect 2822 3222 2825 3388
rect 2830 3162 2833 3318
rect 2838 3182 2841 3388
rect 2878 3372 2881 3468
rect 2886 3452 2889 3478
rect 2894 3382 2897 3538
rect 2910 3482 2913 4108
rect 3048 4103 3050 4107
rect 3054 4103 3057 4107
rect 3062 4103 3064 4107
rect 2918 3382 2921 3498
rect 2878 3312 2881 3338
rect 2910 3312 2913 3338
rect 2874 3218 2878 3221
rect 2854 3152 2857 3188
rect 2878 3152 2881 3158
rect 2774 2482 2777 2628
rect 2782 2542 2785 2608
rect 2814 2532 2817 2568
rect 2758 2342 2761 2358
rect 2778 2278 2782 2281
rect 2750 2272 2753 2278
rect 2806 2232 2809 2388
rect 2814 2312 2817 2358
rect 2702 2081 2705 2128
rect 2702 2078 2710 2081
rect 2726 2072 2729 2098
rect 2702 1942 2705 1948
rect 2726 1932 2729 2068
rect 2822 2052 2825 3078
rect 2846 3032 2849 3128
rect 2862 3102 2865 3148
rect 2874 3128 2878 3131
rect 2846 2892 2849 2918
rect 2846 2652 2849 2658
rect 2830 2532 2833 2568
rect 2838 2522 2841 2528
rect 2830 2352 2833 2368
rect 2750 1882 2753 1888
rect 2702 1872 2705 1878
rect 2830 1858 2838 1861
rect 2694 1692 2697 1758
rect 2710 1612 2713 1628
rect 2698 1518 2702 1521
rect 2710 1462 2713 1578
rect 2726 1532 2729 1688
rect 2698 1458 2702 1461
rect 2726 1392 2729 1528
rect 2718 1272 2721 1288
rect 2702 1248 2710 1251
rect 2702 1122 2705 1248
rect 2698 1048 2702 1051
rect 2694 892 2697 908
rect 2694 842 2697 848
rect 2694 692 2697 728
rect 2702 692 2705 928
rect 2710 812 2713 1208
rect 2726 1132 2729 1378
rect 2734 1362 2737 1558
rect 2742 1532 2745 1548
rect 2746 1478 2750 1481
rect 2766 1382 2769 1598
rect 2734 1272 2737 1298
rect 2718 1112 2721 1118
rect 2718 1072 2721 1078
rect 2726 1062 2729 1128
rect 2726 942 2729 1058
rect 2702 642 2705 688
rect 2718 682 2721 928
rect 2726 872 2729 878
rect 2726 852 2729 858
rect 2726 762 2729 838
rect 2734 752 2737 1228
rect 2742 1202 2745 1358
rect 2750 1282 2753 1288
rect 2742 1142 2745 1168
rect 2766 1152 2769 1308
rect 2742 1002 2745 1138
rect 2750 1052 2753 1068
rect 2742 862 2745 868
rect 2718 502 2721 648
rect 2718 451 2721 458
rect 2714 448 2721 451
rect 2702 442 2705 448
rect 2694 312 2697 348
rect 2702 272 2705 378
rect 2710 302 2713 378
rect 2726 372 2729 658
rect 2738 558 2742 561
rect 2750 432 2753 928
rect 2758 901 2761 1148
rect 2766 1052 2769 1058
rect 2766 912 2769 928
rect 2774 922 2777 1248
rect 2782 1162 2785 1678
rect 2782 982 2785 1158
rect 2790 972 2793 1548
rect 2798 1242 2801 1258
rect 2798 1152 2801 1188
rect 2798 1062 2801 1148
rect 2806 962 2809 1778
rect 2814 1732 2817 1758
rect 2830 1722 2833 1858
rect 2842 1688 2846 1691
rect 2822 1092 2825 1658
rect 2854 1632 2857 2928
rect 2862 2572 2865 2878
rect 2874 2868 2878 2871
rect 2886 2852 2889 3298
rect 2874 2678 2878 2681
rect 2866 2478 2870 2481
rect 2866 2458 2870 2461
rect 2886 2352 2889 2518
rect 2894 2362 2897 2908
rect 2902 2752 2905 3068
rect 2910 3052 2913 3258
rect 2918 3182 2921 3348
rect 2918 2962 2921 3058
rect 2910 2752 2913 2918
rect 2910 2622 2913 2718
rect 2902 2542 2905 2558
rect 2902 2292 2905 2328
rect 2902 2252 2905 2258
rect 2894 2232 2897 2248
rect 2910 1712 2913 2618
rect 2918 2422 2921 2488
rect 2926 2392 2929 3948
rect 2938 3668 2942 3671
rect 2950 3652 2953 3668
rect 2990 3472 2993 3618
rect 2934 3452 2937 3458
rect 2934 3362 2937 3378
rect 2934 3002 2937 3298
rect 2942 3282 2945 3468
rect 2958 3382 2961 3468
rect 2998 3432 3001 3738
rect 3006 3421 3009 3798
rect 3014 3452 3017 3648
rect 3022 3462 3025 3468
rect 3006 3418 3017 3421
rect 3006 3362 3009 3408
rect 2970 3358 2974 3361
rect 2994 3348 2998 3351
rect 2970 3338 2974 3341
rect 2942 3132 2945 3268
rect 2962 3258 2969 3261
rect 2966 3242 2969 3258
rect 2966 2912 2969 3238
rect 2934 2572 2937 2778
rect 2974 2632 2977 3318
rect 2930 2278 2934 2281
rect 2942 2262 2945 2408
rect 2934 2082 2937 2258
rect 2946 2148 2950 2151
rect 2942 1932 2945 1948
rect 2938 1928 2942 1931
rect 2950 1882 2953 2078
rect 2958 1942 2961 2518
rect 2926 1682 2929 1718
rect 2934 1682 2937 1828
rect 2966 1762 2969 2518
rect 2982 2402 2985 3278
rect 3014 3172 3017 3418
rect 2990 2632 2993 3128
rect 2998 3058 3006 3061
rect 2998 2712 3001 3058
rect 3022 2971 3025 3288
rect 3030 3182 3033 4008
rect 3038 3412 3041 4078
rect 3048 3903 3050 3907
rect 3054 3903 3057 3907
rect 3062 3903 3064 3907
rect 3074 3848 3078 3851
rect 3048 3703 3050 3707
rect 3054 3703 3057 3707
rect 3062 3703 3064 3707
rect 3094 3572 3097 3748
rect 3110 3712 3113 3968
rect 3114 3668 3118 3671
rect 3102 3652 3105 3668
rect 3048 3503 3050 3507
rect 3054 3503 3057 3507
rect 3062 3503 3064 3507
rect 3086 3461 3089 3468
rect 3082 3458 3089 3461
rect 3098 3458 3102 3461
rect 3094 3392 3097 3428
rect 3118 3381 3121 3488
rect 3114 3378 3121 3381
rect 3048 3303 3050 3307
rect 3054 3303 3057 3307
rect 3062 3303 3064 3307
rect 3030 3092 3033 3118
rect 3048 3103 3050 3107
rect 3054 3103 3057 3107
rect 3062 3103 3064 3107
rect 3022 2968 3030 2971
rect 3048 2903 3050 2907
rect 3054 2903 3057 2907
rect 3062 2903 3064 2907
rect 2990 2462 2993 2468
rect 2974 2352 2977 2388
rect 2982 2332 2985 2348
rect 2998 2322 3001 2418
rect 2974 2132 2977 2148
rect 2994 1858 2998 1861
rect 2970 1748 2977 1751
rect 2994 1748 2998 1751
rect 2974 1732 2977 1748
rect 3006 1732 3009 2898
rect 3070 2862 3073 3318
rect 3102 3171 3105 3298
rect 3110 3282 3113 3288
rect 3102 3168 3110 3171
rect 3110 2932 3113 3068
rect 3078 2882 3081 2928
rect 3048 2703 3050 2707
rect 3054 2703 3057 2707
rect 3062 2703 3064 2707
rect 3086 2692 3089 2718
rect 2918 1672 2921 1678
rect 2926 1672 2929 1678
rect 2866 1628 2873 1631
rect 2870 1612 2873 1628
rect 2842 1568 2846 1571
rect 2854 1482 2857 1558
rect 2862 1548 2870 1551
rect 2882 1548 2886 1551
rect 2862 1542 2865 1548
rect 2878 1502 2881 1548
rect 2894 1542 2897 1598
rect 2906 1538 2910 1541
rect 2862 1492 2865 1498
rect 2870 1482 2873 1488
rect 2834 1478 2838 1481
rect 2846 1412 2849 1478
rect 2878 1461 2881 1498
rect 2878 1458 2886 1461
rect 2842 1328 2849 1331
rect 2846 1322 2849 1328
rect 2862 1311 2865 1378
rect 2858 1308 2865 1311
rect 2830 1102 2833 1308
rect 2838 1242 2841 1278
rect 2862 1252 2865 1278
rect 2830 1072 2833 1078
rect 2758 898 2769 901
rect 2758 472 2761 888
rect 2766 862 2769 898
rect 2766 652 2769 788
rect 2774 592 2777 688
rect 2782 661 2785 958
rect 2798 948 2806 951
rect 2790 752 2793 948
rect 2798 922 2801 948
rect 2814 941 2817 1068
rect 2810 938 2817 941
rect 2798 742 2801 748
rect 2806 722 2809 938
rect 2822 702 2825 788
rect 2782 658 2790 661
rect 2810 658 2814 661
rect 2790 622 2793 658
rect 2790 522 2793 618
rect 2734 342 2737 408
rect 2750 252 2753 358
rect 2766 322 2769 338
rect 2766 282 2769 288
rect 2758 232 2761 278
rect 2426 138 2430 141
rect 2422 92 2425 98
rect 2462 92 2465 138
rect 2274 68 2278 71
rect 1506 58 1510 61
rect 1810 58 1814 61
rect 2062 52 2065 68
rect 2238 52 2241 68
rect 2286 52 2289 78
rect 2398 72 2401 78
rect 2510 72 2513 138
rect 2594 128 2598 131
rect 2610 118 2614 121
rect 2622 81 2625 228
rect 2630 122 2633 128
rect 2646 102 2649 128
rect 2726 102 2729 218
rect 2774 202 2777 388
rect 2782 322 2785 458
rect 2790 202 2793 438
rect 2798 262 2801 528
rect 2806 462 2809 548
rect 2822 512 2825 698
rect 2830 622 2833 918
rect 2838 702 2841 1158
rect 2846 862 2849 1248
rect 2858 1168 2862 1171
rect 2862 942 2865 988
rect 2854 932 2857 938
rect 2854 862 2857 878
rect 2862 852 2865 858
rect 2862 792 2865 818
rect 2822 472 2825 508
rect 2806 452 2809 458
rect 2822 362 2825 368
rect 2830 352 2833 588
rect 2846 362 2849 768
rect 2862 742 2865 788
rect 2870 572 2873 1378
rect 2878 1192 2881 1438
rect 2894 1322 2897 1358
rect 2902 1352 2905 1528
rect 2934 1402 2937 1678
rect 2982 1662 2985 1698
rect 2966 1442 2969 1648
rect 2998 1472 3001 1538
rect 2902 1262 2905 1348
rect 2922 1328 2926 1331
rect 2918 1298 2926 1301
rect 2918 1282 2921 1298
rect 2890 1258 2894 1261
rect 2914 1258 2918 1261
rect 2926 1252 2929 1268
rect 2890 1248 2894 1251
rect 2886 1232 2889 1248
rect 2878 1022 2881 1168
rect 2902 1092 2905 1098
rect 2886 951 2889 988
rect 2886 948 2894 951
rect 2910 942 2913 1218
rect 2934 1162 2937 1338
rect 2926 942 2929 1128
rect 2934 972 2937 1118
rect 2942 1092 2945 1358
rect 2950 1222 2953 1338
rect 2966 1292 2969 1368
rect 2974 1302 2977 1368
rect 2970 1288 2974 1291
rect 2942 1042 2945 1088
rect 2958 1072 2961 1118
rect 2974 1002 2977 1258
rect 2990 1132 2993 1368
rect 2998 1162 3001 1168
rect 3006 1152 3009 1328
rect 3014 1202 3017 2588
rect 3038 2222 3041 2688
rect 3118 2672 3121 3058
rect 3126 3042 3129 3328
rect 3134 3132 3137 3398
rect 3142 3062 3145 3458
rect 3150 3171 3153 3378
rect 3158 3362 3161 4188
rect 3262 4082 3265 4328
rect 3270 4298 3278 4301
rect 3270 3992 3273 4298
rect 3226 3938 3230 3941
rect 3166 3462 3169 3518
rect 3166 3362 3169 3388
rect 3150 3168 3158 3171
rect 3154 3078 3158 3081
rect 3166 3052 3169 3318
rect 3174 3182 3177 3808
rect 3190 3671 3193 3718
rect 3186 3668 3193 3671
rect 3186 3378 3190 3381
rect 3198 3362 3201 3918
rect 3230 3782 3233 3938
rect 3302 3862 3305 4128
rect 3294 3832 3297 3858
rect 3210 3668 3217 3671
rect 3226 3668 3233 3671
rect 3214 3662 3217 3668
rect 3214 3462 3217 3618
rect 3206 3062 3209 3318
rect 3230 3242 3233 3668
rect 3278 3362 3281 3788
rect 3326 3572 3329 4208
rect 3358 4102 3361 4338
rect 3422 4242 3425 4358
rect 3494 4342 3497 4368
rect 3482 4338 3486 4341
rect 3494 4292 3497 4328
rect 3550 4312 3553 4348
rect 3654 4312 3657 4348
rect 3686 4322 3689 4338
rect 3678 4302 3681 4318
rect 3670 4262 3673 4298
rect 3568 4203 3570 4207
rect 3574 4203 3577 4207
rect 3582 4203 3584 4207
rect 3430 4072 3433 4138
rect 3622 4012 3625 4228
rect 3694 4172 3697 4348
rect 3702 4252 3705 4328
rect 3714 4308 3718 4311
rect 3742 4272 3745 4298
rect 3750 4262 3753 4298
rect 3730 4258 3734 4261
rect 3758 4222 3761 4398
rect 3766 4262 3769 4368
rect 3798 4282 3801 4348
rect 3774 4258 3782 4261
rect 3798 4261 3801 4268
rect 3794 4258 3801 4261
rect 3710 4218 3718 4221
rect 3662 4082 3665 4158
rect 3568 4003 3570 4007
rect 3574 4003 3577 4007
rect 3582 4003 3584 4007
rect 3338 3758 3342 3761
rect 3178 3058 3185 3061
rect 3182 3032 3185 3058
rect 3246 2962 3249 3128
rect 3254 3112 3257 3338
rect 3266 3268 3270 3271
rect 3048 2503 3050 2507
rect 3054 2503 3057 2507
rect 3062 2503 3064 2507
rect 3048 2303 3050 2307
rect 3054 2303 3057 2307
rect 3062 2303 3064 2307
rect 3070 2252 3073 2498
rect 3126 2462 3129 2698
rect 3134 2462 3137 2488
rect 3078 2312 3081 2318
rect 3118 2252 3121 2298
rect 3030 2142 3033 2148
rect 3026 1968 3030 1971
rect 3038 1962 3041 2158
rect 3110 2131 3113 2138
rect 3106 2128 3113 2131
rect 3086 2122 3089 2128
rect 3094 2112 3097 2128
rect 3048 2103 3050 2107
rect 3054 2103 3057 2107
rect 3062 2103 3064 2107
rect 3074 2058 3081 2061
rect 3078 2042 3081 2058
rect 3038 1881 3041 1958
rect 3048 1903 3050 1907
rect 3054 1903 3057 1907
rect 3062 1903 3064 1907
rect 3038 1878 3046 1881
rect 3014 1142 3017 1168
rect 2990 1121 2993 1128
rect 2986 1118 2993 1121
rect 2998 1112 3001 1118
rect 2998 1072 3001 1078
rect 3014 1072 3017 1138
rect 3006 1062 3009 1068
rect 2990 1038 2998 1041
rect 2946 998 2950 1001
rect 2974 952 2977 968
rect 2966 941 2969 948
rect 2962 938 2969 941
rect 2878 862 2881 868
rect 2886 742 2889 898
rect 2926 772 2929 938
rect 2970 868 2974 871
rect 2958 862 2961 868
rect 2934 792 2937 808
rect 2934 752 2937 758
rect 2938 738 2942 741
rect 2942 728 2950 731
rect 2934 722 2937 728
rect 2918 682 2921 688
rect 2862 471 2865 508
rect 2858 468 2865 471
rect 2862 462 2865 468
rect 2818 338 2822 341
rect 2810 318 2814 321
rect 2838 318 2846 321
rect 2838 282 2841 318
rect 2742 152 2745 168
rect 2774 152 2777 198
rect 2862 192 2865 208
rect 2870 192 2873 568
rect 2902 562 2905 578
rect 2878 548 2886 551
rect 2878 462 2881 548
rect 2902 471 2905 558
rect 2930 518 2934 521
rect 2898 468 2905 471
rect 2942 452 2945 728
rect 2958 622 2961 828
rect 2982 792 2985 998
rect 2990 922 2993 1038
rect 2998 951 3001 998
rect 2998 948 3006 951
rect 3002 918 3006 921
rect 2966 712 2969 758
rect 2974 752 2977 758
rect 2990 728 2998 731
rect 2954 548 2958 551
rect 2958 272 2961 468
rect 2966 382 2969 708
rect 2990 592 2993 728
rect 3002 678 3009 681
rect 3006 652 3009 678
rect 3014 562 3017 868
rect 3022 762 3025 1708
rect 3030 1682 3033 1838
rect 3038 1702 3041 1748
rect 3048 1703 3050 1707
rect 3054 1703 3057 1707
rect 3062 1703 3064 1707
rect 3030 1602 3033 1628
rect 3070 1572 3073 1958
rect 3134 1792 3137 2458
rect 3142 2422 3145 2678
rect 3150 2012 3153 2788
rect 3158 1972 3161 2578
rect 3166 2472 3169 2478
rect 3166 2272 3169 2278
rect 3166 2142 3169 2158
rect 3166 2132 3169 2138
rect 3158 1942 3161 1968
rect 3162 1848 3166 1851
rect 3102 1662 3105 1668
rect 3078 1528 3086 1531
rect 3048 1503 3050 1507
rect 3054 1503 3057 1507
rect 3062 1503 3064 1507
rect 3062 1471 3065 1488
rect 3058 1468 3065 1471
rect 3078 1452 3081 1528
rect 3110 1512 3113 1678
rect 3110 1472 3113 1508
rect 3090 1468 3094 1471
rect 3082 1438 3086 1441
rect 3066 1348 3070 1351
rect 3030 1072 3033 1278
rect 3038 1242 3041 1338
rect 3078 1312 3081 1418
rect 3048 1303 3050 1307
rect 3054 1303 3057 1307
rect 3062 1303 3064 1307
rect 3062 1251 3065 1258
rect 3078 1252 3081 1278
rect 3062 1248 3070 1251
rect 3054 1232 3057 1248
rect 3086 1222 3089 1378
rect 3110 1332 3113 1468
rect 3118 1462 3121 1658
rect 3126 1452 3129 1458
rect 3134 1412 3137 1528
rect 3094 1302 3097 1318
rect 3102 1251 3105 1278
rect 3102 1248 3110 1251
rect 3038 1152 3041 1178
rect 3102 1161 3105 1198
rect 3098 1158 3105 1161
rect 3110 1162 3113 1168
rect 3038 1112 3041 1128
rect 3048 1103 3050 1107
rect 3054 1103 3057 1107
rect 3062 1103 3064 1107
rect 3034 1058 3038 1061
rect 3046 922 3049 938
rect 3048 903 3050 907
rect 3054 903 3057 907
rect 3062 903 3064 907
rect 3070 892 3073 1098
rect 3086 962 3089 968
rect 3078 952 3081 958
rect 3102 931 3105 1138
rect 3110 1112 3113 1148
rect 3118 1062 3121 1408
rect 3098 928 3105 931
rect 3106 918 3110 921
rect 3030 872 3033 878
rect 3038 871 3041 878
rect 3038 868 3046 871
rect 3066 848 3070 851
rect 3038 712 3041 728
rect 3048 703 3050 707
rect 3054 703 3057 707
rect 3062 703 3064 707
rect 3070 652 3073 678
rect 3022 442 3025 638
rect 3048 503 3050 507
rect 3054 503 3057 507
rect 3062 503 3064 507
rect 2966 252 2969 378
rect 3022 362 3025 438
rect 3038 432 3041 488
rect 3070 452 3073 548
rect 3086 502 3089 578
rect 3082 398 3086 401
rect 2930 248 2934 251
rect 2754 148 2758 151
rect 2790 112 2793 178
rect 2806 141 2809 148
rect 2802 138 2809 141
rect 2778 108 2782 111
rect 2622 78 2630 81
rect 2522 68 2529 71
rect 2570 68 2574 71
rect 2814 71 2817 98
rect 2814 68 2822 71
rect 2842 68 2846 71
rect 2526 62 2529 68
rect 2870 52 2873 188
rect 2926 101 2929 158
rect 2942 142 2945 228
rect 2950 172 2953 238
rect 2974 192 2977 238
rect 2982 232 2985 338
rect 2978 168 2982 171
rect 2950 142 2953 168
rect 2958 102 2961 168
rect 2926 98 2934 101
rect 2974 51 2977 148
rect 3014 142 3017 358
rect 3026 328 3030 331
rect 3094 322 3097 918
rect 3102 602 3105 898
rect 3110 862 3113 868
rect 3110 542 3113 848
rect 3118 732 3121 1048
rect 3126 1012 3129 1328
rect 3134 1142 3137 1378
rect 3142 1292 3145 1298
rect 3142 1262 3145 1268
rect 3142 1162 3145 1168
rect 3150 1152 3153 1798
rect 3166 1742 3169 1758
rect 3166 1531 3169 1698
rect 3174 1542 3177 2658
rect 3198 2552 3201 2688
rect 3206 2648 3214 2651
rect 3206 2522 3209 2648
rect 3246 2542 3249 2918
rect 3242 2498 3246 2501
rect 3238 2372 3241 2408
rect 3182 1992 3185 2148
rect 3190 1992 3193 2008
rect 3198 1952 3201 1988
rect 3182 1672 3185 1688
rect 3190 1592 3193 1748
rect 3198 1742 3201 1848
rect 3198 1652 3201 1738
rect 3206 1672 3209 1678
rect 3186 1548 3190 1551
rect 3166 1528 3177 1531
rect 3158 1412 3161 1418
rect 3166 1392 3169 1418
rect 3174 1392 3177 1528
rect 3198 1522 3201 1648
rect 3214 1492 3217 2308
rect 3222 2242 3225 2258
rect 3222 2132 3225 2138
rect 3230 2092 3233 2148
rect 3246 2142 3249 2148
rect 3254 2112 3257 3098
rect 3262 2662 3265 2708
rect 3270 2492 3273 3208
rect 3278 2912 3281 3268
rect 3286 3182 3289 3338
rect 3294 3202 3297 3538
rect 3338 3518 3342 3521
rect 3310 3332 3313 3518
rect 3350 3462 3353 3478
rect 3318 3402 3321 3408
rect 3322 3328 3326 3331
rect 3322 3318 3326 3321
rect 3302 3272 3305 3278
rect 3270 2442 3273 2488
rect 3262 2392 3265 2398
rect 3286 2232 3289 2988
rect 3294 2382 3297 3118
rect 3302 2882 3305 2888
rect 3310 2582 3313 3268
rect 3318 3052 3321 3128
rect 3342 2892 3345 3188
rect 3358 3072 3361 3578
rect 3382 3562 3385 3568
rect 3366 3442 3369 3458
rect 3370 3358 3374 3361
rect 3398 3272 3401 3708
rect 3406 3602 3409 3978
rect 3610 3948 3614 3951
rect 3622 3942 3625 4008
rect 3430 3852 3433 3938
rect 3590 3902 3593 3928
rect 3494 3692 3497 3878
rect 3518 3842 3521 3858
rect 3710 3842 3713 4218
rect 3726 4028 3734 4031
rect 3726 3952 3729 4028
rect 3806 4002 3809 4318
rect 3814 4302 3817 4308
rect 3814 4102 3817 4258
rect 3830 4232 3833 4398
rect 3918 4362 3921 4368
rect 3790 3872 3793 3978
rect 3814 3942 3817 4098
rect 3838 3932 3841 4348
rect 3934 4342 3937 4348
rect 3858 4258 3862 4261
rect 3902 4072 3905 4288
rect 3918 4132 3921 4228
rect 3942 4112 3945 4388
rect 3974 4342 3977 4348
rect 3958 4322 3961 4338
rect 3990 4272 3993 4318
rect 3902 3962 3905 4068
rect 3814 3892 3817 3918
rect 3568 3803 3570 3807
rect 3574 3803 3577 3807
rect 3582 3803 3584 3807
rect 3854 3782 3857 3958
rect 3866 3948 3870 3951
rect 3870 3852 3873 3908
rect 3430 3562 3433 3568
rect 3462 3452 3465 3518
rect 3442 3348 3446 3351
rect 3350 2502 3353 2578
rect 3270 2142 3273 2188
rect 3278 2091 3281 2178
rect 3358 2162 3361 2778
rect 3366 2382 3369 3038
rect 3390 2592 3393 2688
rect 3406 2671 3409 3018
rect 3402 2668 3409 2671
rect 3430 2622 3433 3278
rect 3438 2692 3441 3228
rect 3438 2672 3441 2688
rect 3374 2572 3377 2578
rect 3366 2322 3369 2328
rect 3374 2252 3377 2368
rect 3274 2088 3281 2091
rect 3246 1942 3249 1958
rect 3326 1782 3329 2108
rect 3374 2052 3377 2118
rect 3382 2092 3385 2568
rect 3390 2222 3393 2588
rect 3402 2548 3406 2551
rect 3422 2542 3425 2558
rect 3430 2541 3433 2618
rect 3430 2538 3438 2541
rect 3414 2412 3417 2458
rect 3402 2348 3409 2351
rect 3406 2322 3409 2348
rect 3414 2342 3417 2368
rect 3430 2242 3433 2338
rect 3390 2192 3393 2218
rect 3438 2172 3441 2278
rect 3454 2262 3457 3228
rect 3470 2542 3473 3578
rect 3486 3552 3489 3688
rect 3478 3372 3481 3378
rect 3486 3022 3489 3058
rect 3462 2481 3465 2488
rect 3462 2478 3470 2481
rect 3470 2262 3473 2268
rect 3478 2242 3481 2978
rect 3486 2462 3489 2478
rect 3494 2272 3497 2888
rect 3494 2152 3497 2178
rect 3502 2162 3505 3488
rect 3534 3332 3537 3348
rect 3510 2172 3513 2758
rect 3534 2532 3537 2918
rect 3510 2162 3513 2168
rect 3402 2148 3406 2151
rect 3358 1972 3361 2018
rect 3382 1982 3385 2088
rect 3518 1972 3521 1988
rect 3514 1968 3518 1971
rect 3426 1938 3430 1941
rect 3366 1792 3369 1798
rect 3238 1722 3241 1738
rect 3166 1202 3169 1388
rect 3166 1122 3169 1138
rect 3174 1062 3177 1318
rect 3182 1162 3185 1438
rect 3206 1412 3209 1468
rect 3214 1392 3217 1428
rect 3202 1348 3206 1351
rect 3190 1342 3193 1348
rect 3222 1342 3225 1618
rect 3230 1462 3233 1468
rect 3218 1328 3222 1331
rect 3206 1242 3209 1328
rect 3214 1202 3217 1218
rect 3222 1192 3225 1318
rect 3230 1262 3233 1268
rect 3210 1188 3217 1191
rect 3182 1082 3185 1158
rect 3190 1062 3193 1088
rect 3158 1052 3161 1058
rect 3194 1038 3198 1041
rect 3134 892 3137 1028
rect 3166 942 3169 988
rect 3182 952 3185 968
rect 3206 952 3209 1118
rect 3174 871 3177 938
rect 3182 912 3185 948
rect 3170 868 3177 871
rect 3202 868 3206 871
rect 3142 742 3145 868
rect 3214 862 3217 1188
rect 3222 1042 3225 1148
rect 3238 1062 3241 1408
rect 3270 1382 3273 1678
rect 3278 1552 3281 1748
rect 3294 1742 3297 1748
rect 3350 1572 3353 1768
rect 3358 1662 3361 1668
rect 3390 1662 3393 1798
rect 3494 1682 3497 1828
rect 3482 1678 3486 1681
rect 3278 1432 3281 1458
rect 3278 1382 3281 1428
rect 3278 1322 3281 1338
rect 3286 1322 3289 1558
rect 3302 1462 3305 1548
rect 3334 1342 3337 1508
rect 3350 1462 3353 1568
rect 3402 1548 3409 1551
rect 3238 1022 3241 1038
rect 3222 942 3225 948
rect 3222 892 3225 898
rect 3134 712 3137 728
rect 3118 542 3121 548
rect 3102 422 3105 538
rect 3126 452 3129 648
rect 3134 582 3137 698
rect 3150 352 3153 858
rect 3158 782 3161 808
rect 3166 692 3169 798
rect 3198 752 3201 838
rect 3230 802 3233 998
rect 3238 932 3241 938
rect 3238 922 3241 928
rect 3214 752 3217 758
rect 3238 712 3241 898
rect 3246 772 3249 1298
rect 3254 1232 3257 1288
rect 3274 1268 3281 1271
rect 3254 1102 3257 1198
rect 3262 1082 3265 1168
rect 3270 1132 3273 1138
rect 3278 1122 3281 1268
rect 3286 1142 3289 1158
rect 3270 1032 3273 1108
rect 3294 1072 3297 1308
rect 3302 1268 3310 1271
rect 3302 1262 3305 1268
rect 3306 1138 3313 1141
rect 3310 1132 3313 1138
rect 3318 1132 3321 1268
rect 3326 1142 3329 1168
rect 3278 1012 3281 1018
rect 3254 872 3257 978
rect 3262 932 3265 968
rect 3254 762 3257 868
rect 3262 712 3265 928
rect 3274 888 3278 891
rect 3302 792 3305 868
rect 3310 842 3313 1078
rect 3330 1068 3334 1071
rect 3334 992 3337 1018
rect 3334 972 3337 978
rect 3342 941 3345 1198
rect 3350 1072 3353 1318
rect 3358 1202 3361 1228
rect 3366 1212 3369 1508
rect 3374 1372 3377 1548
rect 3406 1522 3409 1548
rect 3386 1458 3390 1461
rect 3358 1162 3361 1168
rect 3358 1052 3361 1068
rect 3350 958 3358 961
rect 3350 952 3353 958
rect 3322 938 3329 941
rect 3342 938 3350 941
rect 3326 802 3329 938
rect 3350 852 3353 878
rect 3166 681 3169 688
rect 3166 678 3174 681
rect 3182 622 3185 648
rect 3158 362 3161 548
rect 3182 522 3185 618
rect 3198 562 3201 708
rect 3266 648 3270 651
rect 3278 641 3281 748
rect 3294 702 3297 748
rect 3334 722 3337 798
rect 3358 692 3361 948
rect 3374 922 3377 1078
rect 3382 1051 3385 1458
rect 3382 1048 3390 1051
rect 3382 882 3385 998
rect 3390 992 3393 998
rect 3390 932 3393 968
rect 3398 932 3401 1258
rect 3406 962 3409 1518
rect 3414 1512 3417 1678
rect 3414 1232 3417 1508
rect 3454 1362 3457 1618
rect 3486 1392 3489 1578
rect 3426 1228 3430 1231
rect 3454 1161 3457 1358
rect 3450 1158 3457 1161
rect 3414 1132 3417 1138
rect 3438 1132 3441 1158
rect 3390 852 3393 868
rect 3398 762 3401 848
rect 3378 748 3385 751
rect 3366 732 3369 748
rect 3382 722 3385 748
rect 3358 672 3361 688
rect 3278 638 3286 641
rect 3238 542 3241 588
rect 3390 572 3393 758
rect 3406 652 3409 828
rect 3414 762 3417 1008
rect 3430 972 3433 1068
rect 3438 932 3441 978
rect 3422 928 3430 931
rect 3422 842 3425 928
rect 3446 892 3449 1138
rect 3454 1112 3457 1118
rect 3446 882 3449 888
rect 3422 822 3425 838
rect 3454 832 3457 1048
rect 3438 762 3441 778
rect 3426 738 3430 741
rect 3438 722 3441 748
rect 3230 538 3238 541
rect 3174 482 3177 518
rect 3206 402 3209 518
rect 3230 452 3233 538
rect 3150 338 3153 348
rect 3174 312 3177 348
rect 3048 303 3050 307
rect 3054 303 3057 307
rect 3062 303 3064 307
rect 3174 262 3177 308
rect 3194 258 3198 261
rect 3206 252 3209 258
rect 3078 222 3081 248
rect 3122 168 3126 171
rect 3030 132 3033 158
rect 3038 142 3041 158
rect 3038 112 3041 138
rect 3110 122 3113 158
rect 3048 103 3050 107
rect 3054 103 3057 107
rect 3062 103 3064 107
rect 3150 92 3153 188
rect 2990 72 2993 88
rect 2998 72 3001 78
rect 3022 62 3025 78
rect 3078 62 3081 78
rect 3050 58 3054 61
rect 3110 52 3113 58
rect 3118 52 3121 68
rect 3150 52 3153 88
rect 3166 82 3169 118
rect 3174 112 3177 228
rect 3214 142 3217 188
rect 3222 142 3225 338
rect 3262 312 3265 558
rect 3310 492 3313 548
rect 3402 538 3406 541
rect 3422 512 3425 548
rect 3430 532 3433 668
rect 3298 448 3302 451
rect 3298 338 3302 341
rect 3230 202 3233 268
rect 3230 171 3233 198
rect 3230 168 3238 171
rect 3254 142 3257 158
rect 3262 112 3265 248
rect 3278 162 3281 178
rect 3254 82 3257 98
rect 3162 78 3166 81
rect 3246 52 3249 68
rect 3270 52 3273 128
rect 3278 92 3281 118
rect 3286 72 3289 338
rect 3298 298 3302 301
rect 3350 262 3353 468
rect 3358 462 3361 508
rect 3398 332 3401 338
rect 3406 332 3409 438
rect 3454 392 3457 828
rect 3462 752 3465 1348
rect 3478 1292 3481 1318
rect 3478 1262 3481 1278
rect 3470 1072 3473 1258
rect 3478 1142 3481 1248
rect 3486 1192 3489 1298
rect 3486 1162 3489 1178
rect 3478 1022 3481 1038
rect 3478 931 3481 968
rect 3474 928 3481 931
rect 3478 812 3481 858
rect 3462 732 3465 748
rect 3478 722 3481 728
rect 3470 502 3473 648
rect 3486 512 3489 1038
rect 3494 532 3497 1588
rect 3502 1552 3505 1718
rect 3510 1592 3513 1728
rect 3526 1592 3529 2508
rect 3542 2362 3545 3588
rect 3550 3072 3553 3658
rect 3568 3603 3570 3607
rect 3574 3603 3577 3607
rect 3582 3603 3584 3607
rect 3568 3403 3570 3407
rect 3574 3403 3577 3407
rect 3582 3403 3584 3407
rect 3568 3203 3570 3207
rect 3574 3203 3577 3207
rect 3582 3203 3584 3207
rect 3568 3003 3570 3007
rect 3574 3003 3577 3007
rect 3582 3003 3584 3007
rect 3568 2803 3570 2807
rect 3574 2803 3577 2807
rect 3582 2803 3584 2807
rect 3568 2603 3570 2607
rect 3574 2603 3577 2607
rect 3582 2603 3584 2607
rect 3558 2332 3561 2528
rect 3590 2522 3593 3608
rect 3742 3552 3745 3658
rect 3614 3452 3617 3518
rect 3590 2472 3593 2498
rect 3598 2452 3601 3428
rect 3702 3261 3705 3308
rect 3698 3258 3705 3261
rect 3638 3111 3641 3118
rect 3638 3108 3646 3111
rect 3638 2622 3641 3108
rect 3670 2861 3673 3138
rect 3666 2858 3673 2861
rect 3654 2552 3657 2558
rect 3626 2518 3630 2521
rect 3642 2468 3646 2471
rect 3568 2403 3570 2407
rect 3574 2403 3577 2407
rect 3582 2403 3584 2407
rect 3590 2352 3593 2408
rect 3606 2341 3609 2348
rect 3602 2338 3609 2341
rect 3568 2203 3570 2207
rect 3574 2203 3577 2207
rect 3582 2203 3584 2207
rect 3550 2122 3553 2138
rect 3646 2112 3649 2128
rect 3582 2032 3585 2048
rect 3568 2003 3570 2007
rect 3574 2003 3577 2007
rect 3582 2003 3584 2007
rect 3630 2002 3633 2108
rect 3630 1912 3633 1998
rect 3558 1762 3561 1808
rect 3568 1803 3570 1807
rect 3574 1803 3577 1807
rect 3582 1803 3584 1807
rect 3630 1752 3633 1758
rect 3542 1662 3545 1738
rect 3566 1732 3569 1748
rect 3550 1682 3553 1698
rect 3568 1603 3570 1607
rect 3574 1603 3577 1607
rect 3582 1603 3584 1607
rect 3610 1548 3614 1551
rect 3526 1542 3529 1548
rect 3502 1312 3505 1528
rect 3606 1462 3609 1468
rect 3518 1302 3521 1408
rect 3568 1403 3570 1407
rect 3574 1403 3577 1407
rect 3582 1403 3584 1407
rect 3614 1372 3617 1448
rect 3526 1332 3529 1348
rect 3502 1072 3505 1248
rect 3510 1222 3513 1298
rect 3550 1262 3553 1268
rect 3582 1252 3585 1358
rect 3598 1332 3601 1348
rect 3590 1322 3593 1328
rect 3542 1232 3545 1248
rect 3568 1203 3570 1207
rect 3574 1203 3577 1207
rect 3582 1203 3584 1207
rect 3542 1162 3545 1198
rect 3558 1132 3561 1188
rect 3590 1142 3593 1278
rect 3598 1252 3601 1328
rect 3510 1081 3513 1108
rect 3526 1102 3529 1118
rect 3510 1078 3518 1081
rect 3502 1042 3505 1048
rect 3502 832 3505 938
rect 3510 822 3513 1028
rect 3534 1012 3537 1068
rect 3518 892 3521 908
rect 3542 892 3545 1098
rect 3550 982 3553 1128
rect 3558 1032 3561 1128
rect 3570 1068 3574 1071
rect 3582 1042 3585 1068
rect 3590 1062 3593 1138
rect 3568 1003 3570 1007
rect 3574 1003 3577 1007
rect 3582 1003 3584 1007
rect 3550 922 3553 938
rect 3526 872 3529 878
rect 3546 828 3553 831
rect 3502 772 3505 818
rect 3510 808 3518 811
rect 3522 808 3526 811
rect 3502 712 3505 758
rect 3422 332 3425 338
rect 3386 278 3390 281
rect 3446 281 3449 368
rect 3446 278 3454 281
rect 3314 238 3321 241
rect 3318 222 3321 238
rect 3318 162 3321 218
rect 3366 122 3369 248
rect 3438 142 3441 268
rect 3462 182 3465 318
rect 3470 202 3473 498
rect 3494 492 3497 528
rect 3502 422 3505 538
rect 3510 482 3513 808
rect 3550 802 3553 828
rect 3558 742 3561 978
rect 3566 942 3569 948
rect 3574 842 3577 968
rect 3590 861 3593 878
rect 3586 858 3593 861
rect 3568 803 3570 807
rect 3574 803 3577 807
rect 3582 803 3584 807
rect 3570 738 3574 741
rect 3598 682 3601 1248
rect 3614 1202 3617 1368
rect 3610 1128 3617 1131
rect 3614 1082 3617 1128
rect 3606 1042 3609 1068
rect 3614 922 3617 928
rect 3622 922 3625 1268
rect 3630 1222 3633 1578
rect 3650 1468 3654 1471
rect 3654 1292 3657 1318
rect 3638 1222 3641 1238
rect 3630 1132 3633 1148
rect 3630 1082 3633 1088
rect 3638 1072 3641 1218
rect 3646 1212 3649 1228
rect 3654 1192 3657 1248
rect 3662 1182 3665 2838
rect 3670 2282 3673 2698
rect 3678 2682 3681 3018
rect 3686 2162 3689 2878
rect 3694 2632 3697 2968
rect 3698 2518 3705 2521
rect 3702 2502 3705 2518
rect 3670 2062 3673 2128
rect 3670 1842 3673 2058
rect 3686 2002 3689 2048
rect 3678 1972 3681 1978
rect 3694 1892 3697 2488
rect 3710 2202 3713 3188
rect 3742 2582 3745 2828
rect 3774 2732 3777 3598
rect 3790 3482 3793 3778
rect 3726 2542 3729 2568
rect 3742 2562 3745 2578
rect 3734 2512 3737 2538
rect 3750 2172 3753 2388
rect 3758 2262 3761 2268
rect 3782 2182 3785 3348
rect 3798 3062 3801 3718
rect 3886 3632 3889 3948
rect 3894 3782 3897 3958
rect 3910 3772 3913 4078
rect 3966 3942 3969 4198
rect 3982 4032 3985 4148
rect 3982 3951 3985 4028
rect 3990 4021 3993 4268
rect 3998 4042 4001 4388
rect 4014 4261 4017 4278
rect 4010 4258 4017 4261
rect 4022 4172 4025 4388
rect 4054 4322 4057 4398
rect 4146 4358 4150 4361
rect 3990 4018 3998 4021
rect 4022 3982 4025 4168
rect 3978 3948 3985 3951
rect 3934 3872 3937 3918
rect 4046 3872 4049 4038
rect 3922 3868 3926 3871
rect 3946 3868 3950 3871
rect 3934 3752 3937 3868
rect 4054 3752 4057 4318
rect 4062 4152 4065 4358
rect 4080 4303 4082 4307
rect 4086 4303 4089 4307
rect 4094 4303 4096 4307
rect 4102 4292 4105 4328
rect 4062 4012 4065 4148
rect 4102 4112 4105 4208
rect 4080 4103 4082 4107
rect 4086 4103 4089 4107
rect 4094 4103 4096 4107
rect 4110 4092 4113 4338
rect 4126 4331 4129 4338
rect 4122 4328 4129 4331
rect 4126 4232 4129 4328
rect 4122 4158 4126 4161
rect 4134 4092 4137 4238
rect 4142 4212 4145 4318
rect 4158 4172 4161 4398
rect 4142 4162 4145 4168
rect 4070 3762 4073 3908
rect 4080 3903 4082 3907
rect 4086 3903 4089 3907
rect 4094 3903 4096 3907
rect 4080 3703 4082 3707
rect 4086 3703 4089 3707
rect 4094 3703 4096 3707
rect 4118 3702 4121 4078
rect 4134 4072 4137 4088
rect 4142 4072 4145 4078
rect 4166 4012 4169 4348
rect 4178 4318 4182 4321
rect 4190 4252 4193 4368
rect 4214 3982 4217 4358
rect 4254 4232 4257 4398
rect 4354 4348 4358 4351
rect 4330 4338 4334 4341
rect 4302 4262 4305 4308
rect 4270 4248 4278 4251
rect 4230 3892 4233 4068
rect 4254 3962 4257 4228
rect 4270 3832 4273 4248
rect 4294 4102 4297 4248
rect 3810 3568 3814 3571
rect 3886 3522 3889 3568
rect 3806 2898 3814 2901
rect 3806 2692 3809 2898
rect 3806 2672 3809 2688
rect 3830 2482 3833 3468
rect 3850 3458 3854 3461
rect 3814 2432 3817 2458
rect 3858 2348 3862 2351
rect 3838 2302 3841 2318
rect 3870 2281 3873 2288
rect 3866 2278 3873 2281
rect 3702 1992 3705 2058
rect 3750 2012 3753 2068
rect 3758 2042 3761 2048
rect 3722 1968 3726 1971
rect 3678 1602 3681 1668
rect 3686 1572 3689 1758
rect 3694 1672 3697 1878
rect 3702 1672 3705 1968
rect 3714 1948 3718 1951
rect 3750 1892 3753 2008
rect 3766 1712 3769 2158
rect 3790 2142 3793 2148
rect 3774 1762 3777 2058
rect 3782 2052 3785 2138
rect 3790 1922 3793 2138
rect 3802 2048 3806 2051
rect 3814 2042 3817 2068
rect 3798 2012 3801 2018
rect 3814 1782 3817 2038
rect 3822 1932 3825 1958
rect 3830 1952 3833 2148
rect 3838 2122 3841 2228
rect 3838 1942 3841 1958
rect 3846 1932 3849 2038
rect 3854 1962 3857 2118
rect 3822 1772 3825 1928
rect 3846 1822 3849 1928
rect 3862 1842 3865 2128
rect 3870 2112 3873 2218
rect 3878 2072 3881 3158
rect 3882 2048 3886 2051
rect 3894 1952 3897 1958
rect 3710 1682 3713 1688
rect 3698 1638 3702 1641
rect 3670 1302 3673 1378
rect 3694 1312 3697 1458
rect 3678 1232 3681 1258
rect 3670 1112 3673 1198
rect 3670 1072 3673 1108
rect 3630 812 3633 928
rect 3638 802 3641 898
rect 3662 892 3665 1048
rect 3686 972 3689 1298
rect 3694 1258 3702 1261
rect 3694 1242 3697 1258
rect 3694 1032 3697 1038
rect 3670 932 3673 958
rect 3650 848 3657 851
rect 3654 782 3657 848
rect 3618 748 3625 751
rect 3606 712 3609 748
rect 3622 732 3625 748
rect 3658 678 3662 681
rect 3654 672 3657 678
rect 3678 662 3681 888
rect 3694 822 3697 938
rect 3702 842 3705 1048
rect 3710 932 3713 938
rect 3622 632 3625 638
rect 3568 603 3570 607
rect 3574 603 3577 607
rect 3582 603 3584 607
rect 3598 562 3601 578
rect 3622 562 3625 628
rect 3662 622 3665 648
rect 3522 438 3529 441
rect 3526 422 3529 438
rect 3568 403 3570 407
rect 3574 403 3577 407
rect 3582 403 3584 407
rect 3482 318 3486 321
rect 3502 262 3505 278
rect 3482 218 3489 221
rect 3510 221 3513 298
rect 3542 292 3545 298
rect 3550 282 3553 288
rect 3506 218 3513 221
rect 3486 212 3489 218
rect 3558 202 3561 308
rect 3568 203 3570 207
rect 3574 203 3577 207
rect 3582 203 3584 207
rect 3446 112 3449 148
rect 3462 122 3465 168
rect 3518 152 3521 178
rect 3534 131 3537 138
rect 3534 128 3542 131
rect 3558 112 3561 178
rect 3570 138 3574 141
rect 3574 112 3577 118
rect 3370 108 3374 111
rect 3582 102 3585 148
rect 3590 142 3593 308
rect 3598 132 3601 558
rect 3662 452 3665 618
rect 3686 611 3689 618
rect 3682 608 3689 611
rect 3694 581 3697 818
rect 3702 752 3705 808
rect 3718 762 3721 1578
rect 3734 1342 3737 1498
rect 3742 1192 3745 1458
rect 3766 1372 3769 1658
rect 3750 1272 3753 1278
rect 3730 1188 3734 1191
rect 3774 1182 3777 1758
rect 3838 1662 3841 1718
rect 3842 1648 3846 1651
rect 3782 1422 3785 1438
rect 3734 1072 3737 1148
rect 3766 1122 3769 1128
rect 3758 1102 3761 1118
rect 3774 1112 3777 1118
rect 3766 1092 3769 1108
rect 3778 1088 3782 1091
rect 3730 948 3737 951
rect 3734 912 3737 948
rect 3742 922 3745 1038
rect 3766 1022 3769 1078
rect 3774 1052 3777 1068
rect 3766 952 3769 1018
rect 3782 952 3785 1068
rect 3790 962 3793 1138
rect 3798 962 3801 1298
rect 3806 1082 3809 1328
rect 3806 962 3809 968
rect 3762 918 3766 921
rect 3726 872 3729 878
rect 3782 862 3785 948
rect 3790 902 3793 908
rect 3794 868 3798 871
rect 3702 592 3705 748
rect 3758 692 3761 768
rect 3774 752 3777 758
rect 3782 742 3785 858
rect 3814 842 3817 1628
rect 3870 1372 3873 1478
rect 3830 1162 3833 1168
rect 3686 578 3697 581
rect 3606 152 3609 398
rect 3650 348 3657 351
rect 3654 342 3657 348
rect 3614 312 3617 318
rect 3662 281 3665 388
rect 3670 322 3673 328
rect 3662 278 3670 281
rect 3662 272 3665 278
rect 3678 272 3681 448
rect 3686 232 3689 578
rect 3698 568 3702 571
rect 3694 432 3697 448
rect 3702 362 3705 438
rect 3698 318 3702 321
rect 3710 302 3713 568
rect 3718 362 3721 368
rect 3718 352 3721 358
rect 3710 272 3713 298
rect 3654 192 3657 218
rect 3654 142 3657 188
rect 3594 118 3598 121
rect 3606 112 3609 128
rect 3662 102 3665 188
rect 3682 158 3686 161
rect 3314 78 3318 81
rect 3430 72 3433 78
rect 3522 68 3526 71
rect 3294 52 3297 58
rect 3486 52 3489 58
rect 3598 52 3601 78
rect 3614 52 3617 88
rect 3702 62 3705 158
rect 3718 82 3721 218
rect 3726 62 3729 678
rect 3734 322 3737 548
rect 3742 482 3745 488
rect 3742 282 3745 408
rect 3734 141 3737 278
rect 3734 138 3742 141
rect 3750 81 3753 688
rect 3782 562 3785 608
rect 3758 342 3761 418
rect 3806 382 3809 698
rect 3814 492 3817 828
rect 3822 812 3825 1048
rect 3838 1012 3841 1348
rect 3878 1282 3881 1458
rect 3902 1402 3905 3558
rect 4030 3462 4033 3658
rect 4080 3503 4082 3507
rect 4086 3503 4089 3507
rect 4094 3503 4096 3507
rect 4102 3502 4105 3668
rect 4190 3652 4193 3688
rect 4262 3662 4265 3748
rect 4286 3732 4289 3928
rect 4294 3762 4297 3918
rect 3938 3458 3942 3461
rect 3918 2482 3921 2528
rect 3930 2448 3934 2451
rect 3950 2362 3953 3298
rect 3958 2652 3961 3188
rect 4050 3138 4054 3141
rect 3998 2462 4001 2768
rect 4042 2668 4049 2671
rect 4038 2482 4041 2488
rect 3998 2362 4001 2458
rect 4014 2372 4017 2408
rect 4010 2348 4014 2351
rect 3970 2338 3974 2341
rect 4022 2202 4025 2228
rect 4046 2182 4049 2668
rect 4054 2432 4057 2728
rect 4070 2412 4073 3498
rect 4102 3388 4110 3391
rect 4080 3303 4082 3307
rect 4086 3303 4089 3307
rect 4094 3303 4096 3307
rect 4102 3222 4105 3388
rect 4118 3142 4121 3268
rect 4080 3103 4082 3107
rect 4086 3103 4089 3107
rect 4094 3103 4096 3107
rect 4080 2903 4082 2907
rect 4086 2903 4089 2907
rect 4094 2903 4096 2907
rect 4080 2703 4082 2707
rect 4086 2703 4089 2707
rect 4094 2703 4096 2707
rect 4080 2503 4082 2507
rect 4086 2503 4089 2507
rect 4094 2503 4096 2507
rect 4080 2303 4082 2307
rect 4086 2303 4089 2307
rect 4094 2303 4096 2307
rect 4090 2268 4094 2271
rect 4086 2212 4089 2258
rect 4046 2022 4049 2158
rect 4080 2103 4082 2107
rect 4086 2103 4089 2107
rect 4094 2103 4096 2107
rect 3962 1958 3966 1961
rect 3966 1912 3969 1918
rect 3918 1742 3921 1748
rect 3942 1522 3945 1908
rect 3958 1872 3961 1878
rect 3974 1792 3977 2008
rect 4050 1998 4054 2001
rect 3982 1832 3985 1958
rect 4038 1932 4041 1948
rect 4022 1928 4030 1931
rect 4022 1832 4025 1928
rect 4062 1922 4065 2048
rect 3958 1672 3961 1728
rect 3954 1668 3958 1671
rect 3966 1662 3969 1668
rect 3890 1358 3894 1361
rect 3846 1252 3849 1278
rect 3854 1102 3857 1248
rect 3886 1242 3889 1258
rect 3846 1092 3849 1098
rect 3830 942 3833 948
rect 3846 902 3849 1048
rect 3854 932 3857 1098
rect 3862 1012 3865 1048
rect 3870 962 3873 1138
rect 3866 868 3870 871
rect 3846 842 3849 848
rect 3830 812 3833 838
rect 3830 802 3833 808
rect 3826 788 3830 791
rect 3822 722 3825 768
rect 3822 532 3825 548
rect 3830 452 3833 758
rect 3838 712 3841 798
rect 3846 718 3854 721
rect 3822 442 3825 448
rect 3846 412 3849 718
rect 3878 712 3881 1088
rect 3886 952 3889 958
rect 3894 931 3897 948
rect 3890 928 3897 931
rect 3894 892 3897 928
rect 3894 692 3897 718
rect 3902 692 3905 1338
rect 3910 1302 3913 1378
rect 3910 852 3913 1228
rect 3930 1168 3934 1171
rect 3918 1042 3921 1048
rect 3926 872 3929 878
rect 3934 862 3937 878
rect 3942 852 3945 1508
rect 3910 772 3913 848
rect 3950 792 3953 1548
rect 3974 1462 3977 1708
rect 3982 1632 3985 1748
rect 3990 1532 3993 1748
rect 4010 1648 4014 1651
rect 3990 1512 3993 1528
rect 3982 1442 3985 1468
rect 3962 1328 3966 1331
rect 3958 1282 3961 1318
rect 3958 982 3961 1238
rect 3966 1212 3969 1318
rect 3982 1262 3985 1438
rect 3970 1208 3977 1211
rect 3974 1202 3977 1208
rect 3966 1102 3969 1148
rect 3966 1062 3969 1098
rect 3854 462 3857 668
rect 3866 598 3873 601
rect 3870 552 3873 598
rect 3902 432 3905 448
rect 3806 372 3809 378
rect 3814 352 3817 368
rect 3762 238 3766 241
rect 3746 78 3753 81
rect 3758 52 3761 208
rect 3774 202 3777 258
rect 3782 222 3785 258
rect 3782 162 3785 208
rect 3766 112 3769 128
rect 3778 108 3785 111
rect 3782 102 3785 108
rect 3766 81 3769 88
rect 3766 78 3774 81
rect 3790 81 3793 298
rect 3814 252 3817 268
rect 3806 112 3809 168
rect 3790 78 3798 81
rect 2974 48 2982 51
rect 3014 48 3022 51
rect 3014 42 3017 48
rect 3302 42 3305 48
rect 3790 42 3793 58
rect 3798 52 3801 58
rect 3814 52 3817 88
rect 3822 72 3825 268
rect 3830 142 3833 148
rect 3838 82 3841 278
rect 3878 171 3881 198
rect 3870 168 3881 171
rect 3854 112 3857 138
rect 3870 112 3873 168
rect 3886 132 3889 188
rect 3886 101 3889 108
rect 3870 98 3889 101
rect 3850 88 3854 91
rect 3870 82 3873 98
rect 3882 78 3886 81
rect 3846 52 3849 78
rect 3894 72 3897 268
rect 3902 132 3905 248
rect 3910 131 3913 458
rect 3918 342 3921 728
rect 3942 522 3945 538
rect 3958 422 3961 978
rect 3966 852 3969 908
rect 3974 791 3977 1178
rect 3982 1082 3985 1088
rect 3982 952 3985 958
rect 3990 952 3993 1468
rect 3998 1442 4001 1528
rect 4006 1362 4009 1598
rect 4014 1462 4017 1468
rect 4022 1362 4025 1568
rect 4054 1532 4057 1898
rect 4070 1882 4073 1908
rect 4080 1903 4082 1907
rect 4086 1903 4089 1907
rect 4094 1903 4096 1907
rect 4030 1422 4033 1458
rect 4014 1282 4017 1358
rect 4022 1222 4025 1348
rect 4030 1332 4033 1338
rect 4030 1282 4033 1298
rect 3974 788 3982 791
rect 3966 452 3969 498
rect 3974 472 3977 598
rect 3954 378 3958 381
rect 3918 222 3921 268
rect 3918 142 3921 178
rect 3910 128 3921 131
rect 3910 112 3913 118
rect 3866 68 3870 71
rect 3854 42 3857 58
rect 3322 28 3326 31
rect 3886 22 3889 28
rect 3902 22 3905 58
rect 3910 22 3913 78
rect 3918 62 3921 128
rect 3926 81 3929 368
rect 3966 281 3969 398
rect 3974 362 3977 468
rect 3998 352 4001 1178
rect 4010 1158 4014 1161
rect 4022 1042 4025 1178
rect 4030 1142 4033 1188
rect 4030 1112 4033 1138
rect 4038 1082 4041 1518
rect 4062 1432 4065 1548
rect 4054 1251 4057 1388
rect 4054 1248 4062 1251
rect 4038 1052 4041 1068
rect 4046 1062 4049 1228
rect 4006 1022 4009 1028
rect 4006 842 4009 848
rect 4014 761 4017 1028
rect 4010 758 4017 761
rect 4010 748 4014 751
rect 4022 742 4025 1018
rect 4030 922 4033 938
rect 4038 922 4041 1038
rect 4034 838 4041 841
rect 4038 822 4041 838
rect 4030 742 4033 748
rect 3994 338 3998 341
rect 3974 332 3977 338
rect 3990 322 3993 328
rect 3966 278 3974 281
rect 3938 258 3945 261
rect 3942 242 3945 258
rect 3942 222 3945 238
rect 3958 182 3961 218
rect 3982 212 3985 258
rect 3946 158 3953 161
rect 3950 152 3953 158
rect 3934 122 3937 138
rect 3946 128 3953 131
rect 3950 112 3953 128
rect 3958 101 3961 148
rect 3950 98 3961 101
rect 3926 78 3934 81
rect 3950 72 3953 98
rect 3934 52 3937 68
rect 3966 62 3969 208
rect 3974 132 3977 138
rect 4006 131 4009 618
rect 4014 502 4017 578
rect 4014 332 4017 348
rect 3998 128 4009 131
rect 3998 92 4001 128
rect 4006 102 4009 118
rect 3974 72 3977 78
rect 3946 28 3950 31
rect 3958 12 3961 28
rect 3966 12 3969 48
rect 4014 42 4017 318
rect 4022 62 4025 508
rect 4030 472 4033 588
rect 4038 542 4041 788
rect 4038 442 4041 458
rect 4038 302 4041 438
rect 4038 162 4041 208
rect 4030 72 4033 108
rect 4038 102 4041 138
rect 4046 72 4049 1048
rect 4054 932 4057 1248
rect 4062 962 4065 1208
rect 4070 1142 4073 1778
rect 4080 1703 4082 1707
rect 4086 1703 4089 1707
rect 4094 1703 4096 1707
rect 4078 1582 4081 1588
rect 4080 1503 4082 1507
rect 4086 1503 4089 1507
rect 4094 1503 4096 1507
rect 4080 1303 4082 1307
rect 4086 1303 4089 1307
rect 4094 1303 4096 1307
rect 4094 1272 4097 1278
rect 4102 1182 4105 1538
rect 4070 1112 4073 1128
rect 4080 1103 4082 1107
rect 4086 1103 4089 1107
rect 4094 1103 4096 1107
rect 4094 1042 4097 1048
rect 4110 972 4113 1678
rect 4118 1522 4121 2978
rect 4142 2472 4145 2518
rect 4146 2358 4150 2361
rect 4158 2332 4161 2338
rect 4126 2152 4129 2288
rect 4134 2192 4137 2258
rect 4130 1878 4137 1881
rect 4134 1872 4137 1878
rect 4142 1742 4145 1948
rect 4166 1932 4169 1958
rect 4118 1052 4121 1478
rect 4134 1232 4137 1448
rect 4142 1312 4145 1608
rect 4154 1578 4158 1581
rect 4174 1572 4177 3388
rect 4214 3272 4217 3538
rect 4206 2652 4209 2708
rect 4186 2538 4190 2541
rect 4190 2512 4193 2538
rect 4182 2452 4185 2498
rect 4214 2392 4217 2418
rect 4210 2368 4217 2371
rect 4198 2262 4201 2268
rect 4190 1941 4193 2078
rect 4198 1952 4201 1978
rect 4190 1938 4201 1941
rect 4182 1702 4185 1748
rect 4182 1622 4185 1648
rect 4170 1548 4174 1551
rect 4166 1502 4169 1518
rect 4154 1458 4158 1461
rect 4134 1162 4137 1168
rect 4126 1112 4129 1138
rect 4090 948 4094 951
rect 4102 942 4105 948
rect 4110 942 4113 968
rect 4070 862 4073 918
rect 4080 903 4082 907
rect 4086 903 4089 907
rect 4094 903 4096 907
rect 4058 728 4062 731
rect 4054 482 4057 528
rect 4054 342 4057 348
rect 4054 232 4057 238
rect 4062 201 4065 718
rect 4070 632 4073 738
rect 4080 703 4082 707
rect 4086 703 4089 707
rect 4094 703 4096 707
rect 4070 592 4073 628
rect 4078 552 4081 578
rect 4080 503 4082 507
rect 4086 503 4089 507
rect 4094 503 4096 507
rect 4070 312 4073 338
rect 4080 303 4082 307
rect 4086 303 4089 307
rect 4094 303 4096 307
rect 4070 232 4073 298
rect 4078 222 4081 238
rect 4054 198 4065 201
rect 4054 132 4057 198
rect 4062 132 4065 168
rect 4086 152 4089 258
rect 4094 222 4097 248
rect 4070 112 4073 128
rect 4080 103 4082 107
rect 4086 103 4089 107
rect 4094 103 4096 107
rect 4102 92 4105 908
rect 4142 842 4145 1198
rect 4150 1092 4153 1458
rect 4158 1182 4161 1398
rect 4166 1192 4169 1448
rect 4174 1392 4177 1518
rect 4182 1372 4185 1538
rect 4190 1402 4193 1658
rect 4198 1512 4201 1938
rect 4206 1572 4209 2158
rect 4214 1502 4217 2368
rect 4186 1368 4193 1371
rect 4174 1262 4177 1268
rect 4158 1172 4161 1178
rect 4158 1122 4161 1128
rect 4182 1112 4185 1188
rect 4190 1092 4193 1368
rect 4210 1338 4214 1341
rect 4198 1152 4201 1218
rect 4206 1162 4209 1228
rect 4214 1112 4217 1318
rect 4214 1082 4217 1088
rect 4190 1002 4193 1008
rect 4158 852 4161 858
rect 4110 592 4113 748
rect 4118 652 4121 788
rect 4110 132 4113 518
rect 4118 112 4121 628
rect 4126 572 4129 788
rect 4134 732 4137 838
rect 4166 832 4169 998
rect 4174 952 4177 958
rect 4190 942 4193 998
rect 4198 952 4201 1068
rect 4134 642 4137 728
rect 4146 668 4150 671
rect 4126 541 4129 548
rect 4126 538 4134 541
rect 4126 112 4129 198
rect 4110 32 4113 98
rect 4134 82 4137 198
rect 4142 72 4145 488
rect 4150 352 4153 668
rect 4158 612 4161 748
rect 4158 542 4161 608
rect 4174 402 4177 928
rect 4182 822 4185 908
rect 4182 442 4185 658
rect 4190 542 4193 938
rect 4210 878 4214 881
rect 4150 272 4153 348
rect 4150 172 4153 178
rect 4150 142 4153 168
rect 4158 162 4161 168
rect 4158 152 4161 158
rect 4166 132 4169 148
rect 4174 132 4177 388
rect 4182 182 4185 398
rect 4198 262 4201 858
rect 4206 782 4209 798
rect 4206 752 4209 768
rect 4214 742 4217 828
rect 4222 622 4225 3588
rect 4262 3122 4265 3238
rect 4230 2592 4233 2738
rect 4230 2572 4233 2588
rect 4254 2302 4257 3028
rect 4262 2232 4265 2888
rect 4310 2572 4313 4308
rect 4322 4228 4329 4231
rect 4326 4072 4329 4228
rect 4334 4172 4337 4338
rect 4350 4332 4353 4338
rect 4350 4262 4353 4328
rect 4358 4322 4361 4328
rect 4358 4241 4361 4318
rect 4354 4238 4361 4241
rect 4358 4072 4361 4238
rect 4366 4052 4369 4388
rect 4374 4042 4377 4398
rect 4442 4358 4446 4361
rect 4490 4348 4494 4351
rect 4382 4252 4385 4258
rect 4322 3758 4329 3761
rect 4318 3642 4321 3748
rect 4326 3692 4329 3758
rect 4334 3642 4337 3818
rect 4350 3752 4353 4038
rect 4370 3938 4374 3941
rect 4398 3862 4401 4348
rect 4406 3872 4409 4338
rect 4414 3952 4417 4178
rect 4422 3882 4425 4328
rect 4430 4192 4433 4278
rect 4430 3972 4433 4188
rect 4438 3942 4441 4118
rect 4322 3638 4329 3641
rect 4318 3342 4321 3478
rect 4326 3212 4329 3638
rect 4318 2958 4326 2961
rect 4318 2942 4321 2958
rect 4306 2558 4310 2561
rect 4326 2542 4329 2578
rect 4334 2531 4337 3148
rect 4334 2528 4342 2531
rect 4326 2501 4329 2528
rect 4322 2498 4329 2501
rect 4334 2492 4337 2528
rect 4346 2368 4350 2371
rect 4274 2348 4278 2351
rect 4310 2322 4313 2328
rect 4258 2118 4265 2121
rect 4262 2082 4265 2118
rect 4250 2068 4254 2071
rect 4270 2062 4273 2068
rect 4230 1612 4233 1748
rect 4246 1701 4249 1988
rect 4258 1918 4262 1921
rect 4254 1882 4257 1888
rect 4286 1852 4289 2178
rect 4302 2062 4305 2148
rect 4294 1921 4297 1948
rect 4294 1918 4302 1921
rect 4242 1698 4249 1701
rect 4238 1612 4241 1618
rect 4234 1598 4238 1601
rect 4234 1568 4238 1571
rect 4230 1542 4233 1548
rect 4230 1452 4233 1468
rect 4238 1462 4241 1468
rect 4230 1322 4233 1408
rect 4246 1392 4249 1638
rect 4254 1632 4257 1738
rect 4254 1562 4257 1628
rect 4262 1562 4265 1568
rect 4254 1402 4257 1538
rect 4278 1522 4281 1578
rect 4262 1458 4270 1461
rect 4262 1372 4265 1458
rect 4238 1352 4241 1358
rect 4238 1202 4241 1228
rect 4254 1162 4257 1258
rect 4270 1171 4273 1378
rect 4278 1182 4281 1298
rect 4270 1168 4281 1171
rect 4234 1128 4238 1131
rect 4238 1072 4241 1078
rect 4230 922 4233 948
rect 4206 292 4209 598
rect 4214 542 4217 618
rect 4230 611 4233 848
rect 4238 682 4241 898
rect 4246 672 4249 1138
rect 4222 608 4233 611
rect 4214 282 4217 328
rect 4222 312 4225 608
rect 4238 562 4241 668
rect 4230 352 4233 558
rect 4238 442 4241 468
rect 4246 372 4249 668
rect 4254 372 4257 1158
rect 4262 1042 4265 1148
rect 4270 952 4273 958
rect 4278 892 4281 1168
rect 4286 862 4289 1738
rect 4310 1722 4313 2308
rect 4326 2272 4329 2348
rect 4338 2328 4342 2331
rect 4326 2192 4329 2268
rect 4350 2122 4353 2248
rect 4318 1762 4321 2058
rect 4342 1902 4345 1928
rect 4350 1752 4353 2078
rect 4358 1692 4361 3768
rect 4374 3622 4377 3858
rect 4374 3051 4377 3138
rect 4370 3048 4377 3051
rect 4366 2362 4369 2418
rect 4382 2342 4385 3748
rect 4438 3732 4441 3838
rect 4374 2308 4382 2311
rect 4374 2262 4377 2308
rect 4374 1762 4377 1788
rect 4370 1678 4374 1681
rect 4306 1638 4310 1641
rect 4390 1592 4393 3288
rect 4406 3082 4409 3198
rect 4406 2122 4409 2368
rect 4398 2002 4401 2118
rect 4406 1972 4409 1978
rect 4398 1751 4401 1958
rect 4398 1748 4406 1751
rect 4402 1648 4406 1651
rect 4398 1571 4401 1578
rect 4394 1568 4401 1571
rect 4346 1548 4353 1551
rect 4402 1548 4406 1551
rect 4294 1538 4302 1541
rect 4294 1372 4297 1538
rect 4302 1392 4305 1528
rect 4310 1458 4318 1461
rect 4310 1452 4313 1458
rect 4298 1248 4302 1251
rect 4294 932 4297 1078
rect 4266 858 4270 861
rect 4294 852 4297 858
rect 4282 848 4286 851
rect 4302 792 4305 1008
rect 4310 922 4313 1448
rect 4318 1262 4321 1348
rect 4326 1212 4329 1418
rect 4322 1128 4329 1131
rect 4326 1022 4329 1128
rect 4334 1052 4337 1458
rect 4350 1442 4353 1548
rect 4342 1122 4345 1328
rect 4342 1082 4345 1088
rect 4318 862 4321 948
rect 4262 742 4265 748
rect 4270 522 4273 528
rect 4230 328 4238 331
rect 4246 331 4249 358
rect 4246 328 4254 331
rect 4218 258 4225 261
rect 4174 81 4177 128
rect 4182 92 4185 178
rect 4190 92 4193 168
rect 4214 152 4217 228
rect 4222 222 4225 258
rect 4230 172 4233 328
rect 4258 198 4262 201
rect 4242 158 4246 161
rect 4174 78 4185 81
rect 4126 68 4134 71
rect 4126 62 4129 68
rect 4174 62 4177 68
rect 4182 51 4185 78
rect 4182 48 4190 51
rect 4198 42 4201 148
rect 4206 142 4209 148
rect 4222 22 4225 148
rect 4262 82 4265 128
rect 4270 92 4273 368
rect 4278 332 4281 728
rect 4310 552 4313 568
rect 4294 462 4297 538
rect 4314 438 4321 441
rect 4278 92 4281 258
rect 4286 242 4289 348
rect 4294 242 4297 248
rect 4270 82 4273 88
rect 4230 52 4233 78
rect 4254 72 4257 78
rect 4270 62 4273 68
rect 4302 42 4305 418
rect 4318 292 4321 438
rect 4334 402 4337 848
rect 4350 822 4353 1388
rect 4358 1262 4361 1308
rect 4358 972 4361 1088
rect 4374 981 4377 1228
rect 4382 1022 4385 1468
rect 4390 1012 4393 1488
rect 4406 1362 4409 1448
rect 4414 1202 4417 3718
rect 4430 2572 4433 3568
rect 4446 3431 4449 4348
rect 4462 4332 4465 4338
rect 4458 4298 4462 4301
rect 4454 4112 4457 4278
rect 4470 4258 4478 4261
rect 4470 4112 4473 4258
rect 4454 3472 4457 4098
rect 4470 3942 4473 4078
rect 4478 4051 4481 4238
rect 4486 4062 4489 4258
rect 4478 4048 4489 4051
rect 4478 3942 4481 3958
rect 4446 3428 4457 3431
rect 4438 3112 4441 3138
rect 4446 2862 4449 3158
rect 4430 2062 4433 2148
rect 4438 1801 4441 2818
rect 4434 1798 4441 1801
rect 4422 1172 4425 1728
rect 4438 1162 4441 1178
rect 4402 1048 4406 1051
rect 4386 988 4390 991
rect 4374 978 4385 981
rect 4362 958 4366 961
rect 4342 472 4345 718
rect 4350 582 4353 628
rect 4358 462 4361 728
rect 4314 258 4321 261
rect 4318 192 4321 258
rect 4318 182 4321 188
rect 4310 112 4313 178
rect 4334 102 4337 128
rect 4342 122 4345 148
rect 4354 138 4358 141
rect 4350 112 4353 128
rect 4342 62 4345 78
rect 4366 32 4369 828
rect 4374 732 4377 738
rect 4374 152 4377 718
rect 4382 32 4385 978
rect 4390 252 4393 558
rect 4398 72 4401 918
rect 4406 862 4409 988
rect 4414 972 4417 1098
rect 4406 282 4409 738
rect 4414 52 4417 928
rect 4422 862 4425 1108
rect 4422 492 4425 698
rect 4422 472 4425 478
rect 4430 82 4433 1068
rect 4438 1042 4441 1148
rect 4438 1002 4441 1028
rect 4438 872 4441 878
rect 4438 362 4441 748
rect 4446 312 4449 2858
rect 4454 2122 4457 3428
rect 4454 1922 4457 1928
rect 4454 1672 4457 1918
rect 4462 1292 4465 3668
rect 4454 1072 4457 1168
rect 4462 1072 4465 1238
rect 4454 1052 4457 1058
rect 4454 842 4457 948
rect 4454 502 4457 548
rect 4462 462 4465 928
rect 4458 448 4462 451
rect 4438 92 4441 128
rect 4470 82 4473 3728
rect 4478 3152 4481 3638
rect 4478 2392 4481 2798
rect 4486 2292 4489 4048
rect 4510 3832 4513 4338
rect 4494 3382 4497 3538
rect 4502 3438 4510 3441
rect 4502 3312 4505 3438
rect 4510 2712 4513 3148
rect 4510 2352 4513 2368
rect 4478 1782 4481 2058
rect 4478 1412 4481 1458
rect 4478 1132 4481 1408
rect 4486 1402 4489 2078
rect 4494 1432 4497 2238
rect 4502 2132 4505 2138
rect 4510 1732 4513 2338
rect 4518 2302 4521 4308
rect 4526 3862 4529 4348
rect 4550 4302 4553 4308
rect 4534 4092 4537 4278
rect 4534 3912 4537 4078
rect 4550 3951 4553 4208
rect 4558 4172 4561 4328
rect 4566 4252 4569 4258
rect 4558 4032 4561 4168
rect 4550 3948 4558 3951
rect 4550 3852 4553 3888
rect 4526 3262 4529 3648
rect 4526 2382 4529 3258
rect 4558 3142 4561 3858
rect 4566 3732 4569 4218
rect 4562 3138 4566 3141
rect 4534 3042 4537 3068
rect 4550 2862 4553 2958
rect 4566 2842 4569 2968
rect 4546 2548 4550 2551
rect 4530 2368 4534 2371
rect 4522 2258 4526 2261
rect 4518 1812 4521 1908
rect 4522 1648 4526 1651
rect 4486 1162 4489 1368
rect 4498 1348 4502 1351
rect 4510 1252 4513 1548
rect 4526 1372 4529 1638
rect 4478 92 4481 1078
rect 4486 962 4489 1078
rect 4534 931 4537 2088
rect 4542 952 4545 2378
rect 4574 2352 4577 4288
rect 4582 3722 4585 4348
rect 4590 3252 4593 4148
rect 4598 3962 4601 4118
rect 4598 3752 4601 3808
rect 4598 2782 4601 2868
rect 4590 2341 4593 2478
rect 4582 2338 4593 2341
rect 4566 2322 4569 2328
rect 4558 2061 4561 2068
rect 4554 2058 4561 2061
rect 4566 1922 4569 2318
rect 4574 2042 4577 2068
rect 4570 1528 4574 1531
rect 4550 1262 4553 1488
rect 4558 1472 4561 1498
rect 4558 1442 4561 1458
rect 4558 1042 4561 1438
rect 4574 1402 4577 1468
rect 4566 1022 4569 1348
rect 4526 928 4537 931
rect 4526 912 4529 928
rect 4486 842 4489 878
rect 4514 858 4521 861
rect 4490 838 4497 841
rect 4486 292 4489 598
rect 4494 332 4497 838
rect 4518 792 4521 858
rect 4502 372 4505 708
rect 4510 452 4513 548
rect 4518 432 4521 618
rect 4486 202 4489 278
rect 4506 148 4513 151
rect 4510 72 4513 148
rect 4526 72 4529 898
rect 4534 142 4537 918
rect 4542 772 4545 928
rect 4550 442 4553 948
rect 4558 932 4561 938
rect 4562 678 4569 681
rect 4566 662 4569 678
rect 4574 562 4577 1378
rect 4570 538 4574 541
rect 4574 472 4577 478
rect 4582 352 4585 2338
rect 4594 1678 4598 1681
rect 4590 1272 4593 1278
rect 4598 1002 4601 1158
rect 4590 662 4593 848
rect 4542 332 4545 338
rect 4542 152 4545 158
rect 4598 122 4601 998
rect 4078 12 4081 18
rect 4534 12 4537 78
rect 1030 8 1038 11
rect 496 3 498 7
rect 502 3 505 7
rect 510 3 512 7
rect 1520 3 1522 7
rect 1526 3 1529 7
rect 1534 3 1536 7
rect 2544 3 2546 7
rect 2550 3 2553 7
rect 2558 3 2560 7
rect 3568 3 3570 7
rect 3574 3 3577 7
rect 3582 3 3584 7
<< m5contact >>
rect 498 4403 502 4407
rect 505 4403 506 4407
rect 506 4403 509 4407
rect 1522 4403 1526 4407
rect 1529 4403 1530 4407
rect 1530 4403 1533 4407
rect 2546 4403 2550 4407
rect 2553 4403 2554 4407
rect 2554 4403 2557 4407
rect 3570 4403 3574 4407
rect 3577 4403 3578 4407
rect 3578 4403 3581 4407
rect 4006 4398 4010 4402
rect 4254 4398 4258 4402
rect 1758 4338 1762 4342
rect 270 4148 274 4152
rect 526 4248 530 4252
rect 470 4238 474 4242
rect 498 4203 502 4207
rect 505 4203 506 4207
rect 506 4203 509 4207
rect 302 3268 306 3272
rect 326 3268 330 3272
rect 498 4003 502 4007
rect 505 4003 506 4007
rect 506 4003 509 4007
rect 286 2068 290 2072
rect 318 2068 322 2072
rect 446 2148 450 2152
rect 478 2078 482 2082
rect 390 1968 394 1972
rect 318 1938 322 1942
rect 302 1548 306 1552
rect 498 3803 502 3807
rect 505 3803 506 3807
rect 506 3803 509 3807
rect 1002 4303 1006 4307
rect 1009 4303 1010 4307
rect 1010 4303 1013 4307
rect 862 4268 866 4272
rect 806 4248 810 4252
rect 678 4228 682 4232
rect 638 4148 642 4152
rect 498 3603 502 3607
rect 505 3603 506 3607
rect 506 3603 509 3607
rect 498 3403 502 3407
rect 505 3403 506 3407
rect 506 3403 509 3407
rect 494 3268 498 3272
rect 498 3203 502 3207
rect 505 3203 506 3207
rect 506 3203 509 3207
rect 1102 4268 1106 4272
rect 1566 4268 1570 4272
rect 1126 4258 1130 4262
rect 1198 4258 1202 4262
rect 1246 4258 1250 4262
rect 942 4238 946 4242
rect 498 3003 502 3007
rect 505 3003 506 3007
rect 506 3003 509 3007
rect 498 2803 502 2807
rect 505 2803 506 2807
rect 506 2803 509 2807
rect 614 2648 618 2652
rect 498 2603 502 2607
rect 505 2603 506 2607
rect 506 2603 509 2607
rect 782 3738 786 3742
rect 646 2748 650 2752
rect 654 2678 658 2682
rect 710 2648 714 2652
rect 750 2658 754 2662
rect 498 2403 502 2407
rect 505 2403 506 2407
rect 506 2403 509 2407
rect 498 2203 502 2207
rect 505 2203 506 2207
rect 506 2203 509 2207
rect 646 2128 650 2132
rect 1046 4148 1050 4152
rect 1310 4158 1314 4162
rect 1254 4128 1258 4132
rect 934 3948 938 3952
rect 790 2678 794 2682
rect 798 2148 802 2152
rect 498 2003 502 2007
rect 505 2003 506 2007
rect 506 2003 509 2007
rect 398 1168 402 1172
rect 498 1803 502 1807
rect 505 1803 506 1807
rect 506 1803 509 1807
rect 550 1688 554 1692
rect 498 1603 502 1607
rect 505 1603 506 1607
rect 506 1603 509 1607
rect 510 1548 514 1552
rect 498 1403 502 1407
rect 505 1403 506 1407
rect 506 1403 509 1407
rect 598 1678 602 1682
rect 822 2658 826 2662
rect 926 3278 930 3282
rect 1002 4103 1006 4107
rect 1009 4103 1010 4107
rect 1010 4103 1013 4107
rect 1002 3903 1006 3907
rect 1009 3903 1010 3907
rect 1010 3903 1013 3907
rect 1002 3703 1006 3707
rect 1009 3703 1010 3707
rect 1010 3703 1013 3707
rect 990 3658 994 3662
rect 1002 3503 1006 3507
rect 1009 3503 1010 3507
rect 1010 3503 1013 3507
rect 1102 3828 1106 3832
rect 1002 3303 1006 3307
rect 1009 3303 1010 3307
rect 1010 3303 1013 3307
rect 966 3268 970 3272
rect 1002 3103 1006 3107
rect 1009 3103 1010 3107
rect 1010 3103 1013 3107
rect 910 3078 914 3082
rect 854 2138 858 2142
rect 886 2748 890 2752
rect 894 2688 898 2692
rect 902 2328 906 2332
rect 870 1988 874 1992
rect 894 2028 898 2032
rect 878 1768 882 1772
rect 862 1758 866 1762
rect 606 1578 610 1582
rect 206 468 210 472
rect 246 648 250 652
rect 182 268 186 272
rect 238 258 242 262
rect 310 658 314 662
rect 286 458 290 462
rect 498 1203 502 1207
rect 505 1203 506 1207
rect 506 1203 509 1207
rect 462 1158 466 1162
rect 486 1158 490 1162
rect 498 1003 502 1007
rect 505 1003 506 1007
rect 506 1003 509 1007
rect 498 803 502 807
rect 505 803 506 807
rect 506 803 509 807
rect 430 648 434 652
rect 498 603 502 607
rect 505 603 506 607
rect 506 603 509 607
rect 558 658 562 662
rect 382 468 386 472
rect 498 403 502 407
rect 505 403 506 407
rect 506 403 509 407
rect 366 248 370 252
rect 498 203 502 207
rect 505 203 506 207
rect 506 203 509 207
rect 262 148 266 152
rect 782 1578 786 1582
rect 1002 2903 1006 2907
rect 1009 2903 1010 2907
rect 1010 2903 1013 2907
rect 1038 2858 1042 2862
rect 1002 2703 1006 2707
rect 1009 2703 1010 2707
rect 1010 2703 1013 2707
rect 1022 2618 1026 2622
rect 918 2478 922 2482
rect 1002 2503 1006 2507
rect 1009 2503 1010 2507
rect 1010 2503 1013 2507
rect 1038 2488 1042 2492
rect 1006 2478 1010 2482
rect 934 2338 938 2342
rect 942 2328 946 2332
rect 918 1968 922 1972
rect 918 1938 922 1942
rect 966 1878 970 1882
rect 974 1788 978 1792
rect 614 268 618 272
rect 606 248 610 252
rect 686 118 690 122
rect 942 868 946 872
rect 1002 2303 1006 2307
rect 1009 2303 1010 2307
rect 1010 2303 1013 2307
rect 990 2118 994 2122
rect 1002 2103 1006 2107
rect 1009 2103 1010 2107
rect 1010 2103 1013 2107
rect 1006 2068 1010 2072
rect 1002 1903 1006 1907
rect 1009 1903 1010 1907
rect 1010 1903 1013 1907
rect 1002 1703 1006 1707
rect 1009 1703 1010 1707
rect 1010 1703 1013 1707
rect 1054 2688 1058 2692
rect 1230 3388 1234 3392
rect 1102 2688 1106 2692
rect 1078 2478 1082 2482
rect 1166 3278 1170 3282
rect 1102 2068 1106 2072
rect 1070 2058 1074 2062
rect 1134 1868 1138 1872
rect 1110 1728 1114 1732
rect 1002 1503 1006 1507
rect 1009 1503 1010 1507
rect 1010 1503 1013 1507
rect 1002 1303 1006 1307
rect 1009 1303 1010 1307
rect 1010 1303 1013 1307
rect 1002 1103 1006 1107
rect 1009 1103 1010 1107
rect 1010 1103 1013 1107
rect 1078 958 1082 962
rect 1070 948 1074 952
rect 1014 938 1018 942
rect 1002 903 1006 907
rect 1009 903 1010 907
rect 1010 903 1013 907
rect 1118 868 1122 872
rect 1002 703 1006 707
rect 1009 703 1010 707
rect 1010 703 1013 707
rect 1002 503 1006 507
rect 1009 503 1010 507
rect 1010 503 1013 507
rect 934 158 938 162
rect 1002 303 1006 307
rect 1009 303 1010 307
rect 1010 303 1013 307
rect 1002 103 1006 107
rect 1009 103 1010 107
rect 1010 103 1013 107
rect 918 58 922 62
rect 1158 1748 1162 1752
rect 1222 2918 1226 2922
rect 1254 2918 1258 2922
rect 1190 2468 1194 2472
rect 1206 2468 1210 2472
rect 1222 1728 1226 1732
rect 1222 1688 1226 1692
rect 1230 1678 1234 1682
rect 1206 1558 1210 1562
rect 1182 1268 1186 1272
rect 1174 1168 1178 1172
rect 1190 848 1194 852
rect 1214 948 1218 952
rect 1198 458 1202 462
rect 1350 3838 1354 3842
rect 1318 3388 1322 3392
rect 1302 3088 1306 3092
rect 1270 2618 1274 2622
rect 1270 2338 1274 2342
rect 1278 1948 1282 1952
rect 1334 2658 1338 2662
rect 1334 2128 1338 2132
rect 1470 4238 1474 4242
rect 1438 4158 1442 4162
rect 1398 4088 1402 4092
rect 1522 4203 1526 4207
rect 1529 4203 1530 4207
rect 1530 4203 1533 4207
rect 1694 4188 1698 4192
rect 1522 4003 1526 4007
rect 1529 4003 1530 4007
rect 1530 4003 1533 4007
rect 1526 3958 1530 3962
rect 1522 3803 1526 3807
rect 1529 3803 1530 3807
rect 1530 3803 1533 3807
rect 1522 3603 1526 3607
rect 1529 3603 1530 3607
rect 1530 3603 1533 3607
rect 1502 3548 1506 3552
rect 1518 3538 1522 3542
rect 1522 3403 1526 3407
rect 1529 3403 1530 3407
rect 1530 3403 1533 3407
rect 1486 3238 1490 3242
rect 1382 2618 1386 2622
rect 1366 2438 1370 2442
rect 1310 1678 1314 1682
rect 1522 3203 1526 3207
rect 1529 3203 1530 3207
rect 1530 3203 1533 3207
rect 1522 3003 1526 3007
rect 1529 3003 1530 3007
rect 1530 3003 1533 3007
rect 1542 2948 1546 2952
rect 1522 2803 1526 2807
rect 1529 2803 1530 2807
rect 1530 2803 1533 2807
rect 1422 2748 1426 2752
rect 1470 2658 1474 2662
rect 1454 2518 1458 2522
rect 1422 2468 1426 2472
rect 1414 2368 1418 2372
rect 1382 1748 1386 1752
rect 1406 848 1410 852
rect 1190 158 1194 162
rect 1454 1558 1458 1562
rect 1462 1418 1466 1422
rect 1454 958 1458 962
rect 1522 2603 1526 2607
rect 1529 2603 1530 2607
rect 1530 2603 1533 2607
rect 1574 3088 1578 3092
rect 1574 2858 1578 2862
rect 1542 2428 1546 2432
rect 1522 2403 1526 2407
rect 1529 2403 1530 2407
rect 1530 2403 1533 2407
rect 1522 2203 1526 2207
rect 1529 2203 1530 2207
rect 1530 2203 1533 2207
rect 1566 2408 1570 2412
rect 1550 2358 1554 2362
rect 1542 2138 1546 2142
rect 1510 2118 1514 2122
rect 1502 1828 1506 1832
rect 1522 2003 1526 2007
rect 1529 2003 1530 2007
rect 1530 2003 1533 2007
rect 1522 1803 1526 1807
rect 1529 1803 1530 1807
rect 1530 1803 1533 1807
rect 1542 1758 1546 1762
rect 1522 1603 1526 1607
rect 1529 1603 1530 1607
rect 1530 1603 1533 1607
rect 1522 1403 1526 1407
rect 1529 1403 1530 1407
rect 1530 1403 1533 1407
rect 1542 1268 1546 1272
rect 1522 1203 1526 1207
rect 1529 1203 1530 1207
rect 1530 1203 1533 1207
rect 1522 1003 1526 1007
rect 1529 1003 1530 1007
rect 1530 1003 1533 1007
rect 1486 938 1490 942
rect 1522 803 1526 807
rect 1529 803 1530 807
rect 1530 803 1533 807
rect 1566 1888 1570 1892
rect 1566 778 1570 782
rect 1522 603 1526 607
rect 1529 603 1530 607
rect 1530 603 1533 607
rect 1522 403 1526 407
rect 1529 403 1530 407
rect 1530 403 1533 407
rect 1614 3138 1618 3142
rect 1590 2268 1594 2272
rect 1598 2238 1602 2242
rect 1670 3088 1674 3092
rect 1670 2748 1674 2752
rect 1638 2438 1642 2442
rect 1590 1328 1594 1332
rect 1654 1478 1658 1482
rect 1646 1418 1650 1422
rect 1654 1258 1658 1262
rect 1654 1248 1658 1252
rect 1622 878 1626 882
rect 1630 618 1634 622
rect 1630 528 1634 532
rect 1606 418 1610 422
rect 1822 4268 1826 4272
rect 1990 4238 1994 4242
rect 1934 4228 1938 4232
rect 1958 4228 1962 4232
rect 1798 4158 1802 4162
rect 1910 4148 1914 4152
rect 1766 4138 1770 4142
rect 1838 4078 1842 4082
rect 1814 3958 1818 3962
rect 1774 3348 1778 3352
rect 1782 3248 1786 3252
rect 1814 3558 1818 3562
rect 1766 2668 1770 2672
rect 1846 3058 1850 3062
rect 1806 2468 1810 2472
rect 1694 2188 1698 2192
rect 1774 2168 1778 2172
rect 1734 2128 1738 2132
rect 1774 2058 1778 2062
rect 1694 2008 1698 2012
rect 1678 1998 1682 2002
rect 1686 1858 1690 1862
rect 1766 1978 1770 1982
rect 1742 1878 1746 1882
rect 1774 1968 1778 1972
rect 1782 1938 1786 1942
rect 1878 3088 1882 3092
rect 1846 1998 1850 2002
rect 1838 1948 1842 1952
rect 1822 1928 1826 1932
rect 1758 1858 1762 1862
rect 1790 1858 1794 1862
rect 1742 1768 1746 1772
rect 1758 1648 1762 1652
rect 1710 1478 1714 1482
rect 1678 1008 1682 1012
rect 1726 1258 1730 1262
rect 1734 918 1738 922
rect 1718 788 1722 792
rect 1742 668 1746 672
rect 1766 1458 1770 1462
rect 1726 538 1730 542
rect 1846 1828 1850 1832
rect 1854 1768 1858 1772
rect 1838 1538 1842 1542
rect 1774 748 1778 752
rect 1686 428 1690 432
rect 1710 358 1714 362
rect 1742 358 1746 362
rect 1598 258 1602 262
rect 1918 3358 1922 3362
rect 1910 3288 1914 3292
rect 1974 4118 1978 4122
rect 2026 4303 2030 4307
rect 2033 4303 2034 4307
rect 2034 4303 2037 4307
rect 2086 4288 2090 4292
rect 2262 4288 2266 4292
rect 2006 4248 2010 4252
rect 2026 4103 2030 4107
rect 2033 4103 2034 4107
rect 2034 4103 2037 4107
rect 2174 4258 2178 4262
rect 2158 4248 2162 4252
rect 2270 4248 2274 4252
rect 2238 4178 2242 4182
rect 2026 3903 2030 3907
rect 2033 3903 2034 3907
rect 2034 3903 2037 3907
rect 2102 3878 2106 3882
rect 2094 3868 2098 3872
rect 2026 3703 2030 3707
rect 2033 3703 2034 3707
rect 2034 3703 2037 3707
rect 1974 3548 1978 3552
rect 2006 3538 2010 3542
rect 2006 3518 2010 3522
rect 1950 3468 1954 3472
rect 1918 2888 1922 2892
rect 1902 2778 1906 2782
rect 1902 2358 1906 2362
rect 1894 2028 1898 2032
rect 1910 1988 1914 1992
rect 1870 1378 1874 1382
rect 1886 1308 1890 1312
rect 1894 1228 1898 1232
rect 1942 1918 1946 1922
rect 1942 1648 1946 1652
rect 1998 2958 2002 2962
rect 1974 2038 1978 2042
rect 1974 1318 1978 1322
rect 1910 1248 1914 1252
rect 1886 1148 1890 1152
rect 1862 1008 1866 1012
rect 1846 738 1850 742
rect 1934 1058 1938 1062
rect 1886 968 1890 972
rect 1878 948 1882 952
rect 1878 768 1882 772
rect 1878 758 1882 762
rect 1870 628 1874 632
rect 1910 748 1914 752
rect 2026 3503 2030 3507
rect 2033 3503 2034 3507
rect 2034 3503 2037 3507
rect 2030 3468 2034 3472
rect 2026 3303 2030 3307
rect 2033 3303 2034 3307
rect 2034 3303 2037 3307
rect 2026 3103 2030 3107
rect 2033 3103 2034 3107
rect 2034 3103 2037 3107
rect 2046 3038 2050 3042
rect 2022 2948 2026 2952
rect 2014 2938 2018 2942
rect 2026 2903 2030 2907
rect 2033 2903 2034 2907
rect 2034 2903 2037 2907
rect 2046 2888 2050 2892
rect 2026 2703 2030 2707
rect 2033 2703 2034 2707
rect 2034 2703 2037 2707
rect 2026 2503 2030 2507
rect 2033 2503 2034 2507
rect 2034 2503 2037 2507
rect 2014 2318 2018 2322
rect 2006 2248 2010 2252
rect 2026 2303 2030 2307
rect 2033 2303 2034 2307
rect 2034 2303 2037 2307
rect 2014 2118 2018 2122
rect 2026 2103 2030 2107
rect 2033 2103 2034 2107
rect 2034 2103 2037 2107
rect 2062 3738 2066 3742
rect 2182 3958 2186 3962
rect 2126 3658 2130 3662
rect 2110 3348 2114 3352
rect 2102 3258 2106 3262
rect 2054 2028 2058 2032
rect 2054 1958 2058 1962
rect 2026 1903 2030 1907
rect 2033 1903 2034 1907
rect 2034 1903 2037 1907
rect 2026 1703 2030 1707
rect 2033 1703 2034 1707
rect 2034 1703 2037 1707
rect 2026 1503 2030 1507
rect 2033 1503 2034 1507
rect 2034 1503 2037 1507
rect 2026 1303 2030 1307
rect 2033 1303 2034 1307
rect 2034 1303 2037 1307
rect 1998 1128 2002 1132
rect 2054 1128 2058 1132
rect 1998 1088 2002 1092
rect 1958 848 1962 852
rect 1950 688 1954 692
rect 1838 358 1842 362
rect 1846 338 1850 342
rect 1830 278 1834 282
rect 1918 348 1922 352
rect 2026 1103 2030 1107
rect 2033 1103 2034 1107
rect 2034 1103 2037 1107
rect 2006 1018 2010 1022
rect 2038 978 2042 982
rect 2022 958 2026 962
rect 2026 903 2030 907
rect 2033 903 2034 907
rect 2034 903 2037 907
rect 2014 858 2018 862
rect 2026 703 2030 707
rect 2033 703 2034 707
rect 2034 703 2037 707
rect 2038 678 2042 682
rect 2014 568 2018 572
rect 1974 478 1978 482
rect 1990 478 1994 482
rect 2054 998 2058 1002
rect 2086 3138 2090 3142
rect 2078 2418 2082 2422
rect 2094 2768 2098 2772
rect 2158 3558 2162 3562
rect 2182 3278 2186 3282
rect 2166 3188 2170 3192
rect 2142 2938 2146 2942
rect 2134 2548 2138 2552
rect 2254 4148 2258 4152
rect 2246 3868 2250 3872
rect 2270 3688 2274 3692
rect 2214 3278 2218 3282
rect 2198 3178 2202 3182
rect 2222 3158 2226 3162
rect 2222 3068 2226 3072
rect 2190 2678 2194 2682
rect 2118 1828 2122 1832
rect 2110 1818 2114 1822
rect 2094 1308 2098 1312
rect 2158 2028 2162 2032
rect 2150 1938 2154 1942
rect 2190 1928 2194 1932
rect 2190 1878 2194 1882
rect 2174 1848 2178 1852
rect 2158 1838 2162 1842
rect 2110 1088 2114 1092
rect 2126 898 2130 902
rect 2054 578 2058 582
rect 2046 538 2050 542
rect 2026 503 2030 507
rect 2033 503 2034 507
rect 2034 503 2037 507
rect 2126 868 2130 872
rect 2126 848 2130 852
rect 2126 598 2130 602
rect 1982 318 1986 322
rect 1522 203 1526 207
rect 1529 203 1530 207
rect 1530 203 1533 207
rect 1870 178 1874 182
rect 1886 158 1890 162
rect 1686 148 1690 152
rect 1510 118 1514 122
rect 1990 118 1994 122
rect 2026 303 2030 307
rect 2033 303 2034 307
rect 2034 303 2037 307
rect 2014 288 2018 292
rect 2126 368 2130 372
rect 2142 1158 2146 1162
rect 2214 2148 2218 2152
rect 2206 1788 2210 1792
rect 2278 3568 2282 3572
rect 2262 3248 2266 3252
rect 2302 3358 2306 3362
rect 2294 3338 2298 3342
rect 2278 3308 2282 3312
rect 2278 3288 2282 3292
rect 2262 3078 2266 3082
rect 2230 2958 2234 2962
rect 2238 2948 2242 2952
rect 2286 2938 2290 2942
rect 2262 2648 2266 2652
rect 2206 1618 2210 1622
rect 2166 1478 2170 1482
rect 2190 1418 2194 1422
rect 2190 948 2194 952
rect 2142 678 2146 682
rect 2270 2448 2274 2452
rect 2246 2388 2250 2392
rect 2238 2278 2242 2282
rect 2238 2098 2242 2102
rect 2238 1918 2242 1922
rect 2398 4258 2402 4262
rect 2350 4138 2354 4142
rect 2358 4118 2362 4122
rect 2390 4058 2394 4062
rect 2334 3718 2338 3722
rect 2326 3658 2330 3662
rect 2326 3588 2330 3592
rect 2334 3438 2338 3442
rect 2350 3418 2354 3422
rect 2366 3678 2370 3682
rect 2358 3398 2362 3402
rect 2318 3108 2322 3112
rect 2318 3058 2322 3062
rect 2310 2878 2314 2882
rect 2350 3378 2354 3382
rect 2342 3368 2346 3372
rect 2358 3298 2362 3302
rect 2350 3218 2354 3222
rect 2342 3038 2346 3042
rect 2414 4228 2418 4232
rect 2478 4268 2482 4272
rect 2510 4248 2514 4252
rect 2430 4178 2434 4182
rect 2438 4078 2442 4082
rect 2470 4058 2474 4062
rect 2654 4248 2658 4252
rect 2546 4203 2550 4207
rect 2553 4203 2554 4207
rect 2554 4203 2557 4207
rect 2758 4188 2762 4192
rect 2662 4088 2666 4092
rect 2630 4078 2634 4082
rect 2630 4068 2634 4072
rect 2590 4058 2594 4062
rect 2502 4048 2506 4052
rect 2622 4048 2626 4052
rect 2406 3938 2410 3942
rect 2422 3518 2426 3522
rect 2414 3388 2418 3392
rect 2430 3388 2434 3392
rect 2382 3318 2386 3322
rect 2406 3318 2410 3322
rect 2390 3308 2394 3312
rect 2382 3168 2386 3172
rect 2390 2668 2394 2672
rect 2334 2488 2338 2492
rect 2302 2408 2306 2412
rect 2294 2378 2298 2382
rect 2254 2048 2258 2052
rect 2254 2008 2258 2012
rect 2246 1738 2250 1742
rect 2374 2368 2378 2372
rect 2366 2328 2370 2332
rect 2382 2258 2386 2262
rect 2310 2178 2314 2182
rect 2334 2078 2338 2082
rect 2302 2058 2306 2062
rect 2302 1988 2306 1992
rect 2318 1918 2322 1922
rect 2286 1728 2290 1732
rect 2278 1468 2282 1472
rect 2254 1328 2258 1332
rect 2246 1268 2250 1272
rect 2246 1248 2250 1252
rect 2230 908 2234 912
rect 2214 878 2218 882
rect 2174 858 2178 862
rect 2158 578 2162 582
rect 2190 668 2194 672
rect 2222 868 2226 872
rect 2230 858 2234 862
rect 2174 488 2178 492
rect 2158 318 2162 322
rect 2150 308 2154 312
rect 2158 258 2162 262
rect 2222 508 2226 512
rect 2222 468 2226 472
rect 2334 1888 2338 1892
rect 2334 1718 2338 1722
rect 2406 2888 2410 2892
rect 2546 4003 2550 4007
rect 2553 4003 2554 4007
rect 2554 4003 2557 4007
rect 2566 3948 2570 3952
rect 2486 3878 2490 3882
rect 2494 3858 2498 3862
rect 2566 3858 2570 3862
rect 2550 3848 2554 3852
rect 2546 3803 2550 3807
rect 2553 3803 2554 3807
rect 2554 3803 2557 3807
rect 2534 3758 2538 3762
rect 2470 3648 2474 3652
rect 2478 3568 2482 3572
rect 2462 3178 2466 3182
rect 2502 3588 2506 3592
rect 2510 3568 2514 3572
rect 2526 3398 2530 3402
rect 2518 3358 2522 3362
rect 2518 3328 2522 3332
rect 2558 3658 2562 3662
rect 2546 3603 2550 3607
rect 2553 3603 2554 3607
rect 2554 3603 2557 3607
rect 2546 3403 2550 3407
rect 2553 3403 2554 3407
rect 2554 3403 2557 3407
rect 2558 3318 2562 3322
rect 2534 3258 2538 3262
rect 2438 3098 2442 3102
rect 2422 2228 2426 2232
rect 2406 2078 2410 2082
rect 2414 2068 2418 2072
rect 2406 2048 2410 2052
rect 2358 2018 2362 2022
rect 2374 1958 2378 1962
rect 2366 1868 2370 1872
rect 2342 1678 2346 1682
rect 2334 1538 2338 1542
rect 2318 1248 2322 1252
rect 2318 968 2322 972
rect 2318 828 2322 832
rect 2262 748 2266 752
rect 2270 708 2274 712
rect 2270 668 2274 672
rect 2342 1308 2346 1312
rect 2358 1358 2362 1362
rect 2342 858 2346 862
rect 2342 838 2346 842
rect 2334 788 2338 792
rect 2326 578 2330 582
rect 2366 948 2370 952
rect 2546 3203 2550 3207
rect 2553 3203 2554 3207
rect 2554 3203 2557 3207
rect 2486 3078 2490 3082
rect 2518 2948 2522 2952
rect 2494 2938 2498 2942
rect 2502 2868 2506 2872
rect 2462 2538 2466 2542
rect 2438 2068 2442 2072
rect 2438 2058 2442 2062
rect 2462 1778 2466 1782
rect 2462 1468 2466 1472
rect 2462 1348 2466 1352
rect 2438 1328 2442 1332
rect 2430 1158 2434 1162
rect 2390 1148 2394 1152
rect 2406 1138 2410 1142
rect 2390 938 2394 942
rect 2414 938 2418 942
rect 2382 878 2386 882
rect 2382 848 2386 852
rect 2406 728 2410 732
rect 2366 558 2370 562
rect 2398 518 2402 522
rect 2546 3003 2550 3007
rect 2553 3003 2554 3007
rect 2554 3003 2557 3007
rect 2574 3268 2578 3272
rect 2622 3468 2626 3472
rect 2654 3518 2658 3522
rect 2646 3458 2650 3462
rect 2546 2803 2550 2807
rect 2553 2803 2554 2807
rect 2554 2803 2557 2807
rect 2534 2718 2538 2722
rect 2546 2603 2550 2607
rect 2553 2603 2554 2607
rect 2554 2603 2557 2607
rect 2510 2458 2514 2462
rect 2546 2403 2550 2407
rect 2553 2403 2554 2407
rect 2554 2403 2557 2407
rect 2590 2478 2594 2482
rect 2546 2203 2550 2207
rect 2553 2203 2554 2207
rect 2554 2203 2557 2207
rect 2590 2158 2594 2162
rect 2590 2078 2594 2082
rect 2526 2068 2530 2072
rect 2546 2003 2550 2007
rect 2553 2003 2554 2007
rect 2554 2003 2557 2007
rect 2494 1928 2498 1932
rect 2630 1868 2634 1872
rect 2546 1803 2550 1807
rect 2553 1803 2554 1807
rect 2554 1803 2557 1807
rect 2494 1728 2498 1732
rect 2478 1458 2482 1462
rect 2478 1438 2482 1442
rect 2478 1108 2482 1112
rect 2478 1098 2482 1102
rect 2494 1088 2498 1092
rect 2622 1748 2626 1752
rect 2526 1678 2530 1682
rect 2630 1668 2634 1672
rect 2546 1603 2550 1607
rect 2553 1603 2554 1607
rect 2554 1603 2557 1607
rect 2558 1548 2562 1552
rect 2534 1428 2538 1432
rect 2546 1403 2550 1407
rect 2553 1403 2554 1407
rect 2554 1403 2557 1407
rect 2462 868 2466 872
rect 2502 958 2506 962
rect 2486 878 2490 882
rect 2470 838 2474 842
rect 2494 868 2498 872
rect 2518 958 2522 962
rect 2510 858 2514 862
rect 2510 838 2514 842
rect 2510 788 2514 792
rect 2494 658 2498 662
rect 2542 1278 2546 1282
rect 2546 1203 2550 1207
rect 2553 1203 2554 1207
rect 2554 1203 2557 1207
rect 2546 1003 2550 1007
rect 2553 1003 2554 1007
rect 2554 1003 2557 1007
rect 2550 968 2554 972
rect 2550 948 2554 952
rect 2574 948 2578 952
rect 2546 803 2550 807
rect 2553 803 2554 807
rect 2554 803 2557 807
rect 2534 798 2538 802
rect 2534 688 2538 692
rect 2462 468 2466 472
rect 2446 378 2450 382
rect 2390 368 2394 372
rect 2294 308 2298 312
rect 2230 238 2234 242
rect 2150 148 2154 152
rect 2198 138 2202 142
rect 2026 103 2030 107
rect 2033 103 2034 107
rect 2034 103 2037 107
rect 2302 248 2306 252
rect 2546 603 2550 607
rect 2553 603 2554 607
rect 2554 603 2557 607
rect 2546 403 2550 407
rect 2553 403 2554 407
rect 2554 403 2557 407
rect 2606 1268 2610 1272
rect 2646 3168 2650 3172
rect 2686 4158 2690 4162
rect 2702 4058 2706 4062
rect 2694 3658 2698 3662
rect 2710 3718 2714 3722
rect 2710 3688 2714 3692
rect 2710 3518 2714 3522
rect 2702 3428 2706 3432
rect 2734 3448 2738 3452
rect 2726 3408 2730 3412
rect 2678 3398 2682 3402
rect 2670 3158 2674 3162
rect 2710 3298 2714 3302
rect 2742 3108 2746 3112
rect 3050 4303 3054 4307
rect 3057 4303 3058 4307
rect 3058 4303 3061 4307
rect 2838 4268 2842 4272
rect 2894 4128 2898 4132
rect 2830 4068 2834 4072
rect 2798 3488 2802 3492
rect 2798 3458 2802 3462
rect 2782 3418 2786 3422
rect 2686 2888 2690 2892
rect 2670 2648 2674 2652
rect 2678 2488 2682 2492
rect 2654 2408 2658 2412
rect 2662 2398 2666 2402
rect 2662 2268 2666 2272
rect 2678 2238 2682 2242
rect 2654 2158 2658 2162
rect 2670 2088 2674 2092
rect 2662 1868 2666 1872
rect 2654 1718 2658 1722
rect 2678 1948 2682 1952
rect 2678 1568 2682 1572
rect 2670 1538 2674 1542
rect 2646 1368 2650 1372
rect 2590 1018 2594 1022
rect 2638 1348 2642 1352
rect 2670 1328 2674 1332
rect 2662 1318 2666 1322
rect 2614 1118 2618 1122
rect 2638 1088 2642 1092
rect 2622 1058 2626 1062
rect 2614 1028 2618 1032
rect 2590 828 2594 832
rect 2598 818 2602 822
rect 2654 1218 2658 1222
rect 2654 1138 2658 1142
rect 2678 1078 2682 1082
rect 2622 978 2626 982
rect 2646 958 2650 962
rect 2590 758 2594 762
rect 2614 718 2618 722
rect 2590 558 2594 562
rect 2590 458 2594 462
rect 2478 338 2482 342
rect 2414 228 2418 232
rect 2350 168 2354 172
rect 2382 148 2386 152
rect 2366 128 2370 132
rect 2374 118 2378 122
rect 2358 88 2362 92
rect 2542 258 2546 262
rect 2502 248 2506 252
rect 2518 238 2522 242
rect 2546 203 2550 207
rect 2553 203 2554 207
rect 2554 203 2557 207
rect 2678 928 2682 932
rect 2662 698 2666 702
rect 2630 448 2634 452
rect 2630 348 2634 352
rect 2678 348 2682 352
rect 2678 328 2682 332
rect 2726 2338 2730 2342
rect 2758 2858 2762 2862
rect 2750 2558 2754 2562
rect 2814 3868 2818 3872
rect 2814 3438 2818 3442
rect 2838 3658 2842 3662
rect 3230 4338 3234 4342
rect 2878 3868 2882 3872
rect 2886 3678 2890 3682
rect 2862 3658 2866 3662
rect 2886 3478 2890 3482
rect 2854 3388 2858 3392
rect 3050 4103 3054 4107
rect 3057 4103 3058 4107
rect 3058 4103 3061 4107
rect 2918 3378 2922 3382
rect 2878 3368 2882 3372
rect 2910 3338 2914 3342
rect 2870 3218 2874 3222
rect 2878 3158 2882 3162
rect 2774 2628 2778 2632
rect 2814 2528 2818 2532
rect 2758 2358 2762 2362
rect 2782 2278 2786 2282
rect 2750 2268 2754 2272
rect 2702 2128 2706 2132
rect 2726 2098 2730 2102
rect 2702 1938 2706 1942
rect 2878 3128 2882 3132
rect 2846 2918 2850 2922
rect 2846 2658 2850 2662
rect 2830 2568 2834 2572
rect 2838 2518 2842 2522
rect 2830 2368 2834 2372
rect 2822 2048 2826 2052
rect 2750 1888 2754 1892
rect 2702 1868 2706 1872
rect 2710 1628 2714 1632
rect 2702 1518 2706 1522
rect 2702 1458 2706 1462
rect 2726 1388 2730 1392
rect 2718 1268 2722 1272
rect 2702 1048 2706 1052
rect 2694 908 2698 912
rect 2694 838 2698 842
rect 2742 1528 2746 1532
rect 2750 1478 2754 1482
rect 2734 1298 2738 1302
rect 2726 1128 2730 1132
rect 2718 1118 2722 1122
rect 2718 1078 2722 1082
rect 2726 938 2730 942
rect 2694 688 2698 692
rect 2726 878 2730 882
rect 2726 848 2730 852
rect 2726 838 2730 842
rect 2750 1278 2754 1282
rect 2742 1138 2746 1142
rect 2750 1048 2754 1052
rect 2750 928 2754 932
rect 2742 868 2746 872
rect 2718 648 2722 652
rect 2702 638 2706 642
rect 2718 458 2722 462
rect 2702 448 2706 452
rect 2702 378 2706 382
rect 2710 378 2714 382
rect 2686 278 2690 282
rect 2734 558 2738 562
rect 2766 1058 2770 1062
rect 2766 928 2770 932
rect 2782 1158 2786 1162
rect 2798 1238 2802 1242
rect 2790 968 2794 972
rect 2846 1688 2850 1692
rect 2870 2868 2874 2872
rect 2870 2678 2874 2682
rect 2870 2478 2874 2482
rect 2862 2458 2866 2462
rect 2910 2748 2914 2752
rect 2894 2358 2898 2362
rect 2886 2348 2890 2352
rect 2902 2288 2906 2292
rect 2902 2258 2906 2262
rect 2894 2228 2898 2232
rect 2942 3668 2946 3672
rect 2950 3648 2954 3652
rect 2958 3468 2962 3472
rect 2990 3468 2994 3472
rect 2934 3458 2938 3462
rect 2934 3378 2938 3382
rect 3022 3458 3026 3462
rect 3006 3408 3010 3412
rect 2974 3358 2978 3362
rect 2998 3348 3002 3352
rect 2966 3338 2970 3342
rect 2958 2518 2962 2522
rect 2926 2388 2930 2392
rect 2934 2278 2938 2282
rect 2934 2258 2938 2262
rect 2950 2148 2954 2152
rect 2934 1928 2938 1932
rect 2934 1828 2938 1832
rect 2926 1718 2930 1722
rect 3050 3903 3054 3907
rect 3057 3903 3058 3907
rect 3058 3903 3061 3907
rect 3070 3848 3074 3852
rect 3050 3703 3054 3707
rect 3057 3703 3058 3707
rect 3058 3703 3061 3707
rect 3110 3668 3114 3672
rect 3050 3503 3054 3507
rect 3057 3503 3058 3507
rect 3058 3503 3061 3507
rect 3118 3488 3122 3492
rect 3086 3468 3090 3472
rect 3094 3458 3098 3462
rect 3094 3428 3098 3432
rect 3050 3303 3054 3307
rect 3057 3303 3058 3307
rect 3058 3303 3061 3307
rect 3050 3103 3054 3107
rect 3057 3103 3058 3107
rect 3058 3103 3061 3107
rect 3050 2903 3054 2907
rect 3057 2903 3058 2907
rect 3058 2903 3061 2907
rect 2990 2468 2994 2472
rect 2998 2418 3002 2422
rect 2982 2398 2986 2402
rect 2974 2388 2978 2392
rect 2982 2328 2986 2332
rect 2974 2148 2978 2152
rect 2998 1858 3002 1862
rect 2966 1758 2970 1762
rect 2998 1748 3002 1752
rect 3110 3278 3114 3282
rect 3086 2718 3090 2722
rect 3050 2703 3054 2707
rect 3057 2703 3058 2707
rect 3058 2703 3061 2707
rect 2974 1728 2978 1732
rect 3006 1728 3010 1732
rect 2918 1678 2922 1682
rect 2926 1668 2930 1672
rect 2870 1608 2874 1612
rect 2838 1568 2842 1572
rect 2878 1548 2882 1552
rect 2862 1538 2866 1542
rect 2902 1538 2906 1542
rect 2862 1498 2866 1502
rect 2838 1478 2842 1482
rect 2870 1478 2874 1482
rect 2846 1318 2850 1322
rect 2862 1278 2866 1282
rect 2838 1158 2842 1162
rect 2822 1088 2826 1092
rect 2830 1068 2834 1072
rect 2782 958 2786 962
rect 2806 958 2810 962
rect 2798 918 2802 922
rect 2798 748 2802 752
rect 2822 698 2826 702
rect 2806 658 2810 662
rect 2758 468 2762 472
rect 2766 288 2770 292
rect 2758 228 2762 232
rect 2422 138 2426 142
rect 2510 138 2514 142
rect 2422 98 2426 102
rect 2398 78 2402 82
rect 2062 68 2066 72
rect 2238 68 2242 72
rect 2278 68 2282 72
rect 1502 58 1506 62
rect 1814 58 1818 62
rect 2590 128 2594 132
rect 2614 118 2618 122
rect 2726 218 2730 222
rect 2630 128 2634 132
rect 2790 438 2794 442
rect 2862 1168 2866 1172
rect 2862 988 2866 992
rect 2854 938 2858 942
rect 2854 878 2858 882
rect 2862 858 2866 862
rect 2862 818 2866 822
rect 2862 788 2866 792
rect 2830 588 2834 592
rect 2806 458 2810 462
rect 2822 358 2826 362
rect 2998 1468 3002 1472
rect 2990 1368 2994 1372
rect 2894 1318 2898 1322
rect 2934 1338 2938 1342
rect 2918 1328 2922 1332
rect 2918 1278 2922 1282
rect 2926 1268 2930 1272
rect 2894 1258 2898 1262
rect 2910 1258 2914 1262
rect 2894 1248 2898 1252
rect 2910 1218 2914 1222
rect 2902 1098 2906 1102
rect 2886 988 2890 992
rect 2974 1298 2978 1302
rect 2974 1288 2978 1292
rect 2950 1218 2954 1222
rect 2958 1118 2962 1122
rect 2998 1158 3002 1162
rect 3222 3938 3226 3942
rect 3166 3518 3170 3522
rect 3166 3388 3170 3392
rect 3158 3078 3162 3082
rect 3190 3718 3194 3722
rect 3182 3378 3186 3382
rect 3294 3828 3298 3832
rect 3214 3658 3218 3662
rect 3654 4348 3658 4352
rect 3478 4338 3482 4342
rect 3550 4308 3554 4312
rect 3678 4298 3682 4302
rect 3670 4258 3674 4262
rect 3570 4203 3574 4207
rect 3577 4203 3578 4207
rect 3578 4203 3581 4207
rect 3710 4308 3714 4312
rect 3742 4268 3746 4272
rect 3726 4258 3730 4262
rect 3798 4278 3802 4282
rect 3798 4268 3802 4272
rect 3782 4258 3786 4262
rect 3570 4003 3574 4007
rect 3577 4003 3578 4007
rect 3578 4003 3581 4007
rect 3334 3758 3338 3762
rect 3230 3238 3234 3242
rect 3270 3268 3274 3272
rect 3050 2503 3054 2507
rect 3057 2503 3058 2507
rect 3058 2503 3061 2507
rect 3050 2303 3054 2307
rect 3057 2303 3058 2307
rect 3058 2303 3061 2307
rect 3134 2488 3138 2492
rect 3078 2318 3082 2322
rect 3070 2248 3074 2252
rect 3038 2218 3042 2222
rect 3030 2138 3034 2142
rect 3030 1968 3034 1972
rect 3110 2138 3114 2142
rect 3086 2128 3090 2132
rect 3094 2108 3098 2112
rect 3050 2103 3054 2107
rect 3057 2103 3058 2107
rect 3058 2103 3061 2107
rect 3078 2038 3082 2042
rect 3050 1903 3054 1907
rect 3057 1903 3058 1907
rect 3058 1903 3061 1907
rect 3014 1138 3018 1142
rect 2990 1128 2994 1132
rect 2998 1108 3002 1112
rect 2998 1078 3002 1082
rect 3006 1068 3010 1072
rect 2950 998 2954 1002
rect 2982 998 2986 1002
rect 2934 968 2938 972
rect 2966 948 2970 952
rect 2910 938 2914 942
rect 2886 898 2890 902
rect 2878 868 2882 872
rect 2966 868 2970 872
rect 2958 858 2962 862
rect 2934 758 2938 762
rect 2934 738 2938 742
rect 2934 728 2938 732
rect 2950 728 2954 732
rect 2918 678 2922 682
rect 2862 508 2866 512
rect 2862 458 2866 462
rect 2814 338 2818 342
rect 2806 318 2810 322
rect 2838 278 2842 282
rect 2862 208 2866 212
rect 2774 198 2778 202
rect 2902 558 2906 562
rect 2926 518 2930 522
rect 2998 918 3002 922
rect 2974 748 2978 752
rect 2966 708 2970 712
rect 2958 548 2962 552
rect 3050 1703 3054 1707
rect 3057 1703 3058 1707
rect 3058 1703 3061 1707
rect 3142 2418 3146 2422
rect 3166 2468 3170 2472
rect 3166 2278 3170 2282
rect 3166 2158 3170 2162
rect 3166 1848 3170 1852
rect 3102 1668 3106 1672
rect 3050 1503 3054 1507
rect 3057 1503 3058 1507
rect 3058 1503 3061 1507
rect 3062 1488 3066 1492
rect 3094 1468 3098 1472
rect 3078 1438 3082 1442
rect 3078 1418 3082 1422
rect 3062 1348 3066 1352
rect 3050 1303 3054 1307
rect 3057 1303 3058 1307
rect 3058 1303 3061 1307
rect 3078 1278 3082 1282
rect 3062 1258 3066 1262
rect 3126 1448 3130 1452
rect 3118 1408 3122 1412
rect 3134 1408 3138 1412
rect 3094 1318 3098 1322
rect 3102 1278 3106 1282
rect 3086 1218 3090 1222
rect 3102 1198 3106 1202
rect 3038 1178 3042 1182
rect 3110 1168 3114 1172
rect 3038 1128 3042 1132
rect 3050 1103 3054 1107
rect 3057 1103 3058 1107
rect 3058 1103 3061 1107
rect 3030 1058 3034 1062
rect 3046 918 3050 922
rect 3050 903 3054 907
rect 3057 903 3058 907
rect 3058 903 3061 907
rect 3086 968 3090 972
rect 3078 948 3082 952
rect 3102 918 3106 922
rect 3030 878 3034 882
rect 3038 878 3042 882
rect 3070 848 3074 852
rect 3022 758 3026 762
rect 3050 703 3054 707
rect 3057 703 3058 707
rect 3058 703 3061 707
rect 3070 648 3074 652
rect 3050 503 3054 507
rect 3057 503 3058 507
rect 3058 503 3061 507
rect 3038 488 3042 492
rect 3078 398 3082 402
rect 3014 358 3018 362
rect 2926 248 2930 252
rect 2974 238 2978 242
rect 2790 178 2794 182
rect 2758 148 2762 152
rect 2806 148 2810 152
rect 2782 108 2786 112
rect 2646 98 2650 102
rect 2814 98 2818 102
rect 2574 68 2578 72
rect 2846 68 2850 72
rect 2526 58 2530 62
rect 2926 158 2930 162
rect 2958 168 2962 172
rect 2974 168 2978 172
rect 2950 138 2954 142
rect 2974 148 2978 152
rect 3030 328 3034 332
rect 3102 898 3106 902
rect 3110 858 3114 862
rect 3142 1288 3146 1292
rect 3142 1268 3146 1272
rect 3142 1168 3146 1172
rect 3166 1738 3170 1742
rect 3246 2498 3250 2502
rect 3238 2368 3242 2372
rect 3190 1988 3194 1992
rect 3198 1988 3202 1992
rect 3182 1688 3186 1692
rect 3206 1678 3210 1682
rect 3182 1548 3186 1552
rect 3174 1538 3178 1542
rect 3158 1418 3162 1422
rect 3246 2148 3250 2152
rect 3222 2128 3226 2132
rect 3342 3518 3346 3522
rect 3350 3478 3354 3482
rect 3318 3398 3322 3402
rect 3326 3328 3330 3332
rect 3318 3318 3322 3322
rect 3302 3278 3306 3282
rect 3270 2438 3274 2442
rect 3262 2388 3266 2392
rect 3302 2878 3306 2882
rect 3342 3188 3346 3192
rect 3318 3128 3322 3132
rect 3382 3568 3386 3572
rect 3366 3438 3370 3442
rect 3366 3358 3370 3362
rect 3614 3948 3618 3952
rect 3814 4308 3818 4312
rect 3918 4358 3922 4362
rect 3838 4348 3842 4352
rect 3934 4338 3938 4342
rect 3854 4258 3858 4262
rect 3974 4338 3978 4342
rect 3902 4068 3906 4072
rect 3518 3838 3522 3842
rect 3570 3803 3574 3807
rect 3577 3803 3578 3807
rect 3578 3803 3581 3807
rect 3862 3948 3866 3952
rect 3430 3568 3434 3572
rect 3438 3348 3442 3352
rect 3350 2578 3354 2582
rect 3294 2378 3298 2382
rect 3278 2178 3282 2182
rect 3230 2088 3234 2092
rect 3438 2688 3442 2692
rect 3430 2618 3434 2622
rect 3390 2588 3394 2592
rect 3374 2568 3378 2572
rect 3382 2568 3386 2572
rect 3366 2318 3370 2322
rect 3374 2118 3378 2122
rect 3246 1958 3250 1962
rect 3406 2548 3410 2552
rect 3414 2408 3418 2412
rect 3414 2368 3418 2372
rect 3390 2188 3394 2192
rect 3478 3368 3482 3372
rect 3470 2538 3474 2542
rect 3462 2488 3466 2492
rect 3470 2268 3474 2272
rect 3454 2258 3458 2262
rect 3486 2458 3490 2462
rect 3534 3328 3538 3332
rect 3510 2168 3514 2172
rect 3502 2158 3506 2162
rect 3398 2148 3402 2152
rect 3494 2148 3498 2152
rect 3382 1978 3386 1982
rect 3518 1968 3522 1972
rect 3422 1938 3426 1942
rect 3366 1788 3370 1792
rect 3326 1778 3330 1782
rect 3294 1748 3298 1752
rect 3238 1718 3242 1722
rect 3214 1488 3218 1492
rect 3182 1438 3186 1442
rect 3174 1388 3178 1392
rect 3150 1148 3154 1152
rect 3166 1138 3170 1142
rect 3198 1348 3202 1352
rect 3230 1458 3234 1462
rect 3190 1338 3194 1342
rect 3222 1338 3226 1342
rect 3214 1328 3218 1332
rect 3206 1238 3210 1242
rect 3214 1218 3218 1222
rect 3230 1258 3234 1262
rect 3222 1188 3226 1192
rect 3190 1088 3194 1092
rect 3182 1078 3186 1082
rect 3158 1058 3162 1062
rect 3174 1058 3178 1062
rect 3198 1038 3202 1042
rect 3166 988 3170 992
rect 3182 948 3186 952
rect 3174 938 3178 942
rect 3182 908 3186 912
rect 3198 868 3202 872
rect 3222 1148 3226 1152
rect 3486 1678 3490 1682
rect 3358 1658 3362 1662
rect 3278 1428 3282 1432
rect 3270 1378 3274 1382
rect 3286 1318 3290 1322
rect 3350 1318 3354 1322
rect 3238 1018 3242 1022
rect 3222 938 3226 942
rect 3222 888 3226 892
rect 3142 738 3146 742
rect 3134 728 3138 732
rect 3118 548 3122 552
rect 3102 538 3106 542
rect 3158 778 3162 782
rect 3238 928 3242 932
rect 3238 918 3242 922
rect 3238 898 3242 902
rect 3214 748 3218 752
rect 3254 1288 3258 1292
rect 3254 1198 3258 1202
rect 3254 1098 3258 1102
rect 3270 1128 3274 1132
rect 3286 1158 3290 1162
rect 3302 1258 3306 1262
rect 3326 1168 3330 1172
rect 3310 1128 3314 1132
rect 3270 1028 3274 1032
rect 3278 1008 3282 1012
rect 3278 888 3282 892
rect 3334 1068 3338 1072
rect 3334 1018 3338 1022
rect 3334 968 3338 972
rect 3358 1228 3362 1232
rect 3406 1518 3410 1522
rect 3382 1458 3386 1462
rect 3358 1168 3362 1172
rect 3374 1078 3378 1082
rect 3358 1068 3362 1072
rect 3350 948 3354 952
rect 3326 798 3330 802
rect 3334 798 3338 802
rect 3302 788 3306 792
rect 3198 708 3202 712
rect 3166 688 3170 692
rect 3262 648 3266 652
rect 3390 998 3394 1002
rect 3494 1588 3498 1592
rect 3486 1578 3490 1582
rect 3454 1358 3458 1362
rect 3430 1228 3434 1232
rect 3446 1138 3450 1142
rect 3414 1128 3418 1132
rect 3438 1128 3442 1132
rect 3414 1008 3418 1012
rect 3390 928 3394 932
rect 3390 868 3394 872
rect 3390 758 3394 762
rect 3366 728 3370 732
rect 3382 718 3386 722
rect 3358 688 3362 692
rect 3438 978 3442 982
rect 3454 1118 3458 1122
rect 3446 878 3450 882
rect 3438 778 3442 782
rect 3422 738 3426 742
rect 3438 718 3442 722
rect 3050 303 3054 307
rect 3057 303 3058 307
rect 3058 303 3061 307
rect 3174 258 3178 262
rect 3198 258 3202 262
rect 3206 248 3210 252
rect 3174 228 3178 232
rect 3118 168 3122 172
rect 3038 138 3042 142
rect 3030 128 3034 132
rect 3110 118 3114 122
rect 3038 108 3042 112
rect 3050 103 3054 107
rect 3057 103 3058 107
rect 3058 103 3061 107
rect 3166 118 3170 122
rect 2990 88 2994 92
rect 3150 88 3154 92
rect 2998 78 3002 82
rect 3022 78 3026 82
rect 3118 68 3122 72
rect 3054 58 3058 62
rect 3078 58 3082 62
rect 3110 58 3114 62
rect 3214 188 3218 192
rect 3310 548 3314 552
rect 3398 538 3402 542
rect 3302 448 3306 452
rect 3294 338 3298 342
rect 3230 268 3234 272
rect 3230 198 3234 202
rect 3254 138 3258 142
rect 3278 178 3282 182
rect 3270 128 3274 132
rect 3254 98 3258 102
rect 3166 78 3170 82
rect 3246 68 3250 72
rect 3278 88 3282 92
rect 3294 298 3298 302
rect 3398 338 3402 342
rect 3478 1318 3482 1322
rect 3478 1278 3482 1282
rect 3486 1178 3490 1182
rect 3478 1138 3482 1142
rect 3478 1038 3482 1042
rect 3478 968 3482 972
rect 3478 858 3482 862
rect 3478 728 3482 732
rect 3570 3603 3574 3607
rect 3577 3603 3578 3607
rect 3578 3603 3581 3607
rect 3570 3403 3574 3407
rect 3577 3403 3578 3407
rect 3578 3403 3581 3407
rect 3570 3203 3574 3207
rect 3577 3203 3578 3207
rect 3578 3203 3581 3207
rect 3550 3068 3554 3072
rect 3570 3003 3574 3007
rect 3577 3003 3578 3007
rect 3578 3003 3581 3007
rect 3570 2803 3574 2807
rect 3577 2803 3578 2807
rect 3578 2803 3581 2807
rect 3570 2603 3574 2607
rect 3577 2603 3578 2607
rect 3578 2603 3581 2607
rect 3614 3518 3618 3522
rect 3590 2518 3594 2522
rect 3590 2498 3594 2502
rect 3638 3118 3642 3122
rect 3654 2548 3658 2552
rect 3630 2518 3634 2522
rect 3638 2468 3642 2472
rect 3598 2448 3602 2452
rect 3570 2403 3574 2407
rect 3577 2403 3578 2407
rect 3578 2403 3581 2407
rect 3606 2348 3610 2352
rect 3570 2203 3574 2207
rect 3577 2203 3578 2207
rect 3578 2203 3581 2207
rect 3646 2108 3650 2112
rect 3582 2028 3586 2032
rect 3570 2003 3574 2007
rect 3577 2003 3578 2007
rect 3578 2003 3581 2007
rect 3630 1998 3634 2002
rect 3570 1803 3574 1807
rect 3577 1803 3578 1807
rect 3578 1803 3581 1807
rect 3558 1758 3562 1762
rect 3630 1758 3634 1762
rect 3570 1603 3574 1607
rect 3577 1603 3578 1607
rect 3578 1603 3581 1607
rect 3526 1588 3530 1592
rect 3502 1548 3506 1552
rect 3606 1548 3610 1552
rect 3526 1538 3530 1542
rect 3606 1468 3610 1472
rect 3570 1403 3574 1407
rect 3577 1403 3578 1407
rect 3578 1403 3581 1407
rect 3510 1298 3514 1302
rect 3550 1268 3554 1272
rect 3590 1328 3594 1332
rect 3542 1248 3546 1252
rect 3582 1248 3586 1252
rect 3570 1203 3574 1207
rect 3577 1203 3578 1207
rect 3578 1203 3581 1207
rect 3558 1188 3562 1192
rect 3542 1158 3546 1162
rect 3590 1138 3594 1142
rect 3510 1108 3514 1112
rect 3526 1098 3530 1102
rect 3502 1038 3506 1042
rect 3510 1028 3514 1032
rect 3502 828 3506 832
rect 3534 1008 3538 1012
rect 3518 908 3522 912
rect 3566 1068 3570 1072
rect 3582 1068 3586 1072
rect 3582 1038 3586 1042
rect 3558 1028 3562 1032
rect 3570 1003 3574 1007
rect 3577 1003 3578 1007
rect 3578 1003 3581 1007
rect 3558 978 3562 982
rect 3550 918 3554 922
rect 3526 868 3530 872
rect 3502 818 3506 822
rect 3526 808 3530 812
rect 3494 528 3498 532
rect 3486 508 3490 512
rect 3454 388 3458 392
rect 3422 338 3426 342
rect 3390 278 3394 282
rect 3366 248 3370 252
rect 3318 218 3322 222
rect 3550 798 3554 802
rect 3566 938 3570 942
rect 3590 878 3594 882
rect 3574 838 3578 842
rect 3570 803 3574 807
rect 3577 803 3578 807
rect 3578 803 3581 807
rect 3566 738 3570 742
rect 3622 1268 3626 1272
rect 3614 1078 3618 1082
rect 3606 1038 3610 1042
rect 3654 1468 3658 1472
rect 3654 1318 3658 1322
rect 3654 1248 3658 1252
rect 3638 1238 3642 1242
rect 3638 1218 3642 1222
rect 3630 1148 3634 1152
rect 3630 1078 3634 1082
rect 3694 2628 3698 2632
rect 3702 2498 3706 2502
rect 3670 2058 3674 2062
rect 3686 2048 3690 2052
rect 3678 1978 3682 1982
rect 3726 2568 3730 2572
rect 3734 2538 3738 2542
rect 3758 2258 3762 2262
rect 4014 4278 4018 4282
rect 4150 4358 4154 4362
rect 3926 3868 3930 3872
rect 3942 3868 3946 3872
rect 4126 4338 4130 4342
rect 4082 4303 4086 4307
rect 4089 4303 4090 4307
rect 4090 4303 4093 4307
rect 4082 4103 4086 4107
rect 4089 4103 4090 4107
rect 4090 4103 4093 4107
rect 4126 4158 4130 4162
rect 4166 4348 4170 4352
rect 4142 4158 4146 4162
rect 4082 3903 4086 3907
rect 4089 3903 4090 3907
rect 4090 3903 4093 3907
rect 3934 3748 3938 3752
rect 4082 3703 4086 3707
rect 4089 3703 4090 3707
rect 4090 3703 4093 3707
rect 4142 4078 4146 4082
rect 4182 4318 4186 4322
rect 4350 4348 4354 4352
rect 4326 4338 4330 4342
rect 3806 3568 3810 3572
rect 3854 3458 3858 3462
rect 3854 2348 3858 2352
rect 3838 2318 3842 2322
rect 3870 2288 3874 2292
rect 3758 2038 3762 2042
rect 3702 1988 3706 1992
rect 3718 1968 3722 1972
rect 3694 1888 3698 1892
rect 3670 1838 3674 1842
rect 3678 1598 3682 1602
rect 3718 1948 3722 1952
rect 3790 2138 3794 2142
rect 3798 2048 3802 2052
rect 3798 2008 3802 2012
rect 3790 1918 3794 1922
rect 3870 2218 3874 2222
rect 3846 2038 3850 2042
rect 3854 1958 3858 1962
rect 3822 1928 3826 1932
rect 3878 2068 3882 2072
rect 3886 2048 3890 2052
rect 3894 1958 3898 1962
rect 3846 1818 3850 1822
rect 3822 1768 3826 1772
rect 3710 1688 3714 1692
rect 3694 1668 3698 1672
rect 3702 1638 3706 1642
rect 3678 1228 3682 1232
rect 3662 1178 3666 1182
rect 3670 1108 3674 1112
rect 3614 918 3618 922
rect 3694 1238 3698 1242
rect 3694 1028 3698 1032
rect 3678 888 3682 892
rect 3654 778 3658 782
rect 3622 728 3626 732
rect 3662 678 3666 682
rect 3654 668 3658 672
rect 3710 938 3714 942
rect 3622 628 3626 632
rect 3570 603 3574 607
rect 3577 603 3578 607
rect 3578 603 3581 607
rect 3686 618 3690 622
rect 3526 418 3530 422
rect 3570 403 3574 407
rect 3577 403 3578 407
rect 3578 403 3581 407
rect 3478 318 3482 322
rect 3558 308 3562 312
rect 3542 298 3546 302
rect 3502 258 3506 262
rect 3550 278 3554 282
rect 3486 208 3490 212
rect 3570 203 3574 207
rect 3577 203 3578 207
rect 3578 203 3581 207
rect 3462 178 3466 182
rect 3518 178 3522 182
rect 3558 178 3562 182
rect 3462 168 3466 172
rect 3446 148 3450 152
rect 3582 148 3586 152
rect 3574 138 3578 142
rect 3574 118 3578 122
rect 3374 108 3378 112
rect 3742 1458 3746 1462
rect 3750 1268 3754 1272
rect 3734 1188 3738 1192
rect 3838 1658 3842 1662
rect 3846 1648 3850 1652
rect 3814 1628 3818 1632
rect 3782 1438 3786 1442
rect 3806 1328 3810 1332
rect 3766 1118 3770 1122
rect 3774 1118 3778 1122
rect 3766 1108 3770 1112
rect 3758 1098 3762 1102
rect 3774 1088 3778 1092
rect 3766 1078 3770 1082
rect 3774 1068 3778 1072
rect 3806 968 3810 972
rect 3790 958 3794 962
rect 3758 918 3762 922
rect 3734 908 3738 912
rect 3726 868 3730 872
rect 3790 908 3794 912
rect 3798 868 3802 872
rect 3758 768 3762 772
rect 3774 748 3778 752
rect 3838 1348 3842 1352
rect 3830 1168 3834 1172
rect 3814 828 3818 832
rect 3654 338 3658 342
rect 3614 318 3618 322
rect 3670 318 3674 322
rect 3662 268 3666 272
rect 3702 568 3706 572
rect 3694 428 3698 432
rect 3702 358 3706 362
rect 3702 318 3706 322
rect 3718 358 3722 362
rect 3710 298 3714 302
rect 3654 218 3658 222
rect 3654 188 3658 192
rect 3662 188 3666 192
rect 3598 118 3602 122
rect 3606 108 3610 112
rect 3686 158 3690 162
rect 3614 88 3618 92
rect 3318 78 3322 82
rect 3598 78 3602 82
rect 3430 68 3434 72
rect 3518 68 3522 72
rect 3294 58 3298 62
rect 3742 488 3746 492
rect 3734 278 3738 282
rect 3782 608 3786 612
rect 4082 3503 4086 3507
rect 4089 3503 4090 3507
rect 4090 3503 4093 3507
rect 3934 3458 3938 3462
rect 3918 2478 3922 2482
rect 3926 2448 3930 2452
rect 4054 3138 4058 3142
rect 4038 2488 4042 2492
rect 3998 2458 4002 2462
rect 4014 2368 4018 2372
rect 4006 2348 4010 2352
rect 3966 2338 3970 2342
rect 4054 2428 4058 2432
rect 4082 3303 4086 3307
rect 4089 3303 4090 3307
rect 4090 3303 4093 3307
rect 4082 3103 4086 3107
rect 4089 3103 4090 3107
rect 4090 3103 4093 3107
rect 4082 2903 4086 2907
rect 4089 2903 4090 2907
rect 4090 2903 4093 2907
rect 4082 2703 4086 2707
rect 4089 2703 4090 2707
rect 4090 2703 4093 2707
rect 4082 2503 4086 2507
rect 4089 2503 4090 2507
rect 4090 2503 4093 2507
rect 4082 2303 4086 2307
rect 4089 2303 4090 2307
rect 4090 2303 4093 2307
rect 4094 2268 4098 2272
rect 4046 2178 4050 2182
rect 4082 2103 4086 2107
rect 4089 2103 4090 2107
rect 4090 2103 4093 2107
rect 4062 2048 4066 2052
rect 3966 1958 3970 1962
rect 3966 1918 3970 1922
rect 3918 1748 3922 1752
rect 3958 1868 3962 1872
rect 4046 1998 4050 2002
rect 4038 1948 4042 1952
rect 3982 1828 3986 1832
rect 3950 1668 3954 1672
rect 3966 1658 3970 1662
rect 3942 1508 3946 1512
rect 3902 1398 3906 1402
rect 3886 1358 3890 1362
rect 3902 1338 3906 1342
rect 3846 1278 3850 1282
rect 3846 1248 3850 1252
rect 3854 1248 3858 1252
rect 3886 1238 3890 1242
rect 3846 1088 3850 1092
rect 3830 938 3834 942
rect 3862 1048 3866 1052
rect 3878 1088 3882 1092
rect 3846 898 3850 902
rect 3862 868 3866 872
rect 3846 838 3850 842
rect 3830 788 3834 792
rect 3822 768 3826 772
rect 3822 528 3826 532
rect 3838 708 3842 712
rect 3822 438 3826 442
rect 3886 948 3890 952
rect 3894 948 3898 952
rect 3894 888 3898 892
rect 3910 1228 3914 1232
rect 3934 1168 3938 1172
rect 3918 1048 3922 1052
rect 3926 868 3930 872
rect 3934 858 3938 862
rect 3982 1628 3986 1632
rect 4014 1648 4018 1652
rect 3990 1528 3994 1532
rect 3990 1508 3994 1512
rect 3982 1438 3986 1442
rect 3958 1328 3962 1332
rect 3958 1318 3962 1322
rect 3974 1198 3978 1202
rect 3974 1178 3978 1182
rect 3966 1098 3970 1102
rect 3958 978 3962 982
rect 3910 768 3914 772
rect 3870 548 3874 552
rect 3910 458 3914 462
rect 3902 448 3906 452
rect 3806 368 3810 372
rect 3814 348 3818 352
rect 3790 298 3794 302
rect 3774 258 3778 262
rect 3766 238 3770 242
rect 3758 208 3762 212
rect 3702 58 3706 62
rect 3766 108 3770 112
rect 3782 98 3786 102
rect 3766 88 3770 92
rect 3838 278 3842 282
rect 3822 268 3826 272
rect 3814 248 3818 252
rect 3814 88 3818 92
rect 3790 58 3794 62
rect 3486 48 3490 52
rect 3830 148 3834 152
rect 3878 198 3882 202
rect 3854 108 3858 112
rect 3886 108 3890 112
rect 3854 88 3858 92
rect 3846 78 3850 82
rect 3870 78 3874 82
rect 3886 78 3890 82
rect 3902 248 3906 252
rect 3982 1088 3986 1092
rect 3982 958 3986 962
rect 4014 1468 4018 1472
rect 4082 1903 4086 1907
rect 4089 1903 4090 1907
rect 4090 1903 4093 1907
rect 4070 1878 4074 1882
rect 4030 1418 4034 1422
rect 4022 1358 4026 1362
rect 4030 1328 4034 1332
rect 4030 1298 4034 1302
rect 4030 1188 4034 1192
rect 3966 498 3970 502
rect 3974 468 3978 472
rect 3958 418 3962 422
rect 3950 378 3954 382
rect 3926 368 3930 372
rect 3918 268 3922 272
rect 3910 118 3914 122
rect 3870 68 3874 72
rect 3798 48 3802 52
rect 3014 38 3018 42
rect 3302 38 3306 42
rect 3854 38 3858 42
rect 3326 28 3330 32
rect 4006 1158 4010 1162
rect 4030 1138 4034 1142
rect 4038 1078 4042 1082
rect 4038 1048 4042 1052
rect 4046 1048 4050 1052
rect 4022 1038 4026 1042
rect 4038 1038 4042 1042
rect 4006 1018 4010 1022
rect 4006 848 4010 852
rect 4006 748 4010 752
rect 4038 818 4042 822
rect 4038 788 4042 792
rect 4030 748 4034 752
rect 4006 618 4010 622
rect 3998 338 4002 342
rect 3974 328 3978 332
rect 3990 318 3994 322
rect 3982 258 3986 262
rect 3942 218 3946 222
rect 3958 218 3962 222
rect 3966 208 3970 212
rect 3950 148 3954 152
rect 3958 148 3962 152
rect 3934 118 3938 122
rect 3950 108 3954 112
rect 3934 68 3938 72
rect 3974 128 3978 132
rect 4014 578 4018 582
rect 4022 508 4026 512
rect 4014 348 4018 352
rect 4014 318 4018 322
rect 4006 118 4010 122
rect 3974 68 3978 72
rect 3942 28 3946 32
rect 3958 28 3962 32
rect 3886 18 3890 22
rect 3902 18 3906 22
rect 4038 458 4042 462
rect 4030 108 4034 112
rect 4038 98 4042 102
rect 4082 1703 4086 1707
rect 4089 1703 4090 1707
rect 4090 1703 4093 1707
rect 4078 1578 4082 1582
rect 4082 1503 4086 1507
rect 4089 1503 4090 1507
rect 4090 1503 4093 1507
rect 4082 1303 4086 1307
rect 4089 1303 4090 1307
rect 4090 1303 4093 1307
rect 4094 1278 4098 1282
rect 4102 1178 4106 1182
rect 4070 1138 4074 1142
rect 4070 1108 4074 1112
rect 4082 1103 4086 1107
rect 4089 1103 4090 1107
rect 4090 1103 4093 1107
rect 4094 1048 4098 1052
rect 4142 2518 4146 2522
rect 4150 2358 4154 2362
rect 4158 2328 4162 2332
rect 4134 1868 4138 1872
rect 4166 1928 4170 1932
rect 4118 1518 4122 1522
rect 4158 1578 4162 1582
rect 4190 2538 4194 2542
rect 4182 2448 4186 2452
rect 4214 2418 4218 2422
rect 4198 2268 4202 2272
rect 4198 1978 4202 1982
rect 4182 1618 4186 1622
rect 4174 1568 4178 1572
rect 4174 1548 4178 1552
rect 4166 1498 4170 1502
rect 4158 1458 4162 1462
rect 4134 1228 4138 1232
rect 4134 1168 4138 1172
rect 4062 958 4066 962
rect 4094 948 4098 952
rect 4102 948 4106 952
rect 4070 918 4074 922
rect 4102 908 4106 912
rect 4082 903 4086 907
rect 4089 903 4090 907
rect 4090 903 4093 907
rect 4062 728 4066 732
rect 4062 718 4066 722
rect 4054 348 4058 352
rect 4054 228 4058 232
rect 4082 703 4086 707
rect 4089 703 4090 707
rect 4090 703 4093 707
rect 4078 578 4082 582
rect 4082 503 4086 507
rect 4089 503 4090 507
rect 4090 503 4093 507
rect 4070 338 4074 342
rect 4082 303 4086 307
rect 4089 303 4090 307
rect 4090 303 4093 307
rect 4070 298 4074 302
rect 4070 228 4074 232
rect 4094 248 4098 252
rect 4086 148 4090 152
rect 4062 128 4066 132
rect 4070 128 4074 132
rect 4082 103 4086 107
rect 4089 103 4090 107
rect 4090 103 4093 107
rect 4206 1568 4210 1572
rect 4174 1258 4178 1262
rect 4166 1188 4170 1192
rect 4158 1168 4162 1172
rect 4158 1118 4162 1122
rect 4182 1108 4186 1112
rect 4206 1338 4210 1342
rect 4198 1218 4202 1222
rect 4214 1088 4218 1092
rect 4190 998 4194 1002
rect 4158 858 4162 862
rect 4134 838 4138 842
rect 4118 628 4122 632
rect 4110 588 4114 592
rect 4110 518 4114 522
rect 4174 958 4178 962
rect 4190 938 4194 942
rect 4174 928 4178 932
rect 4166 828 4170 832
rect 4142 668 4146 672
rect 4134 638 4138 642
rect 4126 568 4130 572
rect 4126 548 4130 552
rect 4142 488 4146 492
rect 4126 198 4130 202
rect 4134 198 4138 202
rect 4046 68 4050 72
rect 4158 608 4162 612
rect 4214 878 4218 882
rect 4190 538 4194 542
rect 4182 398 4186 402
rect 4174 388 4178 392
rect 4150 178 4154 182
rect 4158 168 4162 172
rect 4206 798 4210 802
rect 4206 748 4210 752
rect 4262 3118 4266 3122
rect 4230 2588 4234 2592
rect 4358 4318 4362 4322
rect 4446 4358 4450 4362
rect 4486 4348 4490 4352
rect 4382 4258 4386 4262
rect 4318 3748 4322 3752
rect 4374 3938 4378 3942
rect 4326 2578 4330 2582
rect 4310 2568 4314 2572
rect 4310 2558 4314 2562
rect 4326 2528 4330 2532
rect 4342 2368 4346 2372
rect 4278 2348 4282 2352
rect 4310 2318 4314 2322
rect 4262 2228 4266 2232
rect 4254 2068 4258 2072
rect 4270 2058 4274 2062
rect 4254 1918 4258 1922
rect 4254 1888 4258 1892
rect 4238 1618 4242 1622
rect 4230 1608 4234 1612
rect 4230 1598 4234 1602
rect 4238 1568 4242 1572
rect 4230 1548 4234 1552
rect 4238 1468 4242 1472
rect 4230 1448 4234 1452
rect 4262 1568 4266 1572
rect 4270 1378 4274 1382
rect 4262 1368 4266 1372
rect 4238 1358 4242 1362
rect 4238 1198 4242 1202
rect 4254 1158 4258 1162
rect 4246 1138 4250 1142
rect 4230 1128 4234 1132
rect 4238 1078 4242 1082
rect 4230 918 4234 922
rect 4222 618 4226 622
rect 4238 678 4242 682
rect 4214 328 4218 332
rect 4230 558 4234 562
rect 4238 558 4242 562
rect 4238 468 4242 472
rect 4262 1038 4266 1042
rect 4270 948 4274 952
rect 4334 2328 4338 2332
rect 4342 1928 4346 1932
rect 4366 2358 4370 2362
rect 4382 2338 4386 2342
rect 4374 1788 4378 1792
rect 4358 1688 4362 1692
rect 4374 1678 4378 1682
rect 4302 1638 4306 1642
rect 4406 1968 4410 1972
rect 4406 1648 4410 1652
rect 4390 1588 4394 1592
rect 4398 1578 4402 1582
rect 4406 1548 4410 1552
rect 4310 1448 4314 1452
rect 4294 1248 4298 1252
rect 4302 1008 4306 1012
rect 4294 928 4298 932
rect 4270 858 4274 862
rect 4278 848 4282 852
rect 4294 848 4298 852
rect 4390 1488 4394 1492
rect 4350 1438 4354 1442
rect 4350 1388 4354 1392
rect 4342 1088 4346 1092
rect 4262 748 4266 752
rect 4278 728 4282 732
rect 4270 528 4274 532
rect 4198 258 4202 262
rect 4214 228 4218 232
rect 4182 178 4186 182
rect 4190 168 4194 172
rect 4222 218 4226 222
rect 4254 198 4258 202
rect 4238 158 4242 162
rect 4206 148 4210 152
rect 4222 148 4226 152
rect 4134 68 4138 72
rect 4174 58 4178 62
rect 4110 28 4114 32
rect 4262 128 4266 132
rect 4310 548 4314 552
rect 4302 418 4306 422
rect 4278 258 4282 262
rect 4294 238 4298 242
rect 4230 78 4234 82
rect 4254 78 4258 82
rect 4270 58 4274 62
rect 4406 1358 4410 1362
rect 4462 4328 4466 4332
rect 4462 4298 4466 4302
rect 4486 4258 4490 4262
rect 4454 4108 4458 4112
rect 4478 3938 4482 3942
rect 4454 3468 4458 3472
rect 4422 1728 4426 1732
rect 4414 1198 4418 1202
rect 4438 1178 4442 1182
rect 4406 1048 4410 1052
rect 4382 988 4386 992
rect 4358 968 4362 972
rect 4358 958 4362 962
rect 4350 578 4354 582
rect 4318 288 4322 292
rect 4318 188 4322 192
rect 4310 178 4314 182
rect 4350 138 4354 142
rect 4342 118 4346 122
rect 4350 108 4354 112
rect 4374 738 4378 742
rect 4374 718 4378 722
rect 4398 918 4402 922
rect 4406 858 4410 862
rect 4406 278 4410 282
rect 4430 1068 4434 1072
rect 4422 488 4426 492
rect 4422 468 4426 472
rect 4438 998 4442 1002
rect 4438 878 4442 882
rect 4454 1918 4458 1922
rect 4462 1288 4466 1292
rect 4454 1168 4458 1172
rect 4462 1068 4466 1072
rect 4454 1048 4458 1052
rect 4462 928 4466 932
rect 4454 448 4458 452
rect 4438 88 4442 92
rect 4478 2798 4482 2802
rect 4510 3828 4514 3832
rect 4510 2708 4514 2712
rect 4510 2348 4514 2352
rect 4510 2338 4514 2342
rect 4478 1458 4482 1462
rect 4502 2128 4506 2132
rect 4550 4298 4554 4302
rect 4534 4088 4538 4092
rect 4566 4248 4570 4252
rect 4558 3138 4562 3142
rect 4542 2548 4546 2552
rect 4526 2378 4530 2382
rect 4542 2378 4546 2382
rect 4526 2368 4530 2372
rect 4518 2258 4522 2262
rect 4518 1648 4522 1652
rect 4526 1638 4530 1642
rect 4486 1398 4490 1402
rect 4486 1368 4490 1372
rect 4494 1348 4498 1352
rect 4590 3248 4594 3252
rect 4566 2318 4570 2322
rect 4558 2068 4562 2072
rect 4574 2038 4578 2042
rect 4566 1528 4570 1532
rect 4558 1498 4562 1502
rect 4558 1458 4562 1462
rect 4574 1398 4578 1402
rect 4542 948 4546 952
rect 4526 908 4530 912
rect 4486 838 4490 842
rect 4518 788 4522 792
rect 4518 428 4522 432
rect 4502 368 4506 372
rect 4486 278 4490 282
rect 4470 78 4474 82
rect 4542 768 4546 772
rect 4558 928 4562 932
rect 4566 658 4570 662
rect 4574 538 4578 542
rect 4574 478 4578 482
rect 4590 1678 4594 1682
rect 4590 1268 4594 1272
rect 4542 328 4546 332
rect 4542 158 4546 162
rect 4510 68 4514 72
rect 3966 8 3970 12
rect 4078 8 4082 12
rect 4534 8 4538 12
rect 498 3 502 7
rect 505 3 506 7
rect 506 3 509 7
rect 1522 3 1526 7
rect 1529 3 1530 7
rect 1530 3 1533 7
rect 2546 3 2550 7
rect 2553 3 2554 7
rect 2554 3 2557 7
rect 3570 3 3574 7
rect 3577 3 3578 7
rect 3578 3 3581 7
<< metal5 >>
rect 502 4403 505 4407
rect 501 4402 506 4403
rect 511 4402 512 4407
rect 1526 4403 1529 4407
rect 1525 4402 1530 4403
rect 1535 4402 1536 4407
rect 2550 4403 2553 4407
rect 2549 4402 2554 4403
rect 2559 4402 2560 4407
rect 3574 4403 3577 4407
rect 3573 4402 3578 4403
rect 3583 4402 3584 4407
rect 4010 4398 4254 4401
rect 3922 4358 4150 4361
rect 4446 4352 4449 4358
rect 3658 4348 3838 4351
rect 3842 4348 3977 4351
rect 4170 4348 4350 4351
rect 3974 4342 3977 4348
rect 4482 4348 4486 4351
rect 1762 4338 3230 4341
rect 3482 4338 3934 4341
rect 4130 4338 4326 4341
rect 4386 4328 4462 4331
rect 4186 4318 4358 4321
rect 3554 4308 3710 4311
rect 4550 4308 4573 4311
rect 1006 4303 1009 4307
rect 1005 4302 1010 4303
rect 1015 4302 1016 4307
rect 2030 4303 2033 4307
rect 2029 4302 2034 4303
rect 2039 4302 2040 4307
rect 3054 4303 3057 4307
rect 3053 4302 3058 4303
rect 3063 4302 3064 4307
rect 3814 4301 3817 4308
rect 4086 4303 4089 4307
rect 4085 4302 4090 4303
rect 4095 4302 4096 4307
rect 4550 4302 4553 4308
rect 3682 4298 3817 4301
rect 4462 4292 4465 4298
rect 2090 4288 2262 4291
rect 3802 4278 4014 4281
rect 866 4268 1102 4271
rect 1570 4268 1822 4271
rect 2482 4268 2838 4271
rect 3746 4268 3798 4271
rect 1130 4258 1198 4261
rect 1250 4258 2009 4261
rect 2178 4258 2398 4261
rect 3674 4258 3726 4261
rect 3786 4258 3854 4261
rect 4386 4258 4486 4261
rect 4490 4258 4569 4261
rect 2006 4252 2009 4258
rect 4566 4252 4569 4258
rect 530 4248 806 4251
rect 2162 4248 2270 4251
rect 2514 4248 2654 4251
rect 474 4238 942 4241
rect 1474 4238 1990 4241
rect 682 4228 1934 4231
rect 1962 4228 2414 4231
rect 502 4203 505 4207
rect 501 4202 506 4203
rect 511 4202 512 4207
rect 1526 4203 1529 4207
rect 1525 4202 1530 4203
rect 1535 4202 1536 4207
rect 2550 4203 2553 4207
rect 2549 4202 2554 4203
rect 2559 4202 2560 4207
rect 3574 4203 3577 4207
rect 3573 4202 3578 4203
rect 3583 4202 3584 4207
rect 1698 4188 2758 4191
rect 2242 4178 2430 4181
rect 1314 4158 1438 4161
rect 1802 4158 2686 4161
rect 4130 4158 4142 4161
rect 274 4148 638 4151
rect 1050 4148 1910 4151
rect 1914 4148 2254 4151
rect 1770 4138 2350 4141
rect 1258 4128 2894 4131
rect 1978 4118 2358 4121
rect 4458 4108 4541 4111
rect 1006 4103 1009 4107
rect 1005 4102 1010 4103
rect 1015 4102 1016 4107
rect 2030 4103 2033 4107
rect 2029 4102 2034 4103
rect 2039 4102 2040 4107
rect 3054 4103 3057 4107
rect 3053 4102 3058 4103
rect 3063 4102 3064 4107
rect 4086 4103 4089 4107
rect 4085 4102 4090 4103
rect 4095 4102 4096 4107
rect 1402 4088 2662 4091
rect 4538 4088 4557 4091
rect 1842 4078 2438 4081
rect 2442 4078 2630 4081
rect 2634 4068 2830 4071
rect 4142 4071 4145 4078
rect 3906 4068 4145 4071
rect 2394 4058 2470 4061
rect 2594 4058 2702 4061
rect 2506 4048 2622 4051
rect 502 4003 505 4007
rect 501 4002 506 4003
rect 511 4002 512 4007
rect 1526 4003 1529 4007
rect 1525 4002 1530 4003
rect 1535 4002 1536 4007
rect 2550 4003 2553 4007
rect 2549 4002 2554 4003
rect 2559 4002 2560 4007
rect 3574 4003 3577 4007
rect 3573 4002 3578 4003
rect 3583 4002 3584 4007
rect 1530 3958 1814 3961
rect 2182 3951 2185 3958
rect 938 3948 2566 3951
rect 3618 3948 3862 3951
rect 2410 3938 3222 3941
rect 4378 3938 4478 3941
rect 1006 3903 1009 3907
rect 1005 3902 1010 3903
rect 1015 3902 1016 3907
rect 2030 3903 2033 3907
rect 2029 3902 2034 3903
rect 2039 3902 2040 3907
rect 3054 3903 3057 3907
rect 3053 3902 3058 3903
rect 3063 3902 3064 3907
rect 4086 3903 4089 3907
rect 4085 3902 4090 3903
rect 4095 3902 4096 3907
rect 2106 3878 2486 3881
rect 2098 3868 2246 3871
rect 2818 3868 2878 3871
rect 3930 3868 3942 3871
rect 2498 3858 2566 3861
rect 2554 3848 3070 3851
rect 1354 3838 3518 3841
rect 1106 3828 3294 3831
rect 4510 3822 4513 3828
rect 502 3803 505 3807
rect 501 3802 506 3803
rect 511 3802 512 3807
rect 1526 3803 1529 3807
rect 1525 3802 1530 3803
rect 1535 3802 1536 3807
rect 2550 3803 2553 3807
rect 2549 3802 2554 3803
rect 2559 3802 2560 3807
rect 3574 3803 3577 3807
rect 3573 3802 3578 3803
rect 3583 3802 3584 3807
rect 2538 3758 3334 3761
rect 3938 3748 4318 3751
rect 786 3738 2062 3741
rect 2714 3718 3190 3721
rect 2334 3712 2337 3718
rect 1006 3703 1009 3707
rect 1005 3702 1010 3703
rect 1015 3702 1016 3707
rect 2030 3703 2033 3707
rect 2029 3702 2034 3703
rect 2039 3702 2040 3707
rect 3054 3703 3057 3707
rect 3053 3702 3058 3703
rect 3063 3702 3064 3707
rect 4086 3703 4089 3707
rect 4085 3702 4090 3703
rect 4095 3702 4096 3707
rect 2274 3688 2710 3691
rect 2370 3678 2886 3681
rect 2946 3668 3110 3671
rect 994 3658 2126 3661
rect 2330 3658 2558 3661
rect 2698 3658 2838 3661
rect 2866 3658 3214 3661
rect 2474 3648 2950 3651
rect 502 3603 505 3607
rect 501 3602 506 3603
rect 511 3602 512 3607
rect 1526 3603 1529 3607
rect 1525 3602 1530 3603
rect 1535 3602 1536 3607
rect 2550 3603 2553 3607
rect 2549 3602 2554 3603
rect 2559 3602 2560 3607
rect 3574 3603 3577 3607
rect 3573 3602 3578 3603
rect 3583 3602 3584 3607
rect 2330 3588 2502 3591
rect 2282 3568 2478 3571
rect 2514 3568 3382 3571
rect 3434 3568 3806 3571
rect 1818 3558 2158 3561
rect 1506 3548 1974 3551
rect 1522 3538 2006 3541
rect 2010 3518 2422 3521
rect 2714 3518 3166 3521
rect 3346 3518 3614 3521
rect 2654 3512 2657 3518
rect 1006 3503 1009 3507
rect 1005 3502 1010 3503
rect 1015 3502 1016 3507
rect 2030 3503 2033 3507
rect 2029 3502 2034 3503
rect 2039 3502 2040 3507
rect 3054 3503 3057 3507
rect 3053 3502 3058 3503
rect 3063 3502 3064 3507
rect 4086 3503 4089 3507
rect 4085 3502 4090 3503
rect 4095 3502 4096 3507
rect 2802 3488 3118 3491
rect 2890 3478 3350 3481
rect 1954 3468 2030 3471
rect 2626 3468 2958 3471
rect 2994 3468 3086 3471
rect 4434 3468 4454 3471
rect 2650 3458 2798 3461
rect 3026 3458 3094 3461
rect 3858 3458 3934 3461
rect 2934 3451 2937 3458
rect 2738 3448 2937 3451
rect 2338 3438 2814 3441
rect 2834 3438 3366 3441
rect 2706 3428 3094 3431
rect 2354 3418 2782 3421
rect 2730 3408 3006 3411
rect 502 3403 505 3407
rect 501 3402 506 3403
rect 511 3402 512 3407
rect 1526 3403 1529 3407
rect 1525 3402 1530 3403
rect 1535 3402 1536 3407
rect 2550 3403 2553 3407
rect 2549 3402 2554 3403
rect 2559 3402 2560 3407
rect 3574 3403 3577 3407
rect 3573 3402 3578 3403
rect 3583 3402 3584 3407
rect 2362 3398 2526 3401
rect 2682 3398 3318 3401
rect 1234 3388 1318 3391
rect 1322 3388 2414 3391
rect 2434 3388 2829 3391
rect 2858 3388 3166 3391
rect 2354 3378 2918 3381
rect 2938 3378 3182 3381
rect 2346 3368 2878 3371
rect 2886 3368 3478 3371
rect 1922 3358 2302 3361
rect 2886 3361 2889 3368
rect 2522 3358 2889 3361
rect 2978 3358 3366 3361
rect 1778 3348 2110 3351
rect 3002 3348 3438 3351
rect 2298 3338 2333 3341
rect 2914 3338 2966 3341
rect 2522 3328 2525 3331
rect 3330 3328 3534 3331
rect 2386 3318 2406 3321
rect 2562 3318 3318 3321
rect 2282 3308 2390 3311
rect 1006 3303 1009 3307
rect 1005 3302 1010 3303
rect 1015 3302 1016 3307
rect 2030 3303 2033 3307
rect 2029 3302 2034 3303
rect 2039 3302 2040 3307
rect 3054 3303 3057 3307
rect 3053 3302 3058 3303
rect 3063 3302 3064 3307
rect 4086 3303 4089 3307
rect 4085 3302 4090 3303
rect 4095 3302 4096 3307
rect 2362 3298 2710 3301
rect 1914 3288 2278 3291
rect 930 3278 1166 3281
rect 1170 3278 2182 3281
rect 2218 3278 3110 3281
rect 306 3268 326 3271
rect 330 3268 494 3271
rect 970 3268 2574 3271
rect 3302 3271 3305 3278
rect 3274 3268 3305 3271
rect 2106 3258 2534 3261
rect 1786 3248 2262 3251
rect 4590 3242 4593 3248
rect 1490 3238 3230 3241
rect 2354 3218 2870 3221
rect 502 3203 505 3207
rect 501 3202 506 3203
rect 511 3202 512 3207
rect 1526 3203 1529 3207
rect 1525 3202 1530 3203
rect 1535 3202 1536 3207
rect 2550 3203 2553 3207
rect 2549 3202 2554 3203
rect 2559 3202 2560 3207
rect 3574 3203 3577 3207
rect 3573 3202 3578 3203
rect 3583 3202 3584 3207
rect 2170 3188 3342 3191
rect 2202 3178 2462 3181
rect 2382 3161 2385 3168
rect 2226 3158 2385 3161
rect 2646 3161 2649 3168
rect 2646 3158 2653 3161
rect 2674 3158 2878 3161
rect 1618 3138 2086 3141
rect 4058 3138 4558 3141
rect 2882 3128 3318 3131
rect 3642 3118 4262 3121
rect 2322 3108 2742 3111
rect 1006 3103 1009 3107
rect 1005 3102 1010 3103
rect 1015 3102 1016 3107
rect 2030 3103 2033 3107
rect 2029 3102 2034 3103
rect 2039 3102 2040 3107
rect 3054 3103 3057 3107
rect 3053 3102 3058 3103
rect 3063 3102 3064 3107
rect 4086 3103 4089 3107
rect 4085 3102 4090 3103
rect 4095 3102 4096 3107
rect 2050 3098 2438 3101
rect 1306 3088 1574 3091
rect 1674 3088 1878 3091
rect 914 3078 2262 3081
rect 2490 3078 3158 3081
rect 2226 3068 3550 3071
rect 1850 3058 2318 3061
rect 2050 3038 2342 3041
rect 502 3003 505 3007
rect 501 3002 506 3003
rect 511 3002 512 3007
rect 1526 3003 1529 3007
rect 1525 3002 1530 3003
rect 1535 3002 1536 3007
rect 2550 3003 2553 3007
rect 2549 3002 2554 3003
rect 2559 3002 2560 3007
rect 3574 3003 3577 3007
rect 3573 3002 3578 3003
rect 3583 3002 3584 3007
rect 2002 2958 2230 2961
rect 1546 2948 2022 2951
rect 2242 2948 2518 2951
rect 2018 2938 2142 2941
rect 2290 2938 2494 2941
rect 1226 2918 1254 2921
rect 1258 2918 2846 2921
rect 1006 2903 1009 2907
rect 1005 2902 1010 2903
rect 1015 2902 1016 2907
rect 2030 2903 2033 2907
rect 2029 2902 2034 2903
rect 2039 2902 2040 2907
rect 3054 2903 3057 2907
rect 3053 2902 3058 2903
rect 3063 2902 3064 2907
rect 4086 2903 4089 2907
rect 4085 2902 4090 2903
rect 4095 2902 4096 2907
rect 1922 2888 2046 2891
rect 2410 2888 2686 2891
rect 2314 2878 3302 2881
rect 3306 2878 3949 2881
rect 2506 2868 2870 2871
rect 1042 2858 1574 2861
rect 1578 2858 2758 2861
rect 502 2803 505 2807
rect 501 2802 506 2803
rect 511 2802 512 2807
rect 1526 2803 1529 2807
rect 1525 2802 1530 2803
rect 1535 2802 1536 2807
rect 2550 2803 2553 2807
rect 2549 2802 2554 2803
rect 2559 2802 2560 2807
rect 3574 2803 3577 2807
rect 3573 2802 3578 2803
rect 3583 2802 3584 2807
rect 4478 2802 4481 2807
rect 1906 2778 2097 2781
rect 2094 2772 2097 2778
rect 650 2748 886 2751
rect 1426 2748 1670 2751
rect 1674 2748 2910 2751
rect 2538 2718 3086 2721
rect 4482 2708 4510 2711
rect 1006 2703 1009 2707
rect 1005 2702 1010 2703
rect 1015 2702 1016 2707
rect 2030 2703 2033 2707
rect 2029 2702 2034 2703
rect 2039 2702 2040 2707
rect 3054 2703 3057 2707
rect 3053 2702 3058 2703
rect 3063 2702 3064 2707
rect 4086 2703 4089 2707
rect 4085 2702 4090 2703
rect 4095 2702 4096 2707
rect 898 2688 1054 2691
rect 1058 2688 1102 2691
rect 1106 2688 3438 2691
rect 658 2678 790 2681
rect 2194 2678 2870 2681
rect 1770 2668 2390 2671
rect 754 2658 822 2661
rect 1338 2658 1470 2661
rect 1474 2658 2846 2661
rect 618 2648 710 2651
rect 2266 2648 2670 2651
rect 2778 2628 3694 2631
rect 1026 2618 1270 2621
rect 1274 2618 1382 2621
rect 1386 2618 3430 2621
rect 502 2603 505 2607
rect 501 2602 506 2603
rect 511 2602 512 2607
rect 1526 2603 1529 2607
rect 1525 2602 1530 2603
rect 1535 2602 1536 2607
rect 2550 2603 2553 2607
rect 2549 2602 2554 2603
rect 2559 2602 2560 2607
rect 3574 2603 3577 2607
rect 3573 2602 3578 2603
rect 3583 2602 3584 2607
rect 3394 2588 4230 2591
rect 3354 2578 4326 2581
rect 2834 2568 3374 2571
rect 3386 2568 3726 2571
rect 3810 2568 4310 2571
rect 2754 2558 4310 2561
rect 2130 2548 2134 2551
rect 3410 2548 3654 2551
rect 3858 2548 4542 2551
rect 2466 2538 3470 2541
rect 3738 2538 4190 2541
rect 2818 2528 3741 2531
rect 3746 2528 4326 2531
rect 1458 2518 2838 2521
rect 2962 2518 3590 2521
rect 3634 2518 3661 2521
rect 3666 2518 4142 2521
rect 1006 2503 1009 2507
rect 1005 2502 1010 2503
rect 1015 2502 1016 2507
rect 2030 2503 2033 2507
rect 2029 2502 2034 2503
rect 2039 2502 2040 2507
rect 3054 2503 3057 2507
rect 3053 2502 3058 2503
rect 3063 2502 3064 2507
rect 4086 2503 4089 2507
rect 4085 2502 4090 2503
rect 4095 2502 4096 2507
rect 3250 2498 3590 2501
rect 3594 2498 3702 2501
rect 1042 2488 2334 2491
rect 2682 2488 3134 2491
rect 3466 2488 4038 2491
rect 1010 2478 1078 2481
rect 1082 2478 2590 2481
rect 2874 2478 3918 2481
rect 918 2471 921 2478
rect 918 2468 1190 2471
rect 1210 2468 1422 2471
rect 1426 2468 1806 2471
rect 1810 2468 2990 2471
rect 3170 2468 3638 2471
rect 2514 2458 2862 2461
rect 3490 2458 3998 2461
rect 2274 2448 3598 2451
rect 3930 2448 4182 2451
rect 1370 2438 1638 2441
rect 1642 2438 3270 2441
rect 1546 2428 4054 2431
rect 2082 2418 2998 2421
rect 3146 2418 4214 2421
rect 1570 2408 2302 2411
rect 2658 2408 3414 2411
rect 502 2403 505 2407
rect 501 2402 506 2403
rect 511 2402 512 2407
rect 1526 2403 1529 2407
rect 1525 2402 1530 2403
rect 1535 2402 1536 2407
rect 2550 2403 2553 2407
rect 2549 2402 2554 2403
rect 2559 2402 2560 2407
rect 3574 2403 3577 2407
rect 3573 2402 3578 2403
rect 3583 2402 3584 2407
rect 2666 2398 2982 2401
rect 2250 2388 2926 2391
rect 2978 2388 3262 2391
rect 2298 2378 3294 2381
rect 4530 2378 4542 2381
rect 1414 2361 1417 2368
rect 2370 2368 2374 2371
rect 2834 2368 3238 2371
rect 3418 2368 4014 2371
rect 4346 2368 4526 2371
rect 1414 2358 1550 2361
rect 1554 2358 1902 2361
rect 1906 2358 2758 2361
rect 2898 2358 3725 2361
rect 4154 2358 4366 2361
rect 2890 2348 3606 2351
rect 3858 2348 4006 2351
rect 4282 2348 4510 2351
rect 938 2338 1270 2341
rect 2730 2338 3645 2341
rect 3650 2338 3966 2341
rect 4274 2338 4382 2341
rect 4450 2338 4510 2341
rect 906 2328 942 2331
rect 2370 2328 2982 2331
rect 4162 2328 4334 2331
rect 2018 2318 3078 2321
rect 3370 2318 3838 2321
rect 4314 2318 4566 2321
rect 1006 2303 1009 2307
rect 1005 2302 1010 2303
rect 1015 2302 1016 2307
rect 2030 2303 2033 2307
rect 2029 2302 2034 2303
rect 2039 2302 2040 2307
rect 3054 2303 3057 2307
rect 3053 2302 3058 2303
rect 3063 2302 3064 2307
rect 4086 2303 4089 2307
rect 4085 2302 4090 2303
rect 4095 2302 4096 2307
rect 2850 2288 2902 2291
rect 2906 2288 3870 2291
rect 2242 2278 2782 2281
rect 2938 2278 3166 2281
rect 1594 2268 2662 2271
rect 2754 2268 2937 2271
rect 2934 2262 2937 2268
rect 4098 2268 4198 2271
rect 2386 2258 2902 2261
rect 2938 2258 3454 2261
rect 3470 2261 3473 2268
rect 3470 2258 3758 2261
rect 4522 2258 4525 2261
rect 2010 2248 3070 2251
rect 1602 2238 2678 2241
rect 2426 2228 2894 2231
rect 4178 2228 4262 2231
rect 3042 2218 3870 2221
rect 502 2203 505 2207
rect 501 2202 506 2203
rect 511 2202 512 2207
rect 1526 2203 1529 2207
rect 1525 2202 1530 2203
rect 1535 2202 1536 2207
rect 2550 2203 2553 2207
rect 2549 2202 2554 2203
rect 2559 2202 2560 2207
rect 3574 2203 3577 2207
rect 3573 2202 3578 2203
rect 3583 2202 3584 2207
rect 1698 2188 3390 2191
rect 2314 2178 3278 2181
rect 3282 2178 4046 2181
rect 1778 2168 3510 2171
rect 2594 2158 2654 2161
rect 3170 2158 3502 2161
rect 450 2148 798 2151
rect 2218 2148 2950 2151
rect 2978 2148 3246 2151
rect 3402 2148 3494 2151
rect 858 2138 1542 2141
rect 3034 2138 3110 2141
rect 3794 2138 4505 2141
rect 4502 2132 4505 2138
rect 650 2128 1334 2131
rect 1738 2128 2702 2131
rect 3090 2128 3222 2131
rect 994 2118 1510 2121
rect 2018 2118 3374 2121
rect 3098 2108 3646 2111
rect 1006 2103 1009 2107
rect 1005 2102 1010 2103
rect 1015 2102 1016 2107
rect 2030 2103 2033 2107
rect 2029 2102 2034 2103
rect 2039 2102 2040 2107
rect 3054 2103 3057 2107
rect 3053 2102 3058 2103
rect 3063 2102 3064 2107
rect 4086 2103 4089 2107
rect 4085 2102 4090 2103
rect 4095 2102 4096 2107
rect 2242 2098 2726 2101
rect 2674 2088 3230 2091
rect 482 2078 2334 2081
rect 2410 2078 2590 2081
rect 290 2068 318 2071
rect 322 2068 329 2071
rect 1010 2068 1102 2071
rect 2418 2068 2438 2071
rect 2530 2068 3878 2071
rect 4258 2068 4558 2071
rect 1074 2058 1774 2061
rect 2306 2058 2438 2061
rect 3674 2058 4270 2061
rect 2258 2048 2406 2051
rect 2826 2048 3686 2051
rect 3758 2048 3798 2051
rect 3890 2048 4062 2051
rect 3758 2042 3761 2048
rect 1978 2038 3078 2041
rect 3850 2038 4574 2041
rect 898 2028 1894 2031
rect 1898 2028 2054 2031
rect 2162 2028 3582 2031
rect 2362 2018 3801 2021
rect 3798 2012 3801 2018
rect 1698 2008 2254 2011
rect 502 2003 505 2007
rect 501 2002 506 2003
rect 511 2002 512 2007
rect 1526 2003 1529 2007
rect 1525 2002 1530 2003
rect 1535 2002 1536 2007
rect 2550 2003 2553 2007
rect 2549 2002 2554 2003
rect 2559 2002 2560 2007
rect 3574 2003 3577 2007
rect 3573 2002 3578 2003
rect 3583 2002 3584 2007
rect 1682 1998 1846 2001
rect 3634 1998 4046 2001
rect 874 1988 1910 1991
rect 2306 1988 3190 1991
rect 3202 1988 3702 1991
rect 1770 1978 3382 1981
rect 3682 1978 4198 1981
rect 394 1968 918 1971
rect 3034 1968 3518 1971
rect 3722 1968 4406 1971
rect 1774 1961 1777 1968
rect 1774 1958 2054 1961
rect 2378 1958 2681 1961
rect 3250 1958 3854 1961
rect 3898 1958 3966 1961
rect 2678 1952 2681 1958
rect 1282 1948 1838 1951
rect 3722 1948 4038 1951
rect 322 1938 918 1941
rect 1786 1938 2150 1941
rect 2706 1938 3422 1941
rect 1826 1928 2190 1931
rect 2498 1928 2934 1931
rect 3826 1928 4166 1931
rect 4346 1928 4457 1931
rect 4454 1922 4457 1928
rect 1934 1918 1942 1921
rect 1946 1918 2238 1921
rect 2322 1918 3790 1921
rect 3970 1918 4254 1921
rect 1006 1903 1009 1907
rect 1005 1902 1010 1903
rect 1015 1902 1016 1907
rect 2030 1903 2033 1907
rect 2029 1902 2034 1903
rect 2039 1902 2040 1907
rect 3054 1903 3057 1907
rect 3053 1902 3058 1903
rect 3063 1902 3064 1907
rect 4086 1903 4089 1907
rect 4085 1902 4090 1903
rect 4095 1902 4096 1907
rect 2338 1888 2750 1891
rect 3698 1888 3709 1891
rect 1566 1881 1569 1888
rect 970 1878 1569 1881
rect 1746 1878 2190 1881
rect 4254 1881 4257 1888
rect 4074 1878 4257 1881
rect 1138 1868 2366 1871
rect 2370 1868 2630 1871
rect 2666 1868 2702 1871
rect 3962 1868 4134 1871
rect 1690 1858 1758 1861
rect 1794 1858 2998 1861
rect 2178 1848 3166 1851
rect 2162 1838 3670 1841
rect 1506 1828 1846 1831
rect 1850 1828 2118 1831
rect 2938 1828 3982 1831
rect 2114 1818 3846 1821
rect 502 1803 505 1807
rect 501 1802 506 1803
rect 511 1802 512 1807
rect 1526 1803 1529 1807
rect 1525 1802 1530 1803
rect 1535 1802 1536 1807
rect 2550 1803 2553 1807
rect 2549 1802 2554 1803
rect 2559 1802 2560 1807
rect 3574 1803 3577 1807
rect 3573 1802 3578 1803
rect 3583 1802 3584 1807
rect 978 1788 2206 1791
rect 3370 1788 4141 1791
rect 4146 1788 4374 1791
rect 2466 1778 3326 1781
rect 882 1768 1742 1771
rect 1858 1768 3822 1771
rect 866 1758 1542 1761
rect 2970 1758 2973 1761
rect 3562 1758 3630 1761
rect 1162 1748 1382 1751
rect 2626 1748 2909 1751
rect 2994 1748 2998 1751
rect 3298 1748 3918 1751
rect 2250 1738 3166 1741
rect 1114 1728 1222 1731
rect 2290 1728 2494 1731
rect 2914 1728 2974 1731
rect 3010 1728 4422 1731
rect 2338 1718 2654 1721
rect 2930 1718 3238 1721
rect 1006 1703 1009 1707
rect 1005 1702 1010 1703
rect 1015 1702 1016 1707
rect 2030 1703 2033 1707
rect 2029 1702 2034 1703
rect 2039 1702 2040 1707
rect 3054 1703 3057 1707
rect 3053 1702 3058 1703
rect 3063 1702 3064 1707
rect 4086 1703 4089 1707
rect 4085 1702 4090 1703
rect 4095 1702 4096 1707
rect 554 1688 1222 1691
rect 2850 1688 3182 1691
rect 602 1678 1230 1681
rect 1314 1678 2342 1681
rect 2530 1678 2918 1681
rect 2922 1678 3206 1681
rect 3710 1681 3713 1688
rect 3986 1688 4358 1691
rect 3490 1678 3713 1681
rect 4378 1678 4590 1681
rect 2634 1668 2926 1671
rect 3106 1668 3361 1671
rect 3698 1668 3950 1671
rect 3358 1662 3361 1668
rect 3842 1658 3966 1661
rect 1762 1648 1942 1651
rect 3850 1648 4014 1651
rect 4410 1648 4518 1651
rect 3706 1638 4302 1641
rect 4466 1638 4526 1641
rect 2714 1628 3814 1631
rect 3818 1628 3982 1631
rect 2210 1618 4182 1621
rect 4238 1612 4241 1618
rect 2866 1608 2870 1611
rect 4162 1608 4230 1611
rect 502 1603 505 1607
rect 501 1602 506 1603
rect 511 1602 512 1607
rect 1526 1603 1529 1607
rect 1525 1602 1530 1603
rect 1535 1602 1536 1607
rect 2550 1603 2553 1607
rect 2549 1602 2554 1603
rect 2559 1602 2560 1607
rect 3574 1603 3577 1607
rect 3573 1602 3578 1603
rect 3583 1602 3584 1607
rect 3682 1598 4230 1601
rect 3498 1588 3526 1591
rect 3874 1588 4390 1591
rect 610 1578 782 1581
rect 3490 1578 4078 1581
rect 4162 1578 4398 1581
rect 2682 1568 2838 1571
rect 3922 1568 4174 1571
rect 4242 1568 4262 1571
rect 4206 1562 4209 1568
rect 1210 1558 1454 1561
rect 306 1548 510 1551
rect 2562 1548 2673 1551
rect 2882 1548 3182 1551
rect 3506 1548 3606 1551
rect 4178 1548 4230 1551
rect 2670 1542 2673 1548
rect 4402 1548 4406 1551
rect 1842 1538 2334 1541
rect 2866 1538 2902 1541
rect 3178 1538 3453 1541
rect 3522 1538 3526 1541
rect 2498 1528 2742 1531
rect 2746 1528 3990 1531
rect 4546 1528 4566 1531
rect 2706 1518 3406 1521
rect 4034 1518 4118 1521
rect 3946 1508 3990 1511
rect 1006 1503 1009 1507
rect 1005 1502 1010 1503
rect 1015 1502 1016 1507
rect 2030 1503 2033 1507
rect 2029 1502 2034 1503
rect 2039 1502 2040 1507
rect 3054 1503 3057 1507
rect 3053 1502 3058 1503
rect 3063 1502 3064 1507
rect 4086 1503 4089 1507
rect 4085 1502 4090 1503
rect 4095 1502 4096 1507
rect 4170 1498 4558 1501
rect 2862 1491 2865 1498
rect 2862 1488 3062 1491
rect 3218 1488 4390 1491
rect 1658 1478 1710 1481
rect 2170 1478 2750 1481
rect 2842 1478 2870 1481
rect 2282 1468 2462 1471
rect 3002 1468 3085 1471
rect 3090 1468 3094 1471
rect 3610 1468 3654 1471
rect 4018 1468 4238 1471
rect 1770 1458 2478 1461
rect 2694 1458 2702 1461
rect 2706 1458 3230 1461
rect 3386 1458 3742 1461
rect 4162 1458 4478 1461
rect 4514 1458 4558 1461
rect 2758 1448 3126 1451
rect 4234 1448 4310 1451
rect 2758 1441 2761 1448
rect 2482 1438 2761 1441
rect 3082 1438 3182 1441
rect 3186 1438 3782 1441
rect 3986 1438 4350 1441
rect 2538 1428 3278 1431
rect 1466 1418 1646 1421
rect 2194 1418 3078 1421
rect 3162 1418 4030 1421
rect 3122 1408 3134 1411
rect 502 1403 505 1407
rect 501 1402 506 1403
rect 511 1402 512 1407
rect 1526 1403 1529 1407
rect 1525 1402 1530 1403
rect 1535 1402 1536 1407
rect 2550 1403 2553 1407
rect 2549 1402 2554 1403
rect 2559 1402 2560 1407
rect 3574 1403 3577 1407
rect 3573 1402 3578 1403
rect 3583 1402 3584 1407
rect 3890 1398 3902 1401
rect 3970 1398 4486 1401
rect 4574 1392 4577 1398
rect 2730 1388 2733 1391
rect 3178 1388 4350 1391
rect 3274 1378 4270 1381
rect 1870 1371 1873 1378
rect 1870 1368 2646 1371
rect 2994 1368 4262 1371
rect 4266 1368 4381 1371
rect 4386 1368 4486 1371
rect 3458 1358 3886 1361
rect 4026 1358 4238 1361
rect 2358 1351 2361 1358
rect 4354 1358 4406 1361
rect 2358 1348 2462 1351
rect 3066 1348 3198 1351
rect 3842 1348 4494 1351
rect 2638 1342 2641 1348
rect 2938 1338 3190 1341
rect 3226 1338 3902 1341
rect 4030 1338 4206 1341
rect 4030 1332 4033 1338
rect 1594 1328 2254 1331
rect 2442 1328 2670 1331
rect 2922 1328 3214 1331
rect 3594 1328 3806 1331
rect 3810 1328 3958 1331
rect 1886 1318 1974 1321
rect 2666 1318 2846 1321
rect 2898 1318 3094 1321
rect 3098 1318 3286 1321
rect 3290 1318 3350 1321
rect 3354 1318 3478 1321
rect 3658 1318 3958 1321
rect 1886 1312 1889 1318
rect 2098 1308 2342 1311
rect 1006 1303 1009 1307
rect 1005 1302 1010 1303
rect 1015 1302 1016 1307
rect 2030 1303 2033 1307
rect 2029 1302 2034 1303
rect 2039 1302 2040 1307
rect 3054 1303 3057 1307
rect 3053 1302 3058 1303
rect 3063 1302 3064 1307
rect 4086 1303 4089 1307
rect 4085 1302 4090 1303
rect 4095 1302 4096 1307
rect 2738 1298 2974 1301
rect 3514 1298 4030 1301
rect 2978 1288 3142 1291
rect 3146 1288 3254 1291
rect 3906 1288 4462 1291
rect 2862 1282 2865 1287
rect 2546 1278 2750 1281
rect 2922 1278 3078 1281
rect 3106 1278 3478 1281
rect 3850 1278 4094 1281
rect 1186 1268 1542 1271
rect 2250 1268 2606 1271
rect 2722 1268 2926 1271
rect 3230 1268 3550 1271
rect 3626 1268 3750 1271
rect 1658 1258 1726 1261
rect 2898 1258 2910 1261
rect 3142 1261 3145 1268
rect 3066 1258 3145 1261
rect 3230 1262 3233 1268
rect 3826 1268 4590 1271
rect 3306 1258 4174 1261
rect 1658 1248 1910 1251
rect 2250 1248 2318 1251
rect 2898 1248 3542 1251
rect 3586 1248 3654 1251
rect 3658 1248 3846 1251
rect 3858 1248 4294 1251
rect 2802 1238 3206 1241
rect 3210 1238 3638 1241
rect 3698 1238 3886 1241
rect 1898 1228 3358 1231
rect 3434 1228 3678 1231
rect 3914 1228 4134 1231
rect 2658 1218 2910 1221
rect 2946 1218 2950 1221
rect 3090 1218 3214 1221
rect 3642 1218 4198 1221
rect 502 1203 505 1207
rect 501 1202 506 1203
rect 511 1202 512 1207
rect 1526 1203 1529 1207
rect 1525 1202 1530 1203
rect 1535 1202 1536 1207
rect 2550 1203 2553 1207
rect 2549 1202 2554 1203
rect 2559 1202 2560 1207
rect 3574 1203 3577 1207
rect 3573 1202 3578 1203
rect 3583 1202 3584 1207
rect 3106 1198 3254 1201
rect 3978 1198 4238 1201
rect 4386 1198 4414 1201
rect 3218 1188 3222 1191
rect 3562 1188 3734 1191
rect 4034 1188 4166 1191
rect 3042 1178 3486 1181
rect 3666 1178 3974 1181
rect 4106 1178 4438 1181
rect 402 1168 1174 1171
rect 2866 1168 3069 1171
rect 3146 1168 3326 1171
rect 3362 1168 3830 1171
rect 3938 1168 4134 1171
rect 4162 1168 4454 1171
rect 466 1158 486 1161
rect 2146 1158 2430 1161
rect 2434 1158 2782 1161
rect 2842 1158 2998 1161
rect 3110 1161 3113 1168
rect 3110 1158 3117 1161
rect 3122 1158 3286 1161
rect 3546 1158 4006 1161
rect 4010 1158 4254 1161
rect 1890 1148 2045 1151
rect 2394 1148 3150 1151
rect 3226 1148 3630 1151
rect 2410 1138 2654 1141
rect 2746 1138 3014 1141
rect 3170 1138 3417 1141
rect 3450 1138 3478 1141
rect 3594 1138 4030 1141
rect 4074 1138 4246 1141
rect 3414 1132 3417 1138
rect 1990 1128 1998 1131
rect 2002 1128 2054 1131
rect 2730 1128 2990 1131
rect 3042 1128 3270 1131
rect 3274 1128 3310 1131
rect 3442 1128 4230 1131
rect 2618 1118 2718 1121
rect 2962 1118 3454 1121
rect 3462 1118 3766 1121
rect 3778 1118 4158 1121
rect 2482 1108 2998 1111
rect 3462 1111 3465 1118
rect 3074 1108 3465 1111
rect 3514 1108 3670 1111
rect 3770 1108 4070 1111
rect 4186 1108 4189 1111
rect 1006 1103 1009 1107
rect 1005 1102 1010 1103
rect 1015 1102 1016 1107
rect 2030 1103 2033 1107
rect 2029 1102 2034 1103
rect 2039 1102 2040 1107
rect 3054 1103 3057 1107
rect 3053 1102 3058 1103
rect 3063 1102 3064 1107
rect 4086 1103 4089 1107
rect 4085 1102 4090 1103
rect 4095 1102 4096 1107
rect 2482 1098 2902 1101
rect 3258 1098 3526 1101
rect 3762 1098 3966 1101
rect 2002 1088 2110 1091
rect 2642 1088 2822 1091
rect 3194 1088 3774 1091
rect 3850 1088 3878 1091
rect 3986 1088 4214 1091
rect 4230 1088 4342 1091
rect 2494 1081 2497 1088
rect 2494 1078 2678 1081
rect 3002 1078 3182 1081
rect 3378 1078 3614 1081
rect 3634 1078 3766 1081
rect 2718 1071 2721 1078
rect 3842 1078 4038 1081
rect 4230 1081 4233 1088
rect 4130 1078 4233 1081
rect 4238 1072 4241 1078
rect 2718 1068 2830 1071
rect 3010 1068 3334 1071
rect 3362 1068 3566 1071
rect 3586 1068 3774 1071
rect 4434 1068 4462 1071
rect 1938 1058 2622 1061
rect 3034 1058 3158 1061
rect 3178 1058 4457 1061
rect 2706 1048 2750 1051
rect 2766 1051 2769 1058
rect 4046 1052 4049 1058
rect 4454 1052 4457 1058
rect 2766 1048 3862 1051
rect 3922 1048 4038 1051
rect 4098 1048 4406 1051
rect 3202 1038 3478 1041
rect 3506 1038 3582 1041
rect 3610 1038 4022 1041
rect 4042 1038 4262 1041
rect 2618 1028 3270 1031
rect 3514 1028 3558 1031
rect 3698 1028 4125 1031
rect 2010 1018 2569 1021
rect 2594 1018 3238 1021
rect 3338 1018 4006 1021
rect 1682 1008 1862 1011
rect 2566 1011 2569 1018
rect 2566 1008 3278 1011
rect 3418 1008 3534 1011
rect 3730 1008 4302 1011
rect 502 1003 505 1007
rect 501 1002 506 1003
rect 511 1002 512 1007
rect 1526 1003 1529 1007
rect 1525 1002 1530 1003
rect 1535 1002 1536 1007
rect 2550 1003 2553 1007
rect 2549 1002 2554 1003
rect 2559 1002 2560 1007
rect 3574 1003 3577 1007
rect 3573 1002 3578 1003
rect 3583 1002 3584 1007
rect 2954 998 2982 1001
rect 2986 998 3390 1001
rect 4194 998 4438 1001
rect 2054 991 2057 998
rect 2054 988 2862 991
rect 2890 988 3166 991
rect 3954 988 4382 991
rect 2042 978 2622 981
rect 3334 978 3438 981
rect 3562 978 3958 981
rect 3334 972 3337 978
rect 1890 968 2318 971
rect 2554 968 2790 971
rect 2938 968 3086 971
rect 3482 968 3806 971
rect 4050 968 4358 971
rect 1082 958 1454 961
rect 2026 958 2502 961
rect 2522 958 2646 961
rect 2786 958 2806 961
rect 2834 958 3741 961
rect 3794 958 3982 961
rect 3986 958 4062 961
rect 4066 958 4174 961
rect 4178 958 4358 961
rect 1074 948 1214 951
rect 1882 948 2190 951
rect 2370 948 2550 951
rect 2578 948 2966 951
rect 3082 948 3182 951
rect 3354 948 3886 951
rect 3898 948 4094 951
rect 4106 948 4270 951
rect 4542 942 4545 948
rect 1018 938 1486 941
rect 2394 938 2414 941
rect 2730 938 2854 941
rect 2914 938 3174 941
rect 3186 938 3222 941
rect 3226 938 3566 941
rect 3834 938 4190 941
rect 2682 928 2750 931
rect 2770 928 3238 931
rect 3710 931 3713 938
rect 3394 928 3713 931
rect 4178 928 4294 931
rect 4466 928 4558 931
rect 1726 918 1734 921
rect 1738 918 2109 921
rect 2802 918 2998 921
rect 3050 918 3102 921
rect 3242 918 3550 921
rect 3618 918 3758 921
rect 4074 918 4230 921
rect 4234 918 4398 921
rect 2234 908 2694 911
rect 3186 908 3518 911
rect 3738 908 3790 911
rect 4106 908 4526 911
rect 1006 903 1009 907
rect 1005 902 1010 903
rect 1015 902 1016 907
rect 2030 903 2033 907
rect 2029 902 2034 903
rect 2039 902 2040 907
rect 3054 903 3057 907
rect 3053 902 3058 903
rect 3063 902 3064 907
rect 4086 903 4089 907
rect 4085 902 4090 903
rect 4095 902 4096 907
rect 2130 898 2886 901
rect 2890 898 3041 901
rect 3106 898 3117 901
rect 2094 888 2829 891
rect 2094 881 2097 888
rect 3038 891 3041 898
rect 3242 898 3846 901
rect 3038 888 3213 891
rect 3218 888 3222 891
rect 3282 888 3673 891
rect 3682 888 3894 891
rect 1626 878 2097 881
rect 2114 878 2129 881
rect 2218 878 2382 881
rect 2490 878 2726 881
rect 2858 878 3030 881
rect 3042 878 3181 881
rect 2126 872 2129 878
rect 3450 878 3590 881
rect 3670 881 3673 888
rect 3670 878 4214 881
rect 946 868 1118 871
rect 2226 868 2462 871
rect 2466 868 2494 871
rect 2746 868 2878 871
rect 2970 868 3198 871
rect 3394 868 3526 871
rect 3530 868 3726 871
rect 3802 868 3862 871
rect 4438 871 4441 878
rect 3930 868 4441 871
rect 2018 858 2174 861
rect 2234 858 2342 861
rect 2514 858 2862 861
rect 2962 858 3110 861
rect 3482 858 3934 861
rect 4162 858 4270 861
rect 4294 858 4406 861
rect 4294 852 4297 858
rect 1194 848 1406 851
rect 1962 848 2126 851
rect 2386 848 2726 851
rect 3074 848 3849 851
rect 4010 848 4278 851
rect 3846 842 3849 848
rect 2346 838 2470 841
rect 2514 838 2694 841
rect 2730 838 3574 841
rect 4138 838 4486 841
rect 2322 828 2590 831
rect 2610 828 3502 831
rect 3818 828 4166 831
rect 2602 818 2862 821
rect 3506 818 4038 821
rect 3522 808 3526 811
rect 502 803 505 807
rect 501 802 506 803
rect 511 802 512 807
rect 1526 803 1529 807
rect 1525 802 1530 803
rect 1535 802 1536 807
rect 2550 803 2553 807
rect 2549 802 2554 803
rect 2559 802 2560 807
rect 3574 803 3577 807
rect 3573 802 3578 803
rect 3583 802 3584 807
rect 4206 802 4209 807
rect 2530 798 2534 801
rect 2854 798 3326 801
rect 3338 798 3550 801
rect 1722 788 2334 791
rect 2854 791 2857 798
rect 2514 788 2857 791
rect 2866 788 3302 791
rect 3458 788 3830 791
rect 4042 788 4518 791
rect 1570 778 2845 781
rect 3162 778 3438 781
rect 3442 778 3654 781
rect 1882 768 2605 771
rect 2994 768 3758 771
rect 3826 768 3910 771
rect 3954 768 4542 771
rect 2594 758 2934 761
rect 3026 758 3390 761
rect 1878 751 1881 758
rect 1778 748 1881 751
rect 1914 748 2262 751
rect 2802 748 2974 751
rect 3218 748 3774 751
rect 4010 748 4030 751
rect 4210 748 4262 751
rect 1850 738 2934 741
rect 2938 738 3142 741
rect 3426 738 3566 741
rect 2410 728 2934 731
rect 2946 728 2950 731
rect 3138 728 3366 731
rect 3482 728 3622 731
rect 4066 728 4278 731
rect 4374 731 4377 738
rect 4282 728 4377 731
rect 2618 718 3382 721
rect 3386 718 3438 721
rect 4066 718 4173 721
rect 4378 718 4397 721
rect 2274 708 2966 711
rect 3202 708 3838 711
rect 1006 703 1009 707
rect 1005 702 1010 703
rect 1015 702 1016 707
rect 2030 703 2033 707
rect 2029 702 2034 703
rect 2039 702 2040 707
rect 3054 703 3057 707
rect 3053 702 3058 703
rect 3063 702 3064 707
rect 4086 703 4089 707
rect 4085 702 4090 703
rect 4095 702 4096 707
rect 2666 698 2822 701
rect 1954 688 2041 691
rect 2538 688 2694 691
rect 3170 688 3358 691
rect 2038 682 2041 688
rect 3662 682 3665 687
rect 2146 678 2918 681
rect 4226 678 4238 681
rect 4142 672 4145 677
rect 1746 668 2190 671
rect 2274 668 2733 671
rect 2882 668 3654 671
rect 314 658 558 661
rect 2494 652 2497 658
rect 2738 658 2806 661
rect 4066 658 4566 661
rect 250 648 430 651
rect 2642 648 2718 651
rect 3074 648 3262 651
rect 2706 638 4134 641
rect 1874 628 3622 631
rect 4122 628 4429 631
rect 1634 618 2877 621
rect 2978 618 3686 621
rect 4010 618 4222 621
rect 3786 608 4158 611
rect 502 603 505 607
rect 501 602 506 603
rect 511 602 512 607
rect 1526 603 1529 607
rect 1525 602 1530 603
rect 1535 602 1536 607
rect 2550 603 2553 607
rect 2549 602 2554 603
rect 2559 602 2560 607
rect 3574 603 3577 607
rect 3573 602 3578 603
rect 3583 602 3584 607
rect 2126 592 2129 598
rect 2834 588 4110 591
rect 2058 578 2158 581
rect 2162 578 2326 581
rect 2330 578 4014 581
rect 4082 578 4350 581
rect 3706 568 4126 571
rect 2014 561 2017 568
rect 2014 558 2366 561
rect 2594 558 2734 561
rect 2906 558 4230 561
rect 4234 558 4238 561
rect 2962 548 3118 551
rect 3314 548 3870 551
rect 4130 548 4310 551
rect 1730 538 2046 541
rect 3106 538 3398 541
rect 4194 538 4205 541
rect 4562 538 4574 541
rect 1634 528 3494 531
rect 3826 528 4270 531
rect 2402 518 2926 521
rect 4114 518 4589 521
rect 2226 508 2862 511
rect 3490 508 4022 511
rect 1006 503 1009 507
rect 1005 502 1010 503
rect 1015 502 1016 507
rect 2030 503 2033 507
rect 2029 502 2034 503
rect 2039 502 2040 507
rect 3054 503 3057 507
rect 3053 502 3058 503
rect 3063 502 3064 507
rect 4086 503 4089 507
rect 4085 502 4090 503
rect 4095 502 4096 507
rect 3074 498 3966 501
rect 2178 488 3038 491
rect 4146 488 4422 491
rect 3742 482 3745 488
rect 1978 478 1990 481
rect 1994 478 3069 481
rect 4574 472 4577 478
rect 210 468 382 471
rect 2226 468 2462 471
rect 2762 468 3974 471
rect 4242 468 4422 471
rect 290 458 1198 461
rect 2594 458 2718 461
rect 2722 458 2806 461
rect 2866 458 3910 461
rect 3914 458 4038 461
rect 2634 448 2702 451
rect 3298 448 3302 451
rect 3906 448 4454 451
rect 2794 438 3822 441
rect 1690 428 3694 431
rect 3938 428 4518 431
rect 1610 418 3526 421
rect 3962 418 4302 421
rect 502 403 505 407
rect 501 402 506 403
rect 511 402 512 407
rect 1526 403 1529 407
rect 1525 402 1530 403
rect 1535 402 1536 407
rect 2550 403 2553 407
rect 2549 402 2554 403
rect 2559 402 2560 407
rect 3574 403 3577 407
rect 3573 402 3578 403
rect 3583 402 3584 407
rect 3082 398 3085 401
rect 4186 398 4189 401
rect 3458 388 4174 391
rect 2450 378 2702 381
rect 2714 378 3950 381
rect 2130 368 2390 371
rect 2394 368 3806 371
rect 3930 368 4502 371
rect 1714 358 1742 361
rect 1842 358 2822 361
rect 3018 358 3702 361
rect 1846 348 1918 351
rect 2634 348 2678 351
rect 3718 351 3721 358
rect 3718 348 3814 351
rect 3822 348 4014 351
rect 1846 342 1849 348
rect 2482 338 2681 341
rect 2818 338 3294 341
rect 3402 338 3422 341
rect 3822 341 3825 348
rect 3658 338 3825 341
rect 4054 341 4057 348
rect 4002 338 4057 341
rect 4074 338 4545 341
rect 2678 332 2681 338
rect 4542 332 4545 338
rect 3034 328 3673 331
rect 3978 328 4214 331
rect 3670 322 3673 328
rect 1986 318 2158 321
rect 2810 318 3478 321
rect 3486 318 3614 321
rect 3706 318 3990 321
rect 4018 318 4525 321
rect 2154 308 2294 311
rect 3486 311 3489 318
rect 3314 308 3489 311
rect 3562 308 4073 311
rect 1006 303 1009 307
rect 1005 302 1010 303
rect 1015 302 1016 307
rect 2030 303 2033 307
rect 2029 302 2034 303
rect 2039 302 2040 307
rect 3054 303 3057 307
rect 3053 302 3058 303
rect 3063 302 3064 307
rect 3294 302 3297 307
rect 4070 302 4073 308
rect 4086 303 4089 307
rect 4085 302 4090 303
rect 4095 302 4096 307
rect 3546 298 3710 301
rect 3794 298 3965 301
rect 2018 288 2766 291
rect 2770 288 4318 291
rect 1834 278 2686 281
rect 2842 278 3309 281
rect 3394 278 3550 281
rect 3738 278 3821 281
rect 3842 278 3917 281
rect 4130 278 4406 281
rect 4482 278 4486 281
rect 186 268 614 271
rect 3234 268 3662 271
rect 3826 268 3837 271
rect 3922 268 3981 271
rect 242 258 1598 261
rect 2162 258 2542 261
rect 2546 258 3174 261
rect 3202 258 3502 261
rect 3778 258 3982 261
rect 4202 258 4278 261
rect 370 248 606 251
rect 2306 248 2502 251
rect 2930 248 3206 251
rect 3370 248 3814 251
rect 3906 248 4094 251
rect 2234 238 2518 241
rect 2522 238 2974 241
rect 3770 238 4294 241
rect 2418 228 2758 231
rect 3178 228 4054 231
rect 4074 228 4214 231
rect 2730 218 3318 221
rect 3658 218 3942 221
rect 3962 218 4222 221
rect 2866 208 3486 211
rect 3762 208 3853 211
rect 3954 208 3966 211
rect 502 203 505 207
rect 501 202 506 203
rect 511 202 512 207
rect 1526 203 1529 207
rect 1525 202 1530 203
rect 1535 202 1536 207
rect 2550 203 2553 207
rect 2549 202 2554 203
rect 2559 202 2560 207
rect 3574 203 3577 207
rect 3573 202 3578 203
rect 3583 202 3584 207
rect 2778 198 3230 201
rect 3858 198 3869 201
rect 3882 198 4126 201
rect 4138 198 4254 201
rect 3218 188 3654 191
rect 3666 188 4318 191
rect 1874 178 2790 181
rect 3282 178 3462 181
rect 3466 178 3518 181
rect 3562 178 4150 181
rect 4186 178 4310 181
rect 2354 168 2958 171
rect 2978 168 3118 171
rect 3466 168 4158 171
rect 4194 168 4221 171
rect 938 158 1190 161
rect 1890 158 2926 161
rect 2930 158 3645 161
rect 3650 158 3686 161
rect 3822 158 4238 161
rect 266 148 1686 151
rect 2154 148 2382 151
rect 2762 148 2806 151
rect 2978 148 3446 151
rect 3822 151 3825 158
rect 4542 152 4545 158
rect 3586 148 3825 151
rect 3834 148 3950 151
rect 3962 148 4061 151
rect 4090 148 4206 151
rect 4226 148 4349 151
rect 2202 138 2422 141
rect 2514 138 2950 141
rect 3042 138 3254 141
rect 3566 138 3574 141
rect 3578 138 4350 141
rect 2370 128 2590 131
rect 2634 128 3030 131
rect 3274 128 3974 131
rect 3998 128 4062 131
rect 4074 128 4253 131
rect 690 118 1510 121
rect 1994 118 2374 121
rect 2618 118 3110 121
rect 3170 118 3574 121
rect 3602 118 3910 121
rect 3998 121 4001 128
rect 4266 128 4381 131
rect 3938 118 4001 121
rect 4010 118 4342 121
rect 2786 108 3038 111
rect 3378 108 3606 111
rect 3770 108 3854 111
rect 3890 108 3950 111
rect 4034 108 4045 111
rect 4258 108 4350 111
rect 1006 103 1009 107
rect 1005 102 1010 103
rect 1015 102 1016 107
rect 2030 103 2033 107
rect 2029 102 2034 103
rect 2039 102 2040 107
rect 3054 103 3057 107
rect 3053 102 3058 103
rect 3063 102 3064 107
rect 4086 103 4089 107
rect 4085 102 4090 103
rect 4095 102 4096 107
rect 2426 98 2646 101
rect 2818 98 2845 101
rect 3258 98 3782 101
rect 3842 98 4038 101
rect 2362 88 2365 91
rect 2994 88 3150 91
rect 3282 88 3614 91
rect 3714 88 3766 91
rect 3810 88 3814 91
rect 3858 88 4438 91
rect 2238 78 2398 81
rect 2574 78 2998 81
rect 3026 78 3166 81
rect 3322 78 3593 81
rect 3602 78 3837 81
rect 2238 72 2241 78
rect 2574 72 2577 78
rect 2066 68 2238 71
rect 2282 68 2574 71
rect 2850 68 3118 71
rect 3122 68 3246 71
rect 3434 68 3518 71
rect 3590 71 3593 78
rect 3850 78 3853 81
rect 3862 78 3870 81
rect 3890 78 4230 81
rect 4258 78 4470 81
rect 3862 71 3865 78
rect 3590 68 3865 71
rect 3874 68 3901 71
rect 3930 68 3934 71
rect 3978 68 4046 71
rect 4130 68 4134 71
rect 4158 68 4510 71
rect 922 58 1502 61
rect 1818 58 2526 61
rect 3058 58 3078 61
rect 3114 58 3294 61
rect 3298 58 3702 61
rect 4158 61 4161 68
rect 3794 58 4161 61
rect 4178 58 4205 61
rect 2526 51 2529 58
rect 4210 58 4270 61
rect 2526 48 3486 51
rect 3802 48 4157 51
rect 3018 38 3302 41
rect 3858 38 4269 41
rect 3330 28 3942 31
rect 3962 28 4110 31
rect 3906 18 4557 21
rect 3886 12 3889 18
rect 3970 8 4029 11
rect 4082 8 4534 11
rect 502 3 505 7
rect 501 2 506 3
rect 511 2 512 7
rect 1526 3 1529 7
rect 1525 2 1530 3
rect 1535 2 1536 7
rect 2550 3 2553 7
rect 2549 2 2554 3
rect 2559 2 2560 7
rect 3574 3 3577 7
rect 3573 2 3578 3
rect 3583 2 3584 7
<< m6contact >>
rect 496 4403 498 4407
rect 498 4403 501 4407
rect 506 4403 509 4407
rect 509 4403 511 4407
rect 496 4402 501 4403
rect 506 4402 511 4403
rect 1520 4403 1522 4407
rect 1522 4403 1525 4407
rect 1530 4403 1533 4407
rect 1533 4403 1535 4407
rect 1520 4402 1525 4403
rect 1530 4402 1535 4403
rect 2544 4403 2546 4407
rect 2546 4403 2549 4407
rect 2554 4403 2557 4407
rect 2557 4403 2559 4407
rect 2544 4402 2549 4403
rect 2554 4402 2559 4403
rect 3568 4403 3570 4407
rect 3570 4403 3573 4407
rect 3578 4403 3581 4407
rect 3581 4403 3583 4407
rect 3568 4402 3573 4403
rect 3578 4402 3583 4403
rect 4445 4347 4450 4352
rect 4477 4347 4482 4352
rect 4381 4327 4386 4332
rect 1000 4303 1002 4307
rect 1002 4303 1005 4307
rect 1010 4303 1013 4307
rect 1013 4303 1015 4307
rect 1000 4302 1005 4303
rect 1010 4302 1015 4303
rect 2024 4303 2026 4307
rect 2026 4303 2029 4307
rect 2034 4303 2037 4307
rect 2037 4303 2039 4307
rect 2024 4302 2029 4303
rect 2034 4302 2039 4303
rect 3048 4303 3050 4307
rect 3050 4303 3053 4307
rect 3058 4303 3061 4307
rect 3061 4303 3063 4307
rect 3048 4302 3053 4303
rect 3058 4302 3063 4303
rect 4080 4303 4082 4307
rect 4082 4303 4085 4307
rect 4090 4303 4093 4307
rect 4093 4303 4095 4307
rect 4080 4302 4085 4303
rect 4090 4302 4095 4303
rect 4573 4307 4578 4312
rect 4461 4287 4466 4292
rect 496 4203 498 4207
rect 498 4203 501 4207
rect 506 4203 509 4207
rect 509 4203 511 4207
rect 496 4202 501 4203
rect 506 4202 511 4203
rect 1520 4203 1522 4207
rect 1522 4203 1525 4207
rect 1530 4203 1533 4207
rect 1533 4203 1535 4207
rect 1520 4202 1525 4203
rect 1530 4202 1535 4203
rect 2544 4203 2546 4207
rect 2546 4203 2549 4207
rect 2554 4203 2557 4207
rect 2557 4203 2559 4207
rect 2544 4202 2549 4203
rect 2554 4202 2559 4203
rect 3568 4203 3570 4207
rect 3570 4203 3573 4207
rect 3578 4203 3581 4207
rect 3581 4203 3583 4207
rect 3568 4202 3573 4203
rect 3578 4202 3583 4203
rect 4541 4107 4546 4112
rect 1000 4103 1002 4107
rect 1002 4103 1005 4107
rect 1010 4103 1013 4107
rect 1013 4103 1015 4107
rect 1000 4102 1005 4103
rect 1010 4102 1015 4103
rect 2024 4103 2026 4107
rect 2026 4103 2029 4107
rect 2034 4103 2037 4107
rect 2037 4103 2039 4107
rect 2024 4102 2029 4103
rect 2034 4102 2039 4103
rect 3048 4103 3050 4107
rect 3050 4103 3053 4107
rect 3058 4103 3061 4107
rect 3061 4103 3063 4107
rect 3048 4102 3053 4103
rect 3058 4102 3063 4103
rect 4080 4103 4082 4107
rect 4082 4103 4085 4107
rect 4090 4103 4093 4107
rect 4093 4103 4095 4107
rect 4080 4102 4085 4103
rect 4090 4102 4095 4103
rect 4557 4087 4562 4092
rect 496 4003 498 4007
rect 498 4003 501 4007
rect 506 4003 509 4007
rect 509 4003 511 4007
rect 496 4002 501 4003
rect 506 4002 511 4003
rect 1520 4003 1522 4007
rect 1522 4003 1525 4007
rect 1530 4003 1533 4007
rect 1533 4003 1535 4007
rect 1520 4002 1525 4003
rect 1530 4002 1535 4003
rect 2544 4003 2546 4007
rect 2546 4003 2549 4007
rect 2554 4003 2557 4007
rect 2557 4003 2559 4007
rect 2544 4002 2549 4003
rect 2554 4002 2559 4003
rect 3568 4003 3570 4007
rect 3570 4003 3573 4007
rect 3578 4003 3581 4007
rect 3581 4003 3583 4007
rect 3568 4002 3573 4003
rect 3578 4002 3583 4003
rect 1000 3903 1002 3907
rect 1002 3903 1005 3907
rect 1010 3903 1013 3907
rect 1013 3903 1015 3907
rect 1000 3902 1005 3903
rect 1010 3902 1015 3903
rect 2024 3903 2026 3907
rect 2026 3903 2029 3907
rect 2034 3903 2037 3907
rect 2037 3903 2039 3907
rect 2024 3902 2029 3903
rect 2034 3902 2039 3903
rect 3048 3903 3050 3907
rect 3050 3903 3053 3907
rect 3058 3903 3061 3907
rect 3061 3903 3063 3907
rect 3048 3902 3053 3903
rect 3058 3902 3063 3903
rect 4080 3903 4082 3907
rect 4082 3903 4085 3907
rect 4090 3903 4093 3907
rect 4093 3903 4095 3907
rect 4080 3902 4085 3903
rect 4090 3902 4095 3903
rect 4509 3817 4514 3822
rect 496 3803 498 3807
rect 498 3803 501 3807
rect 506 3803 509 3807
rect 509 3803 511 3807
rect 496 3802 501 3803
rect 506 3802 511 3803
rect 1520 3803 1522 3807
rect 1522 3803 1525 3807
rect 1530 3803 1533 3807
rect 1533 3803 1535 3807
rect 1520 3802 1525 3803
rect 1530 3802 1535 3803
rect 2544 3803 2546 3807
rect 2546 3803 2549 3807
rect 2554 3803 2557 3807
rect 2557 3803 2559 3807
rect 2544 3802 2549 3803
rect 2554 3802 2559 3803
rect 3568 3803 3570 3807
rect 3570 3803 3573 3807
rect 3578 3803 3581 3807
rect 3581 3803 3583 3807
rect 3568 3802 3573 3803
rect 3578 3802 3583 3803
rect 2333 3707 2338 3712
rect 1000 3703 1002 3707
rect 1002 3703 1005 3707
rect 1010 3703 1013 3707
rect 1013 3703 1015 3707
rect 1000 3702 1005 3703
rect 1010 3702 1015 3703
rect 2024 3703 2026 3707
rect 2026 3703 2029 3707
rect 2034 3703 2037 3707
rect 2037 3703 2039 3707
rect 2024 3702 2029 3703
rect 2034 3702 2039 3703
rect 3048 3703 3050 3707
rect 3050 3703 3053 3707
rect 3058 3703 3061 3707
rect 3061 3703 3063 3707
rect 3048 3702 3053 3703
rect 3058 3702 3063 3703
rect 4080 3703 4082 3707
rect 4082 3703 4085 3707
rect 4090 3703 4093 3707
rect 4093 3703 4095 3707
rect 4080 3702 4085 3703
rect 4090 3702 4095 3703
rect 496 3603 498 3607
rect 498 3603 501 3607
rect 506 3603 509 3607
rect 509 3603 511 3607
rect 496 3602 501 3603
rect 506 3602 511 3603
rect 1520 3603 1522 3607
rect 1522 3603 1525 3607
rect 1530 3603 1533 3607
rect 1533 3603 1535 3607
rect 1520 3602 1525 3603
rect 1530 3602 1535 3603
rect 2544 3603 2546 3607
rect 2546 3603 2549 3607
rect 2554 3603 2557 3607
rect 2557 3603 2559 3607
rect 2544 3602 2549 3603
rect 2554 3602 2559 3603
rect 3568 3603 3570 3607
rect 3570 3603 3573 3607
rect 3578 3603 3581 3607
rect 3581 3603 3583 3607
rect 3568 3602 3573 3603
rect 3578 3602 3583 3603
rect 2653 3507 2658 3512
rect 1000 3503 1002 3507
rect 1002 3503 1005 3507
rect 1010 3503 1013 3507
rect 1013 3503 1015 3507
rect 1000 3502 1005 3503
rect 1010 3502 1015 3503
rect 2024 3503 2026 3507
rect 2026 3503 2029 3507
rect 2034 3503 2037 3507
rect 2037 3503 2039 3507
rect 2024 3502 2029 3503
rect 2034 3502 2039 3503
rect 3048 3503 3050 3507
rect 3050 3503 3053 3507
rect 3058 3503 3061 3507
rect 3061 3503 3063 3507
rect 3048 3502 3053 3503
rect 3058 3502 3063 3503
rect 4080 3503 4082 3507
rect 4082 3503 4085 3507
rect 4090 3503 4093 3507
rect 4093 3503 4095 3507
rect 4080 3502 4085 3503
rect 4090 3502 4095 3503
rect 4429 3467 4434 3472
rect 2829 3437 2834 3442
rect 496 3403 498 3407
rect 498 3403 501 3407
rect 506 3403 509 3407
rect 509 3403 511 3407
rect 496 3402 501 3403
rect 506 3402 511 3403
rect 1520 3403 1522 3407
rect 1522 3403 1525 3407
rect 1530 3403 1533 3407
rect 1533 3403 1535 3407
rect 1520 3402 1525 3403
rect 1530 3402 1535 3403
rect 2544 3403 2546 3407
rect 2546 3403 2549 3407
rect 2554 3403 2557 3407
rect 2557 3403 2559 3407
rect 2544 3402 2549 3403
rect 2554 3402 2559 3403
rect 3568 3403 3570 3407
rect 3570 3403 3573 3407
rect 3578 3403 3581 3407
rect 3581 3403 3583 3407
rect 3568 3402 3573 3403
rect 3578 3402 3583 3403
rect 2829 3387 2834 3392
rect 2333 3337 2338 3342
rect 2525 3327 2530 3332
rect 1000 3303 1002 3307
rect 1002 3303 1005 3307
rect 1010 3303 1013 3307
rect 1013 3303 1015 3307
rect 1000 3302 1005 3303
rect 1010 3302 1015 3303
rect 2024 3303 2026 3307
rect 2026 3303 2029 3307
rect 2034 3303 2037 3307
rect 2037 3303 2039 3307
rect 2024 3302 2029 3303
rect 2034 3302 2039 3303
rect 3048 3303 3050 3307
rect 3050 3303 3053 3307
rect 3058 3303 3061 3307
rect 3061 3303 3063 3307
rect 3048 3302 3053 3303
rect 3058 3302 3063 3303
rect 4080 3303 4082 3307
rect 4082 3303 4085 3307
rect 4090 3303 4093 3307
rect 4093 3303 4095 3307
rect 4080 3302 4085 3303
rect 4090 3302 4095 3303
rect 4589 3237 4594 3242
rect 496 3203 498 3207
rect 498 3203 501 3207
rect 506 3203 509 3207
rect 509 3203 511 3207
rect 496 3202 501 3203
rect 506 3202 511 3203
rect 1520 3203 1522 3207
rect 1522 3203 1525 3207
rect 1530 3203 1533 3207
rect 1533 3203 1535 3207
rect 1520 3202 1525 3203
rect 1530 3202 1535 3203
rect 2544 3203 2546 3207
rect 2546 3203 2549 3207
rect 2554 3203 2557 3207
rect 2557 3203 2559 3207
rect 2544 3202 2549 3203
rect 2554 3202 2559 3203
rect 3568 3203 3570 3207
rect 3570 3203 3573 3207
rect 3578 3203 3581 3207
rect 3581 3203 3583 3207
rect 3568 3202 3573 3203
rect 3578 3202 3583 3203
rect 2653 3157 2658 3162
rect 1000 3103 1002 3107
rect 1002 3103 1005 3107
rect 1010 3103 1013 3107
rect 1013 3103 1015 3107
rect 1000 3102 1005 3103
rect 1010 3102 1015 3103
rect 2024 3103 2026 3107
rect 2026 3103 2029 3107
rect 2034 3103 2037 3107
rect 2037 3103 2039 3107
rect 2024 3102 2029 3103
rect 2034 3102 2039 3103
rect 3048 3103 3050 3107
rect 3050 3103 3053 3107
rect 3058 3103 3061 3107
rect 3061 3103 3063 3107
rect 3048 3102 3053 3103
rect 3058 3102 3063 3103
rect 4080 3103 4082 3107
rect 4082 3103 4085 3107
rect 4090 3103 4093 3107
rect 4093 3103 4095 3107
rect 4080 3102 4085 3103
rect 4090 3102 4095 3103
rect 2045 3097 2050 3102
rect 496 3003 498 3007
rect 498 3003 501 3007
rect 506 3003 509 3007
rect 509 3003 511 3007
rect 496 3002 501 3003
rect 506 3002 511 3003
rect 1520 3003 1522 3007
rect 1522 3003 1525 3007
rect 1530 3003 1533 3007
rect 1533 3003 1535 3007
rect 1520 3002 1525 3003
rect 1530 3002 1535 3003
rect 2544 3003 2546 3007
rect 2546 3003 2549 3007
rect 2554 3003 2557 3007
rect 2557 3003 2559 3007
rect 2544 3002 2549 3003
rect 2554 3002 2559 3003
rect 3568 3003 3570 3007
rect 3570 3003 3573 3007
rect 3578 3003 3581 3007
rect 3581 3003 3583 3007
rect 3568 3002 3573 3003
rect 3578 3002 3583 3003
rect 1000 2903 1002 2907
rect 1002 2903 1005 2907
rect 1010 2903 1013 2907
rect 1013 2903 1015 2907
rect 1000 2902 1005 2903
rect 1010 2902 1015 2903
rect 2024 2903 2026 2907
rect 2026 2903 2029 2907
rect 2034 2903 2037 2907
rect 2037 2903 2039 2907
rect 2024 2902 2029 2903
rect 2034 2902 2039 2903
rect 3048 2903 3050 2907
rect 3050 2903 3053 2907
rect 3058 2903 3061 2907
rect 3061 2903 3063 2907
rect 3048 2902 3053 2903
rect 3058 2902 3063 2903
rect 4080 2903 4082 2907
rect 4082 2903 4085 2907
rect 4090 2903 4093 2907
rect 4093 2903 4095 2907
rect 4080 2902 4085 2903
rect 4090 2902 4095 2903
rect 3949 2877 3954 2882
rect 4477 2807 4482 2812
rect 496 2803 498 2807
rect 498 2803 501 2807
rect 506 2803 509 2807
rect 509 2803 511 2807
rect 496 2802 501 2803
rect 506 2802 511 2803
rect 1520 2803 1522 2807
rect 1522 2803 1525 2807
rect 1530 2803 1533 2807
rect 1533 2803 1535 2807
rect 1520 2802 1525 2803
rect 1530 2802 1535 2803
rect 2544 2803 2546 2807
rect 2546 2803 2549 2807
rect 2554 2803 2557 2807
rect 2557 2803 2559 2807
rect 2544 2802 2549 2803
rect 2554 2802 2559 2803
rect 3568 2803 3570 2807
rect 3570 2803 3573 2807
rect 3578 2803 3581 2807
rect 3581 2803 3583 2807
rect 3568 2802 3573 2803
rect 3578 2802 3583 2803
rect 4477 2707 4482 2712
rect 1000 2703 1002 2707
rect 1002 2703 1005 2707
rect 1010 2703 1013 2707
rect 1013 2703 1015 2707
rect 1000 2702 1005 2703
rect 1010 2702 1015 2703
rect 2024 2703 2026 2707
rect 2026 2703 2029 2707
rect 2034 2703 2037 2707
rect 2037 2703 2039 2707
rect 2024 2702 2029 2703
rect 2034 2702 2039 2703
rect 3048 2703 3050 2707
rect 3050 2703 3053 2707
rect 3058 2703 3061 2707
rect 3061 2703 3063 2707
rect 3048 2702 3053 2703
rect 3058 2702 3063 2703
rect 4080 2703 4082 2707
rect 4082 2703 4085 2707
rect 4090 2703 4093 2707
rect 4093 2703 4095 2707
rect 4080 2702 4085 2703
rect 4090 2702 4095 2703
rect 496 2603 498 2607
rect 498 2603 501 2607
rect 506 2603 509 2607
rect 509 2603 511 2607
rect 496 2602 501 2603
rect 506 2602 511 2603
rect 1520 2603 1522 2607
rect 1522 2603 1525 2607
rect 1530 2603 1533 2607
rect 1533 2603 1535 2607
rect 1520 2602 1525 2603
rect 1530 2602 1535 2603
rect 2544 2603 2546 2607
rect 2546 2603 2549 2607
rect 2554 2603 2557 2607
rect 2557 2603 2559 2607
rect 2544 2602 2549 2603
rect 2554 2602 2559 2603
rect 3568 2603 3570 2607
rect 3570 2603 3573 2607
rect 3578 2603 3581 2607
rect 3581 2603 3583 2607
rect 3568 2602 3573 2603
rect 3578 2602 3583 2603
rect 3805 2567 3810 2572
rect 2125 2547 2130 2552
rect 3853 2547 3858 2552
rect 3741 2527 3746 2532
rect 3661 2517 3666 2522
rect 1000 2503 1002 2507
rect 1002 2503 1005 2507
rect 1010 2503 1013 2507
rect 1013 2503 1015 2507
rect 1000 2502 1005 2503
rect 1010 2502 1015 2503
rect 2024 2503 2026 2507
rect 2026 2503 2029 2507
rect 2034 2503 2037 2507
rect 2037 2503 2039 2507
rect 2024 2502 2029 2503
rect 2034 2502 2039 2503
rect 3048 2503 3050 2507
rect 3050 2503 3053 2507
rect 3058 2503 3061 2507
rect 3061 2503 3063 2507
rect 3048 2502 3053 2503
rect 3058 2502 3063 2503
rect 4080 2503 4082 2507
rect 4082 2503 4085 2507
rect 4090 2503 4093 2507
rect 4093 2503 4095 2507
rect 4080 2502 4085 2503
rect 4090 2502 4095 2503
rect 496 2403 498 2407
rect 498 2403 501 2407
rect 506 2403 509 2407
rect 509 2403 511 2407
rect 496 2402 501 2403
rect 506 2402 511 2403
rect 1520 2403 1522 2407
rect 1522 2403 1525 2407
rect 1530 2403 1533 2407
rect 1533 2403 1535 2407
rect 1520 2402 1525 2403
rect 1530 2402 1535 2403
rect 2544 2403 2546 2407
rect 2546 2403 2549 2407
rect 2554 2403 2557 2407
rect 2557 2403 2559 2407
rect 2544 2402 2549 2403
rect 2554 2402 2559 2403
rect 3568 2403 3570 2407
rect 3570 2403 3573 2407
rect 3578 2403 3581 2407
rect 3581 2403 3583 2407
rect 3568 2402 3573 2403
rect 3578 2402 3583 2403
rect 2365 2367 2370 2372
rect 3725 2357 3730 2362
rect 3645 2337 3650 2342
rect 4269 2337 4274 2342
rect 4445 2337 4450 2342
rect 1000 2303 1002 2307
rect 1002 2303 1005 2307
rect 1010 2303 1013 2307
rect 1013 2303 1015 2307
rect 1000 2302 1005 2303
rect 1010 2302 1015 2303
rect 2024 2303 2026 2307
rect 2026 2303 2029 2307
rect 2034 2303 2037 2307
rect 2037 2303 2039 2307
rect 2024 2302 2029 2303
rect 2034 2302 2039 2303
rect 3048 2303 3050 2307
rect 3050 2303 3053 2307
rect 3058 2303 3061 2307
rect 3061 2303 3063 2307
rect 3048 2302 3053 2303
rect 3058 2302 3063 2303
rect 4080 2303 4082 2307
rect 4082 2303 4085 2307
rect 4090 2303 4093 2307
rect 4093 2303 4095 2307
rect 4080 2302 4085 2303
rect 4090 2302 4095 2303
rect 2845 2287 2850 2292
rect 4525 2257 4530 2262
rect 4173 2227 4178 2232
rect 496 2203 498 2207
rect 498 2203 501 2207
rect 506 2203 509 2207
rect 509 2203 511 2207
rect 496 2202 501 2203
rect 506 2202 511 2203
rect 1520 2203 1522 2207
rect 1522 2203 1525 2207
rect 1530 2203 1533 2207
rect 1533 2203 1535 2207
rect 1520 2202 1525 2203
rect 1530 2202 1535 2203
rect 2544 2203 2546 2207
rect 2546 2203 2549 2207
rect 2554 2203 2557 2207
rect 2557 2203 2559 2207
rect 2544 2202 2549 2203
rect 2554 2202 2559 2203
rect 3568 2203 3570 2207
rect 3570 2203 3573 2207
rect 3578 2203 3581 2207
rect 3581 2203 3583 2207
rect 3568 2202 3573 2203
rect 3578 2202 3583 2203
rect 1000 2103 1002 2107
rect 1002 2103 1005 2107
rect 1010 2103 1013 2107
rect 1013 2103 1015 2107
rect 1000 2102 1005 2103
rect 1010 2102 1015 2103
rect 2024 2103 2026 2107
rect 2026 2103 2029 2107
rect 2034 2103 2037 2107
rect 2037 2103 2039 2107
rect 2024 2102 2029 2103
rect 2034 2102 2039 2103
rect 3048 2103 3050 2107
rect 3050 2103 3053 2107
rect 3058 2103 3061 2107
rect 3061 2103 3063 2107
rect 3048 2102 3053 2103
rect 3058 2102 3063 2103
rect 4080 2103 4082 2107
rect 4082 2103 4085 2107
rect 4090 2103 4093 2107
rect 4093 2103 4095 2107
rect 4080 2102 4085 2103
rect 4090 2102 4095 2103
rect 496 2003 498 2007
rect 498 2003 501 2007
rect 506 2003 509 2007
rect 509 2003 511 2007
rect 496 2002 501 2003
rect 506 2002 511 2003
rect 1520 2003 1522 2007
rect 1522 2003 1525 2007
rect 1530 2003 1533 2007
rect 1533 2003 1535 2007
rect 1520 2002 1525 2003
rect 1530 2002 1535 2003
rect 2544 2003 2546 2007
rect 2546 2003 2549 2007
rect 2554 2003 2557 2007
rect 2557 2003 2559 2007
rect 2544 2002 2549 2003
rect 2554 2002 2559 2003
rect 3568 2003 3570 2007
rect 3570 2003 3573 2007
rect 3578 2003 3581 2007
rect 3581 2003 3583 2007
rect 3568 2002 3573 2003
rect 3578 2002 3583 2003
rect 1000 1903 1002 1907
rect 1002 1903 1005 1907
rect 1010 1903 1013 1907
rect 1013 1903 1015 1907
rect 1000 1902 1005 1903
rect 1010 1902 1015 1903
rect 2024 1903 2026 1907
rect 2026 1903 2029 1907
rect 2034 1903 2037 1907
rect 2037 1903 2039 1907
rect 2024 1902 2029 1903
rect 2034 1902 2039 1903
rect 3048 1903 3050 1907
rect 3050 1903 3053 1907
rect 3058 1903 3061 1907
rect 3061 1903 3063 1907
rect 3048 1902 3053 1903
rect 3058 1902 3063 1903
rect 4080 1903 4082 1907
rect 4082 1903 4085 1907
rect 4090 1903 4093 1907
rect 4093 1903 4095 1907
rect 4080 1902 4085 1903
rect 4090 1902 4095 1903
rect 3709 1887 3714 1892
rect 496 1803 498 1807
rect 498 1803 501 1807
rect 506 1803 509 1807
rect 509 1803 511 1807
rect 496 1802 501 1803
rect 506 1802 511 1803
rect 1520 1803 1522 1807
rect 1522 1803 1525 1807
rect 1530 1803 1533 1807
rect 1533 1803 1535 1807
rect 1520 1802 1525 1803
rect 1530 1802 1535 1803
rect 2544 1803 2546 1807
rect 2546 1803 2549 1807
rect 2554 1803 2557 1807
rect 2557 1803 2559 1807
rect 2544 1802 2549 1803
rect 2554 1802 2559 1803
rect 3568 1803 3570 1807
rect 3570 1803 3573 1807
rect 3578 1803 3581 1807
rect 3581 1803 3583 1807
rect 3568 1802 3573 1803
rect 3578 1802 3583 1803
rect 4141 1787 4146 1792
rect 2973 1757 2978 1762
rect 2909 1747 2914 1752
rect 2989 1747 2994 1752
rect 2909 1727 2914 1732
rect 1000 1703 1002 1707
rect 1002 1703 1005 1707
rect 1010 1703 1013 1707
rect 1013 1703 1015 1707
rect 1000 1702 1005 1703
rect 1010 1702 1015 1703
rect 2024 1703 2026 1707
rect 2026 1703 2029 1707
rect 2034 1703 2037 1707
rect 2037 1703 2039 1707
rect 2024 1702 2029 1703
rect 2034 1702 2039 1703
rect 3048 1703 3050 1707
rect 3050 1703 3053 1707
rect 3058 1703 3061 1707
rect 3061 1703 3063 1707
rect 3048 1702 3053 1703
rect 3058 1702 3063 1703
rect 4080 1703 4082 1707
rect 4082 1703 4085 1707
rect 4090 1703 4093 1707
rect 4093 1703 4095 1707
rect 4080 1702 4085 1703
rect 4090 1702 4095 1703
rect 3981 1687 3986 1692
rect 4461 1637 4466 1642
rect 2861 1607 2866 1612
rect 4157 1607 4162 1612
rect 4237 1607 4242 1612
rect 496 1603 498 1607
rect 498 1603 501 1607
rect 506 1603 509 1607
rect 509 1603 511 1607
rect 496 1602 501 1603
rect 506 1602 511 1603
rect 1520 1603 1522 1607
rect 1522 1603 1525 1607
rect 1530 1603 1533 1607
rect 1533 1603 1535 1607
rect 1520 1602 1525 1603
rect 1530 1602 1535 1603
rect 2544 1603 2546 1607
rect 2546 1603 2549 1607
rect 2554 1603 2557 1607
rect 2557 1603 2559 1607
rect 2544 1602 2549 1603
rect 2554 1602 2559 1603
rect 3568 1603 3570 1607
rect 3570 1603 3573 1607
rect 3578 1603 3581 1607
rect 3581 1603 3583 1607
rect 3568 1602 3573 1603
rect 3578 1602 3583 1603
rect 3869 1587 3874 1592
rect 3917 1567 3922 1572
rect 4205 1557 4210 1562
rect 4397 1547 4402 1552
rect 3453 1537 3458 1542
rect 3517 1537 3522 1542
rect 2493 1527 2498 1532
rect 4541 1527 4546 1532
rect 4029 1517 4034 1522
rect 1000 1503 1002 1507
rect 1002 1503 1005 1507
rect 1010 1503 1013 1507
rect 1013 1503 1015 1507
rect 1000 1502 1005 1503
rect 1010 1502 1015 1503
rect 2024 1503 2026 1507
rect 2026 1503 2029 1507
rect 2034 1503 2037 1507
rect 2037 1503 2039 1507
rect 2024 1502 2029 1503
rect 2034 1502 2039 1503
rect 3048 1503 3050 1507
rect 3050 1503 3053 1507
rect 3058 1503 3061 1507
rect 3061 1503 3063 1507
rect 3048 1502 3053 1503
rect 3058 1502 3063 1503
rect 4080 1503 4082 1507
rect 4082 1503 4085 1507
rect 4090 1503 4093 1507
rect 4093 1503 4095 1507
rect 4080 1502 4085 1503
rect 4090 1502 4095 1503
rect 3085 1467 3090 1472
rect 4509 1457 4514 1462
rect 496 1403 498 1407
rect 498 1403 501 1407
rect 506 1403 509 1407
rect 509 1403 511 1407
rect 496 1402 501 1403
rect 506 1402 511 1403
rect 1520 1403 1522 1407
rect 1522 1403 1525 1407
rect 1530 1403 1533 1407
rect 1533 1403 1535 1407
rect 1520 1402 1525 1403
rect 1530 1402 1535 1403
rect 2544 1403 2546 1407
rect 2546 1403 2549 1407
rect 2554 1403 2557 1407
rect 2557 1403 2559 1407
rect 2544 1402 2549 1403
rect 2554 1402 2559 1403
rect 3568 1403 3570 1407
rect 3570 1403 3573 1407
rect 3578 1403 3581 1407
rect 3581 1403 3583 1407
rect 3568 1402 3573 1403
rect 3578 1402 3583 1403
rect 3885 1397 3890 1402
rect 3965 1397 3970 1402
rect 2733 1387 2738 1392
rect 4573 1387 4578 1392
rect 4381 1367 4386 1372
rect 4349 1357 4354 1362
rect 2637 1337 2642 1342
rect 1000 1303 1002 1307
rect 1002 1303 1005 1307
rect 1010 1303 1013 1307
rect 1013 1303 1015 1307
rect 1000 1302 1005 1303
rect 1010 1302 1015 1303
rect 2024 1303 2026 1307
rect 2026 1303 2029 1307
rect 2034 1303 2037 1307
rect 2037 1303 2039 1307
rect 2024 1302 2029 1303
rect 2034 1302 2039 1303
rect 3048 1303 3050 1307
rect 3050 1303 3053 1307
rect 3058 1303 3061 1307
rect 3061 1303 3063 1307
rect 3048 1302 3053 1303
rect 3058 1302 3063 1303
rect 4080 1303 4082 1307
rect 4082 1303 4085 1307
rect 4090 1303 4093 1307
rect 4093 1303 4095 1307
rect 4080 1302 4085 1303
rect 4090 1302 4095 1303
rect 2861 1287 2866 1292
rect 3901 1287 3906 1292
rect 3821 1267 3826 1272
rect 2941 1217 2946 1222
rect 496 1203 498 1207
rect 498 1203 501 1207
rect 506 1203 509 1207
rect 509 1203 511 1207
rect 496 1202 501 1203
rect 506 1202 511 1203
rect 1520 1203 1522 1207
rect 1522 1203 1525 1207
rect 1530 1203 1533 1207
rect 1533 1203 1535 1207
rect 1520 1202 1525 1203
rect 1530 1202 1535 1203
rect 2544 1203 2546 1207
rect 2546 1203 2549 1207
rect 2554 1203 2557 1207
rect 2557 1203 2559 1207
rect 2544 1202 2549 1203
rect 2554 1202 2559 1203
rect 3568 1203 3570 1207
rect 3570 1203 3573 1207
rect 3578 1203 3581 1207
rect 3581 1203 3583 1207
rect 3568 1202 3573 1203
rect 3578 1202 3583 1203
rect 4381 1197 4386 1202
rect 3213 1187 3218 1192
rect 3069 1167 3074 1172
rect 3117 1157 3122 1162
rect 2045 1147 2050 1152
rect 3069 1107 3074 1112
rect 4189 1107 4194 1112
rect 1000 1103 1002 1107
rect 1002 1103 1005 1107
rect 1010 1103 1013 1107
rect 1013 1103 1015 1107
rect 1000 1102 1005 1103
rect 1010 1102 1015 1103
rect 2024 1103 2026 1107
rect 2026 1103 2029 1107
rect 2034 1103 2037 1107
rect 2037 1103 2039 1107
rect 2024 1102 2029 1103
rect 2034 1102 2039 1103
rect 3048 1103 3050 1107
rect 3050 1103 3053 1107
rect 3058 1103 3061 1107
rect 3061 1103 3063 1107
rect 3048 1102 3053 1103
rect 3058 1102 3063 1103
rect 4080 1103 4082 1107
rect 4082 1103 4085 1107
rect 4090 1103 4093 1107
rect 4093 1103 4095 1107
rect 4080 1102 4085 1103
rect 4090 1102 4095 1103
rect 3837 1077 3842 1082
rect 4125 1077 4130 1082
rect 4237 1067 4242 1072
rect 4125 1027 4130 1032
rect 3725 1007 3730 1012
rect 496 1003 498 1007
rect 498 1003 501 1007
rect 506 1003 509 1007
rect 509 1003 511 1007
rect 496 1002 501 1003
rect 506 1002 511 1003
rect 1520 1003 1522 1007
rect 1522 1003 1525 1007
rect 1530 1003 1533 1007
rect 1533 1003 1535 1007
rect 1520 1002 1525 1003
rect 1530 1002 1535 1003
rect 2544 1003 2546 1007
rect 2546 1003 2549 1007
rect 2554 1003 2557 1007
rect 2557 1003 2559 1007
rect 2544 1002 2549 1003
rect 2554 1002 2559 1003
rect 3568 1003 3570 1007
rect 3570 1003 3573 1007
rect 3578 1003 3581 1007
rect 3581 1003 3583 1007
rect 3568 1002 3573 1003
rect 3578 1002 3583 1003
rect 3949 987 3954 992
rect 4045 967 4050 972
rect 2829 957 2834 962
rect 3741 957 3746 962
rect 3181 937 3186 942
rect 4541 937 4546 942
rect 2109 917 2114 922
rect 1000 903 1002 907
rect 1002 903 1005 907
rect 1010 903 1013 907
rect 1013 903 1015 907
rect 1000 902 1005 903
rect 1010 902 1015 903
rect 2024 903 2026 907
rect 2026 903 2029 907
rect 2034 903 2037 907
rect 2037 903 2039 907
rect 2024 902 2029 903
rect 2034 902 2039 903
rect 3048 903 3050 907
rect 3050 903 3053 907
rect 3058 903 3061 907
rect 3061 903 3063 907
rect 3048 902 3053 903
rect 3058 902 3063 903
rect 4080 903 4082 907
rect 4082 903 4085 907
rect 4090 903 4093 907
rect 4093 903 4095 907
rect 4080 902 4085 903
rect 4090 902 4095 903
rect 2829 887 2834 892
rect 3117 897 3122 902
rect 3213 887 3218 892
rect 2109 877 2114 882
rect 3181 877 3186 882
rect 2605 827 2610 832
rect 3517 807 3522 812
rect 4205 807 4210 812
rect 496 803 498 807
rect 498 803 501 807
rect 506 803 509 807
rect 509 803 511 807
rect 496 802 501 803
rect 506 802 511 803
rect 1520 803 1522 807
rect 1522 803 1525 807
rect 1530 803 1533 807
rect 1533 803 1535 807
rect 1520 802 1525 803
rect 1530 802 1535 803
rect 2544 803 2546 807
rect 2546 803 2549 807
rect 2554 803 2557 807
rect 2557 803 2559 807
rect 2544 802 2549 803
rect 2554 802 2559 803
rect 3568 803 3570 807
rect 3570 803 3573 807
rect 3578 803 3581 807
rect 3581 803 3583 807
rect 3568 802 3573 803
rect 3578 802 3583 803
rect 2525 797 2530 802
rect 3453 787 3458 792
rect 2845 777 2850 782
rect 2605 767 2610 772
rect 2989 767 2994 772
rect 3949 767 3954 772
rect 2941 727 2946 732
rect 4173 717 4178 722
rect 4397 717 4402 722
rect 1000 703 1002 707
rect 1002 703 1005 707
rect 1010 703 1013 707
rect 1013 703 1015 707
rect 1000 702 1005 703
rect 1010 702 1015 703
rect 2024 703 2026 707
rect 2026 703 2029 707
rect 2034 703 2037 707
rect 2037 703 2039 707
rect 2024 702 2029 703
rect 2034 702 2039 703
rect 3048 703 3050 707
rect 3050 703 3053 707
rect 3058 703 3061 707
rect 3061 703 3063 707
rect 3048 702 3053 703
rect 3058 702 3063 703
rect 4080 703 4082 707
rect 4082 703 4085 707
rect 4090 703 4093 707
rect 4093 703 4095 707
rect 4080 702 4085 703
rect 4090 702 4095 703
rect 3661 687 3666 692
rect 4141 677 4146 682
rect 4221 677 4226 682
rect 2733 667 2738 672
rect 2877 667 2882 672
rect 2733 657 2738 662
rect 4061 657 4066 662
rect 2493 647 2498 652
rect 2637 647 2642 652
rect 4429 627 4434 632
rect 2877 617 2882 622
rect 2973 617 2978 622
rect 496 603 498 607
rect 498 603 501 607
rect 506 603 509 607
rect 509 603 511 607
rect 496 602 501 603
rect 506 602 511 603
rect 1520 603 1522 607
rect 1522 603 1525 607
rect 1530 603 1533 607
rect 1533 603 1535 607
rect 1520 602 1525 603
rect 1530 602 1535 603
rect 2544 603 2546 607
rect 2546 603 2549 607
rect 2554 603 2557 607
rect 2557 603 2559 607
rect 2544 602 2549 603
rect 2554 602 2559 603
rect 3568 603 3570 607
rect 3570 603 3573 607
rect 3578 603 3581 607
rect 3581 603 3583 607
rect 3568 602 3573 603
rect 3578 602 3583 603
rect 2125 587 2130 592
rect 4205 537 4210 542
rect 4557 537 4562 542
rect 4589 517 4594 522
rect 1000 503 1002 507
rect 1002 503 1005 507
rect 1010 503 1013 507
rect 1013 503 1015 507
rect 1000 502 1005 503
rect 1010 502 1015 503
rect 2024 503 2026 507
rect 2026 503 2029 507
rect 2034 503 2037 507
rect 2037 503 2039 507
rect 2024 502 2029 503
rect 2034 502 2039 503
rect 3048 503 3050 507
rect 3050 503 3053 507
rect 3058 503 3061 507
rect 3061 503 3063 507
rect 3048 502 3053 503
rect 3058 502 3063 503
rect 4080 503 4082 507
rect 4082 503 4085 507
rect 4090 503 4093 507
rect 4093 503 4095 507
rect 4080 502 4085 503
rect 4090 502 4095 503
rect 3069 497 3074 502
rect 3069 477 3074 482
rect 3741 477 3746 482
rect 4573 467 4578 472
rect 3293 447 3298 452
rect 3933 427 3938 432
rect 496 403 498 407
rect 498 403 501 407
rect 506 403 509 407
rect 509 403 511 407
rect 496 402 501 403
rect 506 402 511 403
rect 1520 403 1522 407
rect 1522 403 1525 407
rect 1530 403 1533 407
rect 1533 403 1535 407
rect 1520 402 1525 403
rect 1530 402 1535 403
rect 2544 403 2546 407
rect 2546 403 2549 407
rect 2554 403 2557 407
rect 2557 403 2559 407
rect 2544 402 2549 403
rect 2554 402 2559 403
rect 3568 403 3570 407
rect 3570 403 3573 407
rect 3578 403 3581 407
rect 3581 403 3583 407
rect 3568 402 3573 403
rect 3578 402 3583 403
rect 3085 397 3090 402
rect 4189 397 4194 402
rect 3293 307 3298 312
rect 3309 307 3314 312
rect 4525 317 4530 322
rect 1000 303 1002 307
rect 1002 303 1005 307
rect 1010 303 1013 307
rect 1013 303 1015 307
rect 1000 302 1005 303
rect 1010 302 1015 303
rect 2024 303 2026 307
rect 2026 303 2029 307
rect 2034 303 2037 307
rect 2037 303 2039 307
rect 2024 302 2029 303
rect 2034 302 2039 303
rect 3048 303 3050 307
rect 3050 303 3053 307
rect 3058 303 3061 307
rect 3061 303 3063 307
rect 3048 302 3053 303
rect 3058 302 3063 303
rect 4080 303 4082 307
rect 4082 303 4085 307
rect 4090 303 4093 307
rect 4093 303 4095 307
rect 4080 302 4085 303
rect 4090 302 4095 303
rect 3965 297 3970 302
rect 3309 277 3314 282
rect 3821 277 3826 282
rect 3917 277 3922 282
rect 4125 277 4130 282
rect 4477 277 4482 282
rect 3837 267 3842 272
rect 3981 267 3986 272
rect 3853 207 3858 212
rect 3949 207 3954 212
rect 496 203 498 207
rect 498 203 501 207
rect 506 203 509 207
rect 509 203 511 207
rect 496 202 501 203
rect 506 202 511 203
rect 1520 203 1522 207
rect 1522 203 1525 207
rect 1530 203 1533 207
rect 1533 203 1535 207
rect 1520 202 1525 203
rect 1530 202 1535 203
rect 2544 203 2546 207
rect 2546 203 2549 207
rect 2554 203 2557 207
rect 2557 203 2559 207
rect 2544 202 2549 203
rect 2554 202 2559 203
rect 3568 203 3570 207
rect 3570 203 3573 207
rect 3578 203 3581 207
rect 3581 203 3583 207
rect 3568 202 3573 203
rect 3578 202 3583 203
rect 3853 197 3858 202
rect 3869 197 3874 202
rect 4221 167 4226 172
rect 3645 157 3650 162
rect 4061 147 4066 152
rect 4349 147 4354 152
rect 4541 147 4546 152
rect 4253 127 4258 132
rect 4381 127 4386 132
rect 4045 107 4050 112
rect 4253 107 4258 112
rect 1000 103 1002 107
rect 1002 103 1005 107
rect 1010 103 1013 107
rect 1013 103 1015 107
rect 1000 102 1005 103
rect 1010 102 1015 103
rect 2024 103 2026 107
rect 2026 103 2029 107
rect 2034 103 2037 107
rect 2037 103 2039 107
rect 2024 102 2029 103
rect 2034 102 2039 103
rect 3048 103 3050 107
rect 3050 103 3053 107
rect 3058 103 3061 107
rect 3061 103 3063 107
rect 3048 102 3053 103
rect 3058 102 3063 103
rect 4080 103 4082 107
rect 4082 103 4085 107
rect 4090 103 4093 107
rect 4093 103 4095 107
rect 4080 102 4085 103
rect 4090 102 4095 103
rect 2845 97 2850 102
rect 3837 97 3842 102
rect 2365 87 2370 92
rect 3709 87 3714 92
rect 3805 87 3810 92
rect 3837 77 3842 82
rect 3853 77 3858 82
rect 3901 67 3906 72
rect 3925 67 3930 72
rect 4125 67 4130 72
rect 4205 57 4210 62
rect 4157 47 4162 52
rect 4269 37 4274 42
rect 4557 17 4562 22
rect 3885 7 3890 12
rect 4029 7 4034 12
rect 496 3 498 7
rect 498 3 501 7
rect 506 3 509 7
rect 509 3 511 7
rect 496 2 501 3
rect 506 2 511 3
rect 1520 3 1522 7
rect 1522 3 1525 7
rect 1530 3 1533 7
rect 1533 3 1535 7
rect 1520 2 1525 3
rect 1530 2 1535 3
rect 2544 3 2546 7
rect 2546 3 2549 7
rect 2554 3 2557 7
rect 2557 3 2559 7
rect 2544 2 2549 3
rect 2554 2 2559 3
rect 3568 3 3570 7
rect 3570 3 3573 7
rect 3578 3 3581 7
rect 3581 3 3583 7
rect 3568 2 3573 3
rect 3578 2 3583 3
<< metal6 >>
rect 496 4407 512 4430
rect 501 4402 506 4407
rect 511 4402 512 4407
rect 496 4207 512 4402
rect 501 4202 506 4207
rect 511 4202 512 4207
rect 496 4007 512 4202
rect 501 4002 506 4007
rect 511 4002 512 4007
rect 496 3807 512 4002
rect 501 3802 506 3807
rect 511 3802 512 3807
rect 496 3607 512 3802
rect 501 3602 506 3607
rect 511 3602 512 3607
rect 496 3407 512 3602
rect 501 3402 506 3407
rect 511 3402 512 3407
rect 496 3207 512 3402
rect 501 3202 506 3207
rect 511 3202 512 3207
rect 496 3007 512 3202
rect 501 3002 506 3007
rect 511 3002 512 3007
rect 496 2807 512 3002
rect 501 2802 506 2807
rect 511 2802 512 2807
rect 496 2607 512 2802
rect 501 2602 506 2607
rect 511 2602 512 2607
rect 496 2407 512 2602
rect 501 2402 506 2407
rect 511 2402 512 2407
rect 496 2207 512 2402
rect 501 2202 506 2207
rect 511 2202 512 2207
rect 496 2007 512 2202
rect 501 2002 506 2007
rect 511 2002 512 2007
rect 496 1807 512 2002
rect 501 1802 506 1807
rect 511 1802 512 1807
rect 496 1607 512 1802
rect 501 1602 506 1607
rect 511 1602 512 1607
rect 496 1407 512 1602
rect 501 1402 506 1407
rect 511 1402 512 1407
rect 496 1207 512 1402
rect 501 1202 506 1207
rect 511 1202 512 1207
rect 496 1007 512 1202
rect 501 1002 506 1007
rect 511 1002 512 1007
rect 496 807 512 1002
rect 501 802 506 807
rect 511 802 512 807
rect 496 607 512 802
rect 501 602 506 607
rect 511 602 512 607
rect 496 407 512 602
rect 501 402 506 407
rect 511 402 512 407
rect 496 207 512 402
rect 501 202 506 207
rect 511 202 512 207
rect 496 7 512 202
rect 501 2 506 7
rect 511 2 512 7
rect 496 -30 512 2
rect 1000 4307 1016 4430
rect 1005 4302 1010 4307
rect 1015 4302 1016 4307
rect 1000 4107 1016 4302
rect 1005 4102 1010 4107
rect 1015 4102 1016 4107
rect 1000 3907 1016 4102
rect 1005 3902 1010 3907
rect 1015 3902 1016 3907
rect 1000 3707 1016 3902
rect 1005 3702 1010 3707
rect 1015 3702 1016 3707
rect 1000 3507 1016 3702
rect 1005 3502 1010 3507
rect 1015 3502 1016 3507
rect 1000 3307 1016 3502
rect 1005 3302 1010 3307
rect 1015 3302 1016 3307
rect 1000 3107 1016 3302
rect 1005 3102 1010 3107
rect 1015 3102 1016 3107
rect 1000 2907 1016 3102
rect 1005 2902 1010 2907
rect 1015 2902 1016 2907
rect 1000 2707 1016 2902
rect 1005 2702 1010 2707
rect 1015 2702 1016 2707
rect 1000 2507 1016 2702
rect 1005 2502 1010 2507
rect 1015 2502 1016 2507
rect 1000 2307 1016 2502
rect 1005 2302 1010 2307
rect 1015 2302 1016 2307
rect 1000 2107 1016 2302
rect 1005 2102 1010 2107
rect 1015 2102 1016 2107
rect 1000 1907 1016 2102
rect 1005 1902 1010 1907
rect 1015 1902 1016 1907
rect 1000 1707 1016 1902
rect 1005 1702 1010 1707
rect 1015 1702 1016 1707
rect 1000 1507 1016 1702
rect 1005 1502 1010 1507
rect 1015 1502 1016 1507
rect 1000 1307 1016 1502
rect 1005 1302 1010 1307
rect 1015 1302 1016 1307
rect 1000 1107 1016 1302
rect 1005 1102 1010 1107
rect 1015 1102 1016 1107
rect 1000 907 1016 1102
rect 1005 902 1010 907
rect 1015 902 1016 907
rect 1000 707 1016 902
rect 1005 702 1010 707
rect 1015 702 1016 707
rect 1000 507 1016 702
rect 1005 502 1010 507
rect 1015 502 1016 507
rect 1000 307 1016 502
rect 1005 302 1010 307
rect 1015 302 1016 307
rect 1000 107 1016 302
rect 1005 102 1010 107
rect 1015 102 1016 107
rect 1000 -30 1016 102
rect 1520 4407 1536 4430
rect 1525 4402 1530 4407
rect 1535 4402 1536 4407
rect 1520 4207 1536 4402
rect 1525 4202 1530 4207
rect 1535 4202 1536 4207
rect 1520 4007 1536 4202
rect 1525 4002 1530 4007
rect 1535 4002 1536 4007
rect 1520 3807 1536 4002
rect 1525 3802 1530 3807
rect 1535 3802 1536 3807
rect 1520 3607 1536 3802
rect 1525 3602 1530 3607
rect 1535 3602 1536 3607
rect 1520 3407 1536 3602
rect 1525 3402 1530 3407
rect 1535 3402 1536 3407
rect 1520 3207 1536 3402
rect 1525 3202 1530 3207
rect 1535 3202 1536 3207
rect 1520 3007 1536 3202
rect 1525 3002 1530 3007
rect 1535 3002 1536 3007
rect 1520 2807 1536 3002
rect 1525 2802 1530 2807
rect 1535 2802 1536 2807
rect 1520 2607 1536 2802
rect 1525 2602 1530 2607
rect 1535 2602 1536 2607
rect 1520 2407 1536 2602
rect 1525 2402 1530 2407
rect 1535 2402 1536 2407
rect 1520 2207 1536 2402
rect 1525 2202 1530 2207
rect 1535 2202 1536 2207
rect 1520 2007 1536 2202
rect 1525 2002 1530 2007
rect 1535 2002 1536 2007
rect 1520 1807 1536 2002
rect 1525 1802 1530 1807
rect 1535 1802 1536 1807
rect 1520 1607 1536 1802
rect 1525 1602 1530 1607
rect 1535 1602 1536 1607
rect 1520 1407 1536 1602
rect 1525 1402 1530 1407
rect 1535 1402 1536 1407
rect 1520 1207 1536 1402
rect 1525 1202 1530 1207
rect 1535 1202 1536 1207
rect 1520 1007 1536 1202
rect 1525 1002 1530 1007
rect 1535 1002 1536 1007
rect 1520 807 1536 1002
rect 1525 802 1530 807
rect 1535 802 1536 807
rect 1520 607 1536 802
rect 1525 602 1530 607
rect 1535 602 1536 607
rect 1520 407 1536 602
rect 1525 402 1530 407
rect 1535 402 1536 407
rect 1520 207 1536 402
rect 1525 202 1530 207
rect 1535 202 1536 207
rect 1520 7 1536 202
rect 1525 2 1530 7
rect 1535 2 1536 7
rect 1520 -30 1536 2
rect 2024 4307 2040 4430
rect 2029 4302 2034 4307
rect 2039 4302 2040 4307
rect 2024 4107 2040 4302
rect 2029 4102 2034 4107
rect 2039 4102 2040 4107
rect 2024 3907 2040 4102
rect 2029 3902 2034 3907
rect 2039 3902 2040 3907
rect 2024 3707 2040 3902
rect 2544 4407 2560 4430
rect 2549 4402 2554 4407
rect 2559 4402 2560 4407
rect 2544 4207 2560 4402
rect 2549 4202 2554 4207
rect 2559 4202 2560 4207
rect 2544 4007 2560 4202
rect 2549 4002 2554 4007
rect 2559 4002 2560 4007
rect 2544 3807 2560 4002
rect 2549 3802 2554 3807
rect 2559 3802 2560 3807
rect 2029 3702 2034 3707
rect 2039 3702 2040 3707
rect 2024 3507 2040 3702
rect 2029 3502 2034 3507
rect 2039 3502 2040 3507
rect 2024 3307 2040 3502
rect 2333 3342 2338 3707
rect 2544 3607 2560 3802
rect 2549 3602 2554 3607
rect 2559 3602 2560 3607
rect 2544 3407 2560 3602
rect 3048 4307 3064 4430
rect 3053 4302 3058 4307
rect 3063 4302 3064 4307
rect 3048 4107 3064 4302
rect 3053 4102 3058 4107
rect 3063 4102 3064 4107
rect 3048 3907 3064 4102
rect 3053 3902 3058 3907
rect 3063 3902 3064 3907
rect 3048 3707 3064 3902
rect 3053 3702 3058 3707
rect 3063 3702 3064 3707
rect 2549 3402 2554 3407
rect 2559 3402 2560 3407
rect 2029 3302 2034 3307
rect 2039 3302 2040 3307
rect 2024 3107 2040 3302
rect 2029 3102 2034 3107
rect 2039 3102 2040 3107
rect 2024 2907 2040 3102
rect 2029 2902 2034 2907
rect 2039 2902 2040 2907
rect 2024 2707 2040 2902
rect 2029 2702 2034 2707
rect 2039 2702 2040 2707
rect 2024 2507 2040 2702
rect 2029 2502 2034 2507
rect 2039 2502 2040 2507
rect 2024 2307 2040 2502
rect 2029 2302 2034 2307
rect 2039 2302 2040 2307
rect 2024 2107 2040 2302
rect 2029 2102 2034 2107
rect 2039 2102 2040 2107
rect 2024 1907 2040 2102
rect 2029 1902 2034 1907
rect 2039 1902 2040 1907
rect 2024 1707 2040 1902
rect 2029 1702 2034 1707
rect 2039 1702 2040 1707
rect 2024 1507 2040 1702
rect 2029 1502 2034 1507
rect 2039 1502 2040 1507
rect 2024 1307 2040 1502
rect 2029 1302 2034 1307
rect 2039 1302 2040 1307
rect 2024 1107 2040 1302
rect 2045 1152 2050 3097
rect 2029 1102 2034 1107
rect 2039 1102 2040 1107
rect 2024 907 2040 1102
rect 2029 902 2034 907
rect 2039 902 2040 907
rect 2024 707 2040 902
rect 2109 882 2114 917
rect 2029 702 2034 707
rect 2039 702 2040 707
rect 2024 507 2040 702
rect 2125 592 2130 2547
rect 2029 502 2034 507
rect 2039 502 2040 507
rect 2024 307 2040 502
rect 2029 302 2034 307
rect 2039 302 2040 307
rect 2024 107 2040 302
rect 2029 102 2034 107
rect 2039 102 2040 107
rect 2024 -30 2040 102
rect 2365 92 2370 2367
rect 2493 652 2498 1527
rect 2525 802 2530 3327
rect 2544 3207 2560 3402
rect 2549 3202 2554 3207
rect 2559 3202 2560 3207
rect 2544 3007 2560 3202
rect 2653 3162 2658 3507
rect 3048 3507 3064 3702
rect 3053 3502 3058 3507
rect 3063 3502 3064 3507
rect 2829 3392 2834 3437
rect 3048 3307 3064 3502
rect 3053 3302 3058 3307
rect 3063 3302 3064 3307
rect 2549 3002 2554 3007
rect 2559 3002 2560 3007
rect 2544 2807 2560 3002
rect 2549 2802 2554 2807
rect 2559 2802 2560 2807
rect 2544 2607 2560 2802
rect 2549 2602 2554 2607
rect 2559 2602 2560 2607
rect 2544 2407 2560 2602
rect 2549 2402 2554 2407
rect 2559 2402 2560 2407
rect 2544 2207 2560 2402
rect 3048 3107 3064 3302
rect 3053 3102 3058 3107
rect 3063 3102 3064 3107
rect 3048 2907 3064 3102
rect 3053 2902 3058 2907
rect 3063 2902 3064 2907
rect 3048 2707 3064 2902
rect 3053 2702 3058 2707
rect 3063 2702 3064 2707
rect 3048 2507 3064 2702
rect 3053 2502 3058 2507
rect 3063 2502 3064 2507
rect 3048 2307 3064 2502
rect 3053 2302 3058 2307
rect 3063 2302 3064 2307
rect 2549 2202 2554 2207
rect 2559 2202 2560 2207
rect 2544 2007 2560 2202
rect 2549 2002 2554 2007
rect 2559 2002 2560 2007
rect 2544 1807 2560 2002
rect 2549 1802 2554 1807
rect 2559 1802 2560 1807
rect 2544 1607 2560 1802
rect 2549 1602 2554 1607
rect 2559 1602 2560 1607
rect 2544 1407 2560 1602
rect 2549 1402 2554 1407
rect 2559 1402 2560 1407
rect 2544 1207 2560 1402
rect 2549 1202 2554 1207
rect 2559 1202 2560 1207
rect 2544 1007 2560 1202
rect 2549 1002 2554 1007
rect 2559 1002 2560 1007
rect 2544 807 2560 1002
rect 2549 802 2554 807
rect 2559 802 2560 807
rect 2544 607 2560 802
rect 2605 772 2610 827
rect 2637 652 2642 1337
rect 2733 672 2738 1387
rect 2829 892 2834 957
rect 2733 662 2738 667
rect 2845 782 2850 2287
rect 3048 2107 3064 2302
rect 3053 2102 3058 2107
rect 3063 2102 3064 2107
rect 3048 1907 3064 2102
rect 3053 1902 3058 1907
rect 3063 1902 3064 1907
rect 2909 1732 2914 1747
rect 2861 1292 2866 1607
rect 2549 602 2554 607
rect 2559 602 2560 607
rect 2544 407 2560 602
rect 2549 402 2554 407
rect 2559 402 2560 407
rect 2544 207 2560 402
rect 2549 202 2554 207
rect 2559 202 2560 207
rect 2544 7 2560 202
rect 2845 102 2850 777
rect 2941 732 2946 1217
rect 2877 622 2882 667
rect 2973 622 2978 1757
rect 2989 772 2994 1747
rect 3048 1707 3064 1902
rect 3053 1702 3058 1707
rect 3063 1702 3064 1707
rect 3048 1507 3064 1702
rect 3568 4407 3584 4430
rect 3573 4402 3578 4407
rect 3583 4402 3584 4407
rect 3568 4207 3584 4402
rect 3573 4202 3578 4207
rect 3583 4202 3584 4207
rect 3568 4007 3584 4202
rect 3573 4002 3578 4007
rect 3583 4002 3584 4007
rect 3568 3807 3584 4002
rect 3573 3802 3578 3807
rect 3583 3802 3584 3807
rect 3568 3607 3584 3802
rect 3573 3602 3578 3607
rect 3583 3602 3584 3607
rect 3568 3407 3584 3602
rect 3573 3402 3578 3407
rect 3583 3402 3584 3407
rect 3568 3207 3584 3402
rect 3573 3202 3578 3207
rect 3583 3202 3584 3207
rect 3568 3007 3584 3202
rect 3573 3002 3578 3007
rect 3583 3002 3584 3007
rect 3568 2807 3584 3002
rect 4080 4307 4096 4430
rect 4085 4302 4090 4307
rect 4095 4302 4096 4307
rect 4080 4107 4096 4302
rect 4085 4102 4090 4107
rect 4095 4102 4096 4107
rect 4080 3907 4096 4102
rect 4085 3902 4090 3907
rect 4095 3902 4096 3907
rect 4080 3707 4096 3902
rect 4085 3702 4090 3707
rect 4095 3702 4096 3707
rect 4080 3507 4096 3702
rect 4085 3502 4090 3507
rect 4095 3502 4096 3507
rect 4080 3307 4096 3502
rect 4085 3302 4090 3307
rect 4095 3302 4096 3307
rect 4080 3107 4096 3302
rect 4085 3102 4090 3107
rect 4095 3102 4096 3107
rect 4080 2907 4096 3102
rect 4085 2902 4090 2907
rect 4095 2902 4096 2907
rect 3573 2802 3578 2807
rect 3583 2802 3584 2807
rect 3568 2607 3584 2802
rect 3573 2602 3578 2607
rect 3583 2602 3584 2607
rect 3568 2407 3584 2602
rect 3573 2402 3578 2407
rect 3583 2402 3584 2407
rect 3568 2207 3584 2402
rect 3573 2202 3578 2207
rect 3583 2202 3584 2207
rect 3568 2007 3584 2202
rect 3573 2002 3578 2007
rect 3583 2002 3584 2007
rect 3568 1807 3584 2002
rect 3573 1802 3578 1807
rect 3583 1802 3584 1807
rect 3568 1607 3584 1802
rect 3573 1602 3578 1607
rect 3583 1602 3584 1607
rect 3053 1502 3058 1507
rect 3063 1502 3064 1507
rect 3048 1307 3064 1502
rect 3053 1302 3058 1307
rect 3063 1302 3064 1307
rect 3048 1107 3064 1302
rect 3069 1112 3074 1167
rect 3053 1102 3058 1107
rect 3063 1102 3064 1107
rect 3048 907 3064 1102
rect 3053 902 3058 907
rect 3063 902 3064 907
rect 3048 707 3064 902
rect 3053 702 3058 707
rect 3063 702 3064 707
rect 3048 507 3064 702
rect 3053 502 3058 507
rect 3063 502 3064 507
rect 3048 307 3064 502
rect 3069 482 3074 497
rect 3085 402 3090 1467
rect 3117 902 3122 1157
rect 3181 882 3186 937
rect 3213 892 3218 1187
rect 3453 792 3458 1537
rect 3517 812 3522 1537
rect 3568 1407 3584 1602
rect 3573 1402 3578 1407
rect 3583 1402 3584 1407
rect 3568 1207 3584 1402
rect 3573 1202 3578 1207
rect 3583 1202 3584 1207
rect 3568 1007 3584 1202
rect 3573 1002 3578 1007
rect 3583 1002 3584 1007
rect 3568 807 3584 1002
rect 3573 802 3578 807
rect 3583 802 3584 807
rect 3568 607 3584 802
rect 3573 602 3578 607
rect 3583 602 3584 607
rect 3293 312 3298 447
rect 3568 407 3584 602
rect 3573 402 3578 407
rect 3583 402 3584 407
rect 3053 302 3058 307
rect 3063 302 3064 307
rect 3048 107 3064 302
rect 3309 282 3314 307
rect 3053 102 3058 107
rect 3063 102 3064 107
rect 2549 2 2554 7
rect 2559 2 2560 7
rect 2544 -30 2560 2
rect 3048 -30 3064 102
rect 3568 207 3584 402
rect 3573 202 3578 207
rect 3583 202 3584 207
rect 3568 7 3584 202
rect 3645 162 3650 2337
rect 3661 692 3666 2517
rect 3709 92 3714 1887
rect 3725 1012 3730 2357
rect 3741 962 3746 2527
rect 3741 482 3746 957
rect 3805 92 3810 2567
rect 3821 282 3826 1267
rect 3837 272 3842 1077
rect 3853 212 3858 2547
rect 3869 202 3874 1587
rect 3837 82 3842 97
rect 3853 82 3858 197
rect 3885 12 3890 1397
rect 3901 72 3906 1287
rect 3917 282 3922 1567
rect 3949 992 3954 2877
rect 4080 2707 4096 2902
rect 4085 2702 4090 2707
rect 4095 2702 4096 2707
rect 4080 2507 4096 2702
rect 4085 2502 4090 2507
rect 4095 2502 4096 2507
rect 4080 2307 4096 2502
rect 4085 2302 4090 2307
rect 4095 2302 4096 2307
rect 4080 2107 4096 2302
rect 4085 2102 4090 2107
rect 4095 2102 4096 2107
rect 4080 1907 4096 2102
rect 4085 1902 4090 1907
rect 4095 1902 4096 1907
rect 4080 1707 4096 1902
rect 4085 1702 4090 1707
rect 4095 1702 4096 1707
rect 3933 72 3938 427
rect 3949 212 3954 767
rect 3965 302 3970 1397
rect 3981 272 3986 1687
rect 3930 67 3938 72
rect 4029 12 4034 1517
rect 4080 1507 4096 1702
rect 4085 1502 4090 1507
rect 4095 1502 4096 1507
rect 4080 1307 4096 1502
rect 4085 1302 4090 1307
rect 4095 1302 4096 1307
rect 4080 1107 4096 1302
rect 4085 1102 4090 1107
rect 4095 1102 4096 1107
rect 4045 112 4050 967
rect 4080 907 4096 1102
rect 4125 1032 4130 1077
rect 4085 902 4090 907
rect 4095 902 4096 907
rect 4080 707 4096 902
rect 4085 702 4090 707
rect 4095 702 4096 707
rect 4061 152 4066 657
rect 4080 507 4096 702
rect 4141 682 4146 1787
rect 4085 502 4090 507
rect 4095 502 4096 507
rect 4080 307 4096 502
rect 4085 302 4090 307
rect 4095 302 4096 307
rect 4080 107 4096 302
rect 4085 102 4090 107
rect 4095 102 4096 107
rect 3573 2 3578 7
rect 3583 2 3584 7
rect 3568 -30 3584 2
rect 4080 -30 4096 102
rect 4125 72 4130 277
rect 4157 52 4162 1607
rect 4173 722 4178 2227
rect 4189 402 4194 1107
rect 4205 812 4210 1557
rect 4237 1072 4242 1607
rect 4205 62 4210 537
rect 4221 172 4226 677
rect 4253 112 4258 127
rect 4269 42 4274 2337
rect 4381 1372 4386 4327
rect 4349 152 4354 1357
rect 4381 132 4386 1197
rect 4397 722 4402 1547
rect 4429 632 4434 3467
rect 4445 2342 4450 4347
rect 4461 1642 4466 4287
rect 4477 2812 4482 4347
rect 4477 282 4482 2707
rect 4509 1462 4514 3817
rect 4525 322 4530 2257
rect 4541 1532 4546 4107
rect 4541 152 4546 937
rect 4557 542 4562 4087
rect 4557 22 4562 537
rect 4573 1392 4578 4307
rect 4573 472 4578 1387
rect 4589 522 4594 3237
use BUFX2  BUFX2_49
timestamp 1693479267
transform -1 0 28 0 -1 105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_7
timestamp 1693479267
transform -1 0 100 0 -1 105
box -2 -3 74 103
use BUFX2  BUFX2_71
timestamp 1693479267
transform -1 0 124 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_482
timestamp 1693479267
transform -1 0 100 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_480
timestamp 1693479267
transform -1 0 196 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_448
timestamp 1693479267
transform 1 0 124 0 -1 105
box -2 -3 98 103
use NAND3X1  NAND3X1_23
timestamp 1693479267
transform 1 0 196 0 1 105
box -2 -3 34 103
use BUFX2  BUFX2_13
timestamp 1693479267
transform -1 0 244 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_170
timestamp 1693479267
transform -1 0 340 0 -1 105
box -2 -3 98 103
use NAND3X1  NAND3X1_22
timestamp 1693479267
transform 1 0 228 0 1 105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_41
timestamp 1693479267
transform 1 0 260 0 1 105
box -2 -3 74 103
use BUFX2  BUFX2_51
timestamp 1693479267
transform -1 0 364 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_452
timestamp 1693479267
transform 1 0 364 0 -1 105
box -2 -3 98 103
use NAND3X1  NAND3X1_30
timestamp 1693479267
transform -1 0 364 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_31
timestamp 1693479267
transform 1 0 364 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_484
timestamp 1693479267
transform 1 0 396 0 1 105
box -2 -3 98 103
use BUFX2  BUFX2_45
timestamp 1693479267
transform 1 0 460 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_17
timestamp 1693479267
transform -1 0 508 0 -1 105
box -2 -3 26 103
use FILL  FILL_0_0_0
timestamp 1693479267
transform -1 0 516 0 -1 105
box -2 -3 10 103
use FILL  FILL_1_0_0
timestamp 1693479267
transform 1 0 492 0 1 105
box -2 -3 10 103
use FILL  FILL_1_0_1
timestamp 1693479267
transform 1 0 500 0 1 105
box -2 -3 10 103
use BUFX2  BUFX2_46
timestamp 1693479267
transform 1 0 508 0 1 105
box -2 -3 26 103
use FILL  FILL_0_0_1
timestamp 1693479267
transform -1 0 524 0 -1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_174
timestamp 1693479267
transform -1 0 620 0 -1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_661
timestamp 1693479267
transform 1 0 532 0 1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_389
timestamp 1693479267
transform 1 0 556 0 1 105
box -2 -3 26 103
use OR2X2  OR2X2_47
timestamp 1693479267
transform -1 0 612 0 1 105
box -2 -3 34 103
use BUFX2  BUFX2_52
timestamp 1693479267
transform 1 0 620 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_453
timestamp 1693479267
transform 1 0 644 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_837
timestamp 1693479267
transform 1 0 612 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_834
timestamp 1693479267
transform 1 0 644 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_660
timestamp 1693479267
transform -1 0 700 0 1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_387
timestamp 1693479267
transform -1 0 724 0 1 105
box -2 -3 26 103
use BUFX2  BUFX2_41
timestamp 1693479267
transform -1 0 764 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_42
timestamp 1693479267
transform -1 0 788 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_665
timestamp 1693479267
transform -1 0 812 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_477
timestamp 1693479267
transform -1 0 740 0 1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_485
timestamp 1693479267
transform -1 0 836 0 1 105
box -2 -3 98 103
use BUFX2  BUFX2_54
timestamp 1693479267
transform -1 0 836 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_455
timestamp 1693479267
transform 1 0 836 0 -1 105
box -2 -3 98 103
use NAND3X1  NAND3X1_32
timestamp 1693479267
transform 1 0 836 0 1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_216
timestamp 1693479267
transform 1 0 868 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_838
timestamp 1693479267
transform 1 0 900 0 1 105
box -2 -3 34 103
use BUFX2  BUFX2_53
timestamp 1693479267
transform 1 0 932 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_43
timestamp 1693479267
transform 1 0 956 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_44
timestamp 1693479267
transform 1 0 980 0 -1 105
box -2 -3 26 103
use FILL  FILL_0_1_0
timestamp 1693479267
transform 1 0 1004 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_1_1
timestamp 1693479267
transform 1 0 1012 0 -1 105
box -2 -3 10 103
use NAND3X1  NAND3X1_36
timestamp 1693479267
transform -1 0 964 0 1 105
box -2 -3 34 103
use FILL  FILL_1_1_0
timestamp 1693479267
transform -1 0 972 0 1 105
box -2 -3 10 103
use FILL  FILL_1_1_1
timestamp 1693479267
transform -1 0 980 0 1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_487
timestamp 1693479267
transform -1 0 1076 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_486
timestamp 1693479267
transform 1 0 1020 0 -1 105
box -2 -3 98 103
use NAND3X1  NAND3X1_34
timestamp 1693479267
transform -1 0 1108 0 1 105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_51
timestamp 1693479267
transform 1 0 1108 0 1 105
box -2 -3 58 103
use BUFX2  BUFX2_9
timestamp 1693479267
transform -1 0 1140 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_168
timestamp 1693479267
transform 1 0 1140 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_836
timestamp 1693479267
transform 1 0 1164 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_663
timestamp 1693479267
transform -1 0 1220 0 1 105
box -2 -3 26 103
use BUFX2  BUFX2_11
timestamp 1693479267
transform 1 0 1236 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_171
timestamp 1693479267
transform 1 0 1260 0 -1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_664
timestamp 1693479267
transform 1 0 1220 0 1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_454
timestamp 1693479267
transform 1 0 1244 0 1 105
box -2 -3 98 103
use BUFX2  BUFX2_14
timestamp 1693479267
transform 1 0 1356 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_8
timestamp 1693479267
transform 1 0 1380 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_10
timestamp 1693479267
transform 1 0 1404 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_48
timestamp 1693479267
transform 1 0 1340 0 1 105
box -2 -3 26 103
use BUFX2  BUFX2_5
timestamp 1693479267
transform 1 0 1364 0 1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_167
timestamp 1693479267
transform -1 0 1484 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_172
timestamp 1693479267
transform 1 0 1428 0 -1 105
box -2 -3 98 103
use FILL  FILL_1_2_0
timestamp 1693479267
transform 1 0 1484 0 1 105
box -2 -3 10 103
use FILL  FILL_1_2_1
timestamp 1693479267
transform 1 0 1492 0 1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_173
timestamp 1693479267
transform 1 0 1500 0 1 105
box -2 -3 98 103
use FILL  FILL_0_2_0
timestamp 1693479267
transform 1 0 1524 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_2_1
timestamp 1693479267
transform 1 0 1532 0 -1 105
box -2 -3 10 103
use BUFX2  BUFX2_15
timestamp 1693479267
transform 1 0 1540 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_16
timestamp 1693479267
transform 1 0 1564 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_267
timestamp 1693479267
transform 1 0 1588 0 -1 105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_14
timestamp 1693479267
transform 1 0 1596 0 1 105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_269
timestamp 1693479267
transform 1 0 1684 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_262
timestamp 1693479267
transform 1 0 1668 0 1 105
box -2 -3 98 103
use MUX2X1  MUX2X1_3
timestamp 1693479267
transform -1 0 1828 0 -1 105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_266
timestamp 1693479267
transform 1 0 1764 0 1 105
box -2 -3 98 103
use INVX1  INVX1_330
timestamp 1693479267
transform 1 0 1828 0 -1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_307
timestamp 1693479267
transform 1 0 1844 0 -1 105
box -2 -3 34 103
use INVX1  INVX1_342
timestamp 1693479267
transform -1 0 1892 0 -1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_279
timestamp 1693479267
transform 1 0 1892 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_282
timestamp 1693479267
transform 1 0 1916 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_241
timestamp 1693479267
transform -1 0 1884 0 1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_268
timestamp 1693479267
transform 1 0 1884 0 1 105
box -2 -3 98 103
use NOR2X1  NOR2X1_146
timestamp 1693479267
transform -1 0 1964 0 -1 105
box -2 -3 26 103
use INVX2  INVX2_46
timestamp 1693479267
transform -1 0 1980 0 -1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_448
timestamp 1693479267
transform 1 0 1980 0 -1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_244
timestamp 1693479267
transform 1 0 2004 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_343
timestamp 1693479267
transform 1 0 1980 0 1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_321
timestamp 1693479267
transform 1 0 1996 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_280
timestamp 1693479267
transform -1 0 2068 0 1 105
box -2 -3 26 103
use FILL  FILL_1_3_1
timestamp 1693479267
transform -1 0 2044 0 1 105
box -2 -3 10 103
use FILL  FILL_1_3_0
timestamp 1693479267
transform -1 0 2036 0 1 105
box -2 -3 10 103
use AND2X2  AND2X2_37
timestamp 1693479267
transform -1 0 2076 0 -1 105
box -2 -3 34 103
use FILL  FILL_0_3_1
timestamp 1693479267
transform -1 0 2044 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_3_0
timestamp 1693479267
transform -1 0 2036 0 -1 105
box -2 -3 10 103
use OAI22X1  OAI22X1_22
timestamp 1693479267
transform -1 0 2140 0 -1 105
box -2 -3 42 103
use NOR2X1  NOR2X1_245
timestamp 1693479267
transform 1 0 2076 0 -1 105
box -2 -3 26 103
use MUX2X1  MUX2X1_15
timestamp 1693479267
transform -1 0 2164 0 1 105
box -2 -3 50 103
use MUX2X1  MUX2X1_16
timestamp 1693479267
transform 1 0 2068 0 1 105
box -2 -3 50 103
use NOR2X1  NOR2X1_243
timestamp 1693479267
transform -1 0 2164 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_111
timestamp 1693479267
transform -1 0 2196 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_291
timestamp 1693479267
transform -1 0 2220 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_281
timestamp 1693479267
transform 1 0 2220 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_277
timestamp 1693479267
transform -1 0 2188 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_320
timestamp 1693479267
transform -1 0 2220 0 1 105
box -2 -3 34 103
use INVX1  INVX1_341
timestamp 1693479267
transform -1 0 2236 0 1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_4
timestamp 1693479267
transform 1 0 2244 0 -1 105
box -2 -3 50 103
use NAND2X1  NAND2X1_244
timestamp 1693479267
transform -1 0 2316 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_308
timestamp 1693479267
transform -1 0 2348 0 -1 105
box -2 -3 34 103
use AOI22X1  AOI22X1_74
timestamp 1693479267
transform -1 0 2276 0 1 105
box -2 -3 42 103
use NAND2X1  NAND2X1_278
timestamp 1693479267
transform -1 0 2300 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_511
timestamp 1693479267
transform -1 0 2332 0 1 105
box -2 -3 34 103
use INVX1  INVX1_331
timestamp 1693479267
transform -1 0 2364 0 -1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_156
timestamp 1693479267
transform -1 0 2388 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_51
timestamp 1693479267
transform 1 0 2388 0 -1 105
box -2 -3 34 103
use BUFX4  BUFX4_41
timestamp 1693479267
transform -1 0 2452 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_145
timestamp 1693479267
transform 1 0 2332 0 1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_144
timestamp 1693479267
transform -1 0 2380 0 1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_449
timestamp 1693479267
transform -1 0 2404 0 1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_293
timestamp 1693479267
transform 1 0 2404 0 1 105
box -2 -3 26 103
use BUFX4  BUFX4_43
timestamp 1693479267
transform 1 0 2452 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_328
timestamp 1693479267
transform -1 0 2508 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_347
timestamp 1693479267
transform -1 0 2540 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_502
timestamp 1693479267
transform 1 0 2428 0 1 105
box -2 -3 34 103
use AOI22X1  AOI22X1_89
timestamp 1693479267
transform -1 0 2500 0 1 105
box -2 -3 42 103
use NAND2X1  NAND2X1_294
timestamp 1693479267
transform -1 0 2524 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_324
timestamp 1693479267
transform 1 0 2524 0 1 105
box -2 -3 34 103
use FILL  FILL_1_4_1
timestamp 1693479267
transform -1 0 2572 0 1 105
box -2 -3 10 103
use FILL  FILL_1_4_0
timestamp 1693479267
transform -1 0 2564 0 1 105
box -2 -3 10 103
use NAND2X1  NAND2X1_386
timestamp 1693479267
transform 1 0 2556 0 -1 105
box -2 -3 26 103
use FILL  FILL_0_4_1
timestamp 1693479267
transform 1 0 2548 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_4_0
timestamp 1693479267
transform 1 0 2540 0 -1 105
box -2 -3 10 103
use AOI21X1  AOI21X1_96
timestamp 1693479267
transform -1 0 2628 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_292
timestamp 1693479267
transform -1 0 2596 0 1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_329
timestamp 1693479267
transform 1 0 2580 0 -1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_166
timestamp 1693479267
transform -1 0 2652 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_403
timestamp 1693479267
transform 1 0 2628 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_400
timestamp 1693479267
transform -1 0 2628 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_387
timestamp 1693479267
transform 1 0 2660 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_368
timestamp 1693479267
transform 1 0 2684 0 -1 105
box -2 -3 18 103
use BUFX4  BUFX4_42
timestamp 1693479267
transform 1 0 2700 0 -1 105
box -2 -3 34 103
use MUX2X1  MUX2X1_31
timestamp 1693479267
transform -1 0 2700 0 1 105
box -2 -3 50 103
use NAND2X1  NAND2X1_381
timestamp 1693479267
transform -1 0 2724 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_396
timestamp 1693479267
transform 1 0 2724 0 1 105
box -2 -3 34 103
use INVX1  INVX1_333
timestamp 1693479267
transform 1 0 2732 0 -1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_310
timestamp 1693479267
transform 1 0 2748 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_248
timestamp 1693479267
transform 1 0 2780 0 -1 105
box -2 -3 26 103
use MUX2X1  MUX2X1_6
timestamp 1693479267
transform 1 0 2804 0 -1 105
box -2 -3 50 103
use OAI21X1  OAI21X1_395
timestamp 1693479267
transform -1 0 2788 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_415
timestamp 1693479267
transform 1 0 2788 0 1 105
box -2 -3 26 103
use INVX1  INVX1_366
timestamp 1693479267
transform 1 0 2812 0 1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_397
timestamp 1693479267
transform 1 0 2828 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_348
timestamp 1693479267
transform 1 0 2852 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_330
timestamp 1693479267
transform 1 0 2884 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_353
timestamp 1693479267
transform 1 0 2908 0 -1 105
box -2 -3 18 103
use INVX1  INVX1_332
timestamp 1693479267
transform 1 0 2924 0 -1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_382
timestamp 1693479267
transform 1 0 2860 0 1 105
box -2 -3 26 103
use INVX8  INVX8_8
timestamp 1693479267
transform -1 0 2924 0 1 105
box -2 -3 42 103
use NAND2X1  NAND2X1_416
timestamp 1693479267
transform -1 0 2948 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_309
timestamp 1693479267
transform 1 0 2940 0 -1 105
box -2 -3 34 103
use OR2X2  OR2X2_21
timestamp 1693479267
transform 1 0 2972 0 -1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_100
timestamp 1693479267
transform -1 0 3036 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_418
timestamp 1693479267
transform 1 0 2948 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_364
timestamp 1693479267
transform 1 0 2980 0 1 105
box -2 -3 34 103
use INVX1  INVX1_354
timestamp 1693479267
transform 1 0 3012 0 1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_414
timestamp 1693479267
transform -1 0 3060 0 1 105
box -2 -3 34 103
use FILL  FILL_1_5_1
timestamp 1693479267
transform 1 0 3068 0 1 105
box -2 -3 10 103
use FILL  FILL_1_5_0
timestamp 1693479267
transform 1 0 3060 0 1 105
box -2 -3 10 103
use FILL  FILL_0_5_1
timestamp 1693479267
transform -1 0 3076 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_5_0
timestamp 1693479267
transform -1 0 3068 0 -1 105
box -2 -3 10 103
use NAND2X1  NAND2X1_304
timestamp 1693479267
transform 1 0 3036 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_402
timestamp 1693479267
transform 1 0 3076 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_250
timestamp 1693479267
transform 1 0 3100 0 -1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_287
timestamp 1693479267
transform -1 0 3100 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_349
timestamp 1693479267
transform -1 0 3140 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_117
timestamp 1693479267
transform -1 0 3148 0 -1 105
box -2 -3 26 103
use INVX2  INVX2_41
timestamp 1693479267
transform -1 0 3164 0 -1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_499
timestamp 1693479267
transform 1 0 3164 0 -1 105
box -2 -3 26 103
use INVX2  INVX2_40
timestamp 1693479267
transform -1 0 3204 0 -1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_510
timestamp 1693479267
transform 1 0 3204 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_303
timestamp 1693479267
transform 1 0 3228 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_402
timestamp 1693479267
transform -1 0 3164 0 1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_404
timestamp 1693479267
transform 1 0 3164 0 1 105
box -2 -3 26 103
use OR2X2  OR2X2_19
timestamp 1693479267
transform 1 0 3188 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_351
timestamp 1693479267
transform 1 0 3220 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_285
timestamp 1693479267
transform -1 0 3276 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_305
timestamp 1693479267
transform 1 0 3276 0 -1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_170
timestamp 1693479267
transform -1 0 3324 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_249
timestamp 1693479267
transform 1 0 3324 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_583
timestamp 1693479267
transform -1 0 3284 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_433
timestamp 1693479267
transform 1 0 3284 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_432
timestamp 1693479267
transform -1 0 3348 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_112
timestamp 1693479267
transform 1 0 3348 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_242
timestamp 1693479267
transform -1 0 3396 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_245
timestamp 1693479267
transform 1 0 3396 0 -1 105
box -2 -3 26 103
use INVX2  INVX2_38
timestamp 1693479267
transform 1 0 3420 0 -1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_524
timestamp 1693479267
transform -1 0 3460 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_399
timestamp 1693479267
transform -1 0 3380 0 1 105
box -2 -3 34 103
use MUX2X1  MUX2X1_37
timestamp 1693479267
transform -1 0 3428 0 1 105
box -2 -3 50 103
use AOI21X1  AOI21X1_120
timestamp 1693479267
transform 1 0 3428 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_291
timestamp 1693479267
transform -1 0 3484 0 -1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_111
timestamp 1693479267
transform 1 0 3484 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_243
timestamp 1693479267
transform 1 0 3508 0 -1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_127
timestamp 1693479267
transform -1 0 3556 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_526
timestamp 1693479267
transform -1 0 3484 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_584
timestamp 1693479267
transform -1 0 3516 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_247
timestamp 1693479267
transform -1 0 3540 0 1 105
box -2 -3 26 103
use FILL  FILL_1_6_0
timestamp 1693479267
transform 1 0 3588 0 1 105
box -2 -3 10 103
use FILL  FILL_0_6_1
timestamp 1693479267
transform 1 0 3588 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_6_0
timestamp 1693479267
transform 1 0 3580 0 -1 105
box -2 -3 10 103
use NAND2X1  NAND2X1_306
timestamp 1693479267
transform 1 0 3556 0 -1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_192
timestamp 1693479267
transform 1 0 3628 0 1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_118
timestamp 1693479267
transform 1 0 3604 0 1 105
box -2 -3 26 103
use FILL  FILL_1_6_1
timestamp 1693479267
transform 1 0 3596 0 1 105
box -2 -3 10 103
use NOR2X1  NOR2X1_303
timestamp 1693479267
transform 1 0 3636 0 -1 105
box -2 -3 26 103
use INVX2  INVX2_39
timestamp 1693479267
transform 1 0 3620 0 -1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_307
timestamp 1693479267
transform 1 0 3596 0 -1 105
box -2 -3 26 103
use MUX2X1  MUX2X1_36
timestamp 1693479267
transform -1 0 3588 0 1 105
box -2 -3 50 103
use NAND2X1  NAND2X1_518
timestamp 1693479267
transform -1 0 3684 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_246
timestamp 1693479267
transform 1 0 3684 0 -1 105
box -2 -3 26 103
use MUX2X1  MUX2X1_50
timestamp 1693479267
transform 1 0 3708 0 -1 105
box -2 -3 50 103
use MUX2X1  MUX2X1_5
timestamp 1693479267
transform -1 0 3700 0 1 105
box -2 -3 50 103
use OAI21X1  OAI21X1_606
timestamp 1693479267
transform -1 0 3732 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_105
timestamp 1693479267
transform -1 0 3756 0 1 105
box -2 -3 26 103
use OR2X2  OR2X2_58
timestamp 1693479267
transform 1 0 3756 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_753
timestamp 1693479267
transform 1 0 3788 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_953
timestamp 1693479267
transform -1 0 3852 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_115
timestamp 1693479267
transform 1 0 3756 0 1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_106
timestamp 1693479267
transform 1 0 3780 0 1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_302
timestamp 1693479267
transform 1 0 3804 0 1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_107
timestamp 1693479267
transform -1 0 3852 0 1 105
box -2 -3 26 103
use AOI22X1  AOI22X1_155
timestamp 1693479267
transform -1 0 3892 0 -1 105
box -2 -3 42 103
use OAI22X1  OAI22X1_23
timestamp 1693479267
transform -1 0 3932 0 -1 105
box -2 -3 42 103
use OAI21X1  OAI21X1_521
timestamp 1693479267
transform -1 0 3964 0 -1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_90
timestamp 1693479267
transform 1 0 3852 0 1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_145
timestamp 1693479267
transform 1 0 3884 0 1 105
box -2 -3 34 103
use OAI22X1  OAI22X1_31
timestamp 1693479267
transform -1 0 3956 0 1 105
box -2 -3 42 103
use OAI21X1  OAI21X1_971
timestamp 1693479267
transform -1 0 3996 0 -1 105
box -2 -3 34 103
use BUFX4  BUFX4_117
timestamp 1693479267
transform 1 0 3996 0 -1 105
box -2 -3 34 103
use OAI22X1  OAI22X1_34
timestamp 1693479267
transform -1 0 4068 0 -1 105
box -2 -3 42 103
use AOI21X1  AOI21X1_121
timestamp 1693479267
transform -1 0 3988 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_330
timestamp 1693479267
transform -1 0 4020 0 1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_42
timestamp 1693479267
transform 1 0 4020 0 1 105
box -2 -3 34 103
use FILL  FILL_1_7_1
timestamp 1693479267
transform 1 0 4084 0 1 105
box -2 -3 10 103
use FILL  FILL_1_7_0
timestamp 1693479267
transform 1 0 4076 0 1 105
box -2 -3 10 103
use NAND2X1  NAND2X1_251
timestamp 1693479267
transform -1 0 4076 0 1 105
box -2 -3 26 103
use FILL  FILL_0_7_0
timestamp 1693479267
transform -1 0 4092 0 -1 105
box -2 -3 10 103
use INVX1  INVX1_729
timestamp 1693479267
transform 1 0 4068 0 -1 105
box -2 -3 18 103
use AOI22X1  AOI22X1_70
timestamp 1693479267
transform -1 0 4164 0 1 105
box -2 -3 42 103
use OAI21X1  OAI21X1_588
timestamp 1693479267
transform 1 0 4092 0 1 105
box -2 -3 34 103
use AND2X2  AND2X2_41
timestamp 1693479267
transform 1 0 4116 0 -1 105
box -2 -3 34 103
use INVX1  INVX1_739
timestamp 1693479267
transform -1 0 4116 0 -1 105
box -2 -3 18 103
use FILL  FILL_0_7_1
timestamp 1693479267
transform -1 0 4100 0 -1 105
box -2 -3 10 103
use AOI22X1  AOI22X1_98
timestamp 1693479267
transform -1 0 4188 0 -1 105
box -2 -3 42 103
use INVX8  INVX8_7
timestamp 1693479267
transform 1 0 4188 0 -1 105
box -2 -3 42 103
use OAI21X1  OAI21X1_1039
timestamp 1693479267
transform -1 0 4260 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_589
timestamp 1693479267
transform -1 0 4196 0 1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_122
timestamp 1693479267
transform 1 0 4196 0 1 105
box -2 -3 34 103
use OAI22X1  OAI22X1_7
timestamp 1693479267
transform 1 0 4228 0 1 105
box -2 -3 42 103
use OR2X2  OR2X2_30
timestamp 1693479267
transform -1 0 4292 0 -1 105
box -2 -3 34 103
use BUFX4  BUFX4_127
timestamp 1693479267
transform 1 0 4292 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_280
timestamp 1693479267
transform 1 0 4324 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_143
timestamp 1693479267
transform -1 0 4300 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_113
timestamp 1693479267
transform 1 0 4300 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_607
timestamp 1693479267
transform -1 0 4356 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_373
timestamp 1693479267
transform 1 0 4348 0 -1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_288
timestamp 1693479267
transform -1 0 4396 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_577
timestamp 1693479267
transform 1 0 4396 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_522
timestamp 1693479267
transform -1 0 4452 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_331
timestamp 1693479267
transform 1 0 4356 0 1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_133
timestamp 1693479267
transform 1 0 4388 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_292
timestamp 1693479267
transform -1 0 4444 0 1 105
box -2 -3 26 103
use OAI22X1  OAI22X1_38
timestamp 1693479267
transform -1 0 4484 0 1 105
box -2 -3 42 103
use NAND2X1  NAND2X1_523
timestamp 1693479267
transform 1 0 4452 0 -1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_216
timestamp 1693479267
transform 1 0 4476 0 -1 105
box -2 -3 26 103
use BUFX4  BUFX4_173
timestamp 1693479267
transform -1 0 4532 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_290
timestamp 1693479267
transform 1 0 4532 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_580
timestamp 1693479267
transform 1 0 4484 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_114
timestamp 1693479267
transform -1 0 4540 0 1 105
box -2 -3 26 103
use BUFX4  BUFX4_254
timestamp 1693479267
transform 1 0 4540 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_578
timestamp 1693479267
transform 1 0 4556 0 -1 105
box -2 -3 34 103
use FILL  FILL_1_1
timestamp 1693479267
transform -1 0 4596 0 -1 105
box -2 -3 10 103
use FILL  FILL_1_2
timestamp 1693479267
transform -1 0 4604 0 -1 105
box -2 -3 10 103
use FILL  FILL_2_1
timestamp 1693479267
transform 1 0 4572 0 1 105
box -2 -3 10 103
use FILL  FILL_2_2
timestamp 1693479267
transform 1 0 4580 0 1 105
box -2 -3 10 103
use FILL  FILL_2_3
timestamp 1693479267
transform 1 0 4588 0 1 105
box -2 -3 10 103
use FILL  FILL_2_4
timestamp 1693479267
transform 1 0 4596 0 1 105
box -2 -3 10 103
use BUFX2  BUFX2_47
timestamp 1693479267
transform -1 0 28 0 -1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_450
timestamp 1693479267
transform 1 0 28 0 -1 305
box -2 -3 98 103
use AOI21X1  AOI21X1_215
timestamp 1693479267
transform -1 0 156 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_829
timestamp 1693479267
transform 1 0 156 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_171
timestamp 1693479267
transform -1 0 220 0 -1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_27
timestamp 1693479267
transform -1 0 252 0 -1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_26
timestamp 1693479267
transform 1 0 252 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_169
timestamp 1693479267
transform 1 0 284 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_653
timestamp 1693479267
transform 1 0 316 0 -1 305
box -2 -3 26 103
use NAND3X1  NAND3X1_182
timestamp 1693479267
transform -1 0 372 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_173
timestamp 1693479267
transform 1 0 372 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_659
timestamp 1693479267
transform 1 0 404 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_833
timestamp 1693479267
transform -1 0 460 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_658
timestamp 1693479267
transform -1 0 484 0 -1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_385
timestamp 1693479267
transform 1 0 484 0 -1 305
box -2 -3 26 103
use FILL  FILL_2_0_0
timestamp 1693479267
transform 1 0 508 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_0_1
timestamp 1693479267
transform 1 0 516 0 -1 305
box -2 -3 10 103
use INVX1  INVX1_476
timestamp 1693479267
transform 1 0 524 0 -1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_649
timestamp 1693479267
transform 1 0 540 0 -1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_383
timestamp 1693479267
transform -1 0 588 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_826
timestamp 1693479267
transform 1 0 588 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_650
timestamp 1693479267
transform -1 0 644 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_655
timestamp 1693479267
transform 1 0 644 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_835
timestamp 1693479267
transform 1 0 668 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_662
timestamp 1693479267
transform 1 0 700 0 -1 305
box -2 -3 26 103
use XOR2X1  XOR2X1_8
timestamp 1693479267
transform 1 0 724 0 -1 305
box -2 -3 58 103
use OAI21X1  OAI21X1_174
timestamp 1693479267
transform -1 0 812 0 -1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_33
timestamp 1693479267
transform -1 0 844 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_827
timestamp 1693479267
transform 1 0 844 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_170
timestamp 1693479267
transform -1 0 908 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_176
timestamp 1693479267
transform -1 0 940 0 -1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_37
timestamp 1693479267
transform -1 0 972 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_175
timestamp 1693479267
transform 1 0 972 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_1_0
timestamp 1693479267
transform -1 0 1012 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_1_1
timestamp 1693479267
transform -1 0 1020 0 -1 305
box -2 -3 10 103
use NAND3X1  NAND3X1_35
timestamp 1693479267
transform -1 0 1052 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_652
timestamp 1693479267
transform -1 0 1076 0 -1 305
box -2 -3 26 103
use NAND3X1  NAND3X1_24
timestamp 1693479267
transform -1 0 1108 0 -1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_25
timestamp 1693479267
transform 1 0 1108 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_481
timestamp 1693479267
transform 1 0 1140 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_449
timestamp 1693479267
transform 1 0 1236 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_263
timestamp 1693479267
transform 1 0 1332 0 -1 305
box -2 -3 98 103
use XNOR2X1  XNOR2X1_35
timestamp 1693479267
transform 1 0 1428 0 -1 305
box -2 -3 58 103
use CLKBUF1  CLKBUF1_26
timestamp 1693479267
transform -1 0 1556 0 -1 305
box -2 -3 74 103
use FILL  FILL_2_2_0
timestamp 1693479267
transform 1 0 1556 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_2_1
timestamp 1693479267
transform 1 0 1564 0 -1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_264
timestamp 1693479267
transform 1 0 1572 0 -1 305
box -2 -3 98 103
use XNOR2X1  XNOR2X1_34
timestamp 1693479267
transform -1 0 1724 0 -1 305
box -2 -3 58 103
use NOR2X1  NOR2X1_40
timestamp 1693479267
transform -1 0 1748 0 -1 305
box -2 -3 26 103
use INVX2  INVX2_13
timestamp 1693479267
transform 1 0 1748 0 -1 305
box -2 -3 18 103
use XNOR2X1  XNOR2X1_44
timestamp 1693479267
transform -1 0 1820 0 -1 305
box -2 -3 58 103
use AOI22X1  AOI22X1_52
timestamp 1693479267
transform -1 0 1860 0 -1 305
box -2 -3 42 103
use AOI22X1  AOI22X1_50
timestamp 1693479267
transform 1 0 1860 0 -1 305
box -2 -3 42 103
use AOI22X1  AOI22X1_51
timestamp 1693479267
transform -1 0 1940 0 -1 305
box -2 -3 42 103
use NOR2X1  NOR2X1_96
timestamp 1693479267
transform -1 0 1964 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_237
timestamp 1693479267
transform -1 0 1988 0 -1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_98
timestamp 1693479267
transform 1 0 1988 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_236
timestamp 1693479267
transform -1 0 2036 0 -1 305
box -2 -3 26 103
use FILL  FILL_2_3_0
timestamp 1693479267
transform -1 0 2044 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_3_1
timestamp 1693479267
transform -1 0 2052 0 -1 305
box -2 -3 10 103
use NOR2X1  NOR2X1_312
timestamp 1693479267
transform -1 0 2076 0 -1 305
box -2 -3 26 103
use INVX2  INVX2_37
timestamp 1693479267
transform 1 0 2076 0 -1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_239
timestamp 1693479267
transform -1 0 2116 0 -1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_97
timestamp 1693479267
transform -1 0 2140 0 -1 305
box -2 -3 26 103
use INVX2  INVX2_36
timestamp 1693479267
transform 1 0 2140 0 -1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_536
timestamp 1693479267
transform -1 0 2180 0 -1 305
box -2 -3 26 103
use NAND3X1  NAND3X1_99
timestamp 1693479267
transform 1 0 2180 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_530
timestamp 1693479267
transform 1 0 2212 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_491
timestamp 1693479267
transform 1 0 2236 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_98
timestamp 1693479267
transform 1 0 2268 0 -1 305
box -2 -3 34 103
use AND2X2  AND2X2_35
timestamp 1693479267
transform -1 0 2332 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_233
timestamp 1693479267
transform 1 0 2332 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_493
timestamp 1693479267
transform 1 0 2356 0 -1 305
box -2 -3 34 103
use OAI22X1  OAI22X1_11
timestamp 1693479267
transform 1 0 2388 0 -1 305
box -2 -3 42 103
use OAI21X1  OAI21X1_487
timestamp 1693479267
transform 1 0 2428 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_147
timestamp 1693479267
transform 1 0 2460 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_548
timestamp 1693479267
transform 1 0 2484 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_91
timestamp 1693479267
transform 1 0 2516 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_4_0
timestamp 1693479267
transform 1 0 2548 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_4_1
timestamp 1693479267
transform 1 0 2556 0 -1 305
box -2 -3 10 103
use INVX2  INVX2_53
timestamp 1693479267
transform 1 0 2564 0 -1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_474
timestamp 1693479267
transform 1 0 2580 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_512
timestamp 1693479267
transform -1 0 2636 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_41
timestamp 1693479267
transform 1 0 2636 0 -1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_91
timestamp 1693479267
transform -1 0 2700 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_326
timestamp 1693479267
transform 1 0 2700 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_383
timestamp 1693479267
transform 1 0 2732 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_93
timestamp 1693479267
transform -1 0 2788 0 -1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_30
timestamp 1693479267
transform 1 0 2788 0 -1 305
box -2 -3 50 103
use NAND2X1  NAND2X1_380
timestamp 1693479267
transform -1 0 2860 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_430
timestamp 1693479267
transform -1 0 2892 0 -1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_22
timestamp 1693479267
transform 1 0 2892 0 -1 305
box -2 -3 50 103
use NAND2X1  NAND2X1_326
timestamp 1693479267
transform 1 0 2940 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_405
timestamp 1693479267
transform -1 0 2988 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_340
timestamp 1693479267
transform 1 0 2988 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_454
timestamp 1693479267
transform -1 0 3036 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_401
timestamp 1693479267
transform 1 0 3036 0 -1 305
box -2 -3 26 103
use FILL  FILL_2_5_0
timestamp 1693479267
transform -1 0 3068 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_5_1
timestamp 1693479267
transform -1 0 3076 0 -1 305
box -2 -3 10 103
use NAND2X1  NAND2X1_455
timestamp 1693479267
transform -1 0 3100 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_471
timestamp 1693479267
transform -1 0 3124 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_341
timestamp 1693479267
transform -1 0 3148 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_415
timestamp 1693479267
transform -1 0 3180 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_352
timestamp 1693479267
transform 1 0 3180 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_431
timestamp 1693479267
transform -1 0 3244 0 -1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_33
timestamp 1693479267
transform 1 0 3244 0 -1 305
box -2 -3 50 103
use NAND2X1  NAND2X1_417
timestamp 1693479267
transform -1 0 3316 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_388
timestamp 1693479267
transform -1 0 3340 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_401
timestamp 1693479267
transform 1 0 3340 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_367
timestamp 1693479267
transform -1 0 3388 0 -1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_503
timestamp 1693479267
transform 1 0 3388 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_490
timestamp 1693479267
transform 1 0 3412 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_531
timestamp 1693479267
transform -1 0 3468 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_464
timestamp 1693479267
transform 1 0 3468 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_518
timestamp 1693479267
transform 1 0 3492 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_350
timestamp 1693479267
transform -1 0 3556 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_478
timestamp 1693479267
transform 1 0 3556 0 -1 305
box -2 -3 26 103
use FILL  FILL_2_6_0
timestamp 1693479267
transform 1 0 3580 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_6_1
timestamp 1693479267
transform 1 0 3588 0 -1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_400
timestamp 1693479267
transform 1 0 3596 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_517
timestamp 1693479267
transform -1 0 3660 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_496
timestamp 1693479267
transform -1 0 3684 0 -1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_191
timestamp 1693479267
transform 1 0 3684 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_608
timestamp 1693479267
transform -1 0 3740 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_116
timestamp 1693479267
transform -1 0 3764 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_561
timestamp 1693479267
transform 1 0 3764 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_563
timestamp 1693479267
transform 1 0 3796 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_117
timestamp 1693479267
transform 1 0 3828 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_564
timestamp 1693479267
transform -1 0 3892 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_281
timestamp 1693479267
transform 1 0 3892 0 -1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_282
timestamp 1693479267
transform -1 0 3940 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_562
timestamp 1693479267
transform 1 0 3940 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_500
timestamp 1693479267
transform -1 0 3996 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_571
timestamp 1693479267
transform 1 0 3996 0 -1 305
box -2 -3 34 103
use OAI22X1  OAI22X1_8
timestamp 1693479267
transform 1 0 4028 0 -1 305
box -2 -3 42 103
use FILL  FILL_2_7_0
timestamp 1693479267
transform 1 0 4068 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_7_1
timestamp 1693479267
transform 1 0 4076 0 -1 305
box -2 -3 10 103
use OAI22X1  OAI22X1_29
timestamp 1693479267
transform 1 0 4084 0 -1 305
box -2 -3 42 103
use AOI21X1  AOI21X1_129
timestamp 1693479267
transform 1 0 4124 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_593
timestamp 1693479267
transform 1 0 4156 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_119
timestamp 1693479267
transform -1 0 4220 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_573
timestamp 1693479267
transform 1 0 4220 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_602
timestamp 1693479267
transform 1 0 4252 0 -1 305
box -2 -3 34 103
use INVX2  INVX2_64
timestamp 1693479267
transform -1 0 4300 0 -1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_525
timestamp 1693479267
transform -1 0 4324 0 -1 305
box -2 -3 26 103
use AOI22X1  AOI22X1_99
timestamp 1693479267
transform 1 0 4324 0 -1 305
box -2 -3 42 103
use NAND2X1  NAND2X1_519
timestamp 1693479267
transform 1 0 4364 0 -1 305
box -2 -3 26 103
use NAND3X1  NAND3X1_138
timestamp 1693479267
transform 1 0 4388 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_581
timestamp 1693479267
transform -1 0 4452 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_293
timestamp 1693479267
transform 1 0 4452 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_123
timestamp 1693479267
transform 1 0 4476 0 -1 305
box -2 -3 34 103
use OAI22X1  OAI22X1_32
timestamp 1693479267
transform -1 0 4548 0 -1 305
box -2 -3 42 103
use BUFX4  BUFX4_115
timestamp 1693479267
transform 1 0 4548 0 -1 305
box -2 -3 34 103
use FILL  FILL_3_1
timestamp 1693479267
transform -1 0 4588 0 -1 305
box -2 -3 10 103
use FILL  FILL_3_2
timestamp 1693479267
transform -1 0 4596 0 -1 305
box -2 -3 10 103
use FILL  FILL_3_3
timestamp 1693479267
transform -1 0 4604 0 -1 305
box -2 -3 10 103
use NAND2X1  NAND2X1_656
timestamp 1693479267
transform 1 0 4 0 1 305
box -2 -3 26 103
use INVX1  INVX1_474
timestamp 1693479267
transform 1 0 28 0 1 305
box -2 -3 18 103
use INVX1  INVX1_475
timestamp 1693479267
transform 1 0 44 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_830
timestamp 1693479267
transform -1 0 92 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_828
timestamp 1693479267
transform 1 0 92 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_654
timestamp 1693479267
transform -1 0 148 0 1 305
box -2 -3 26 103
use INVX1  INVX1_473
timestamp 1693479267
transform -1 0 164 0 1 305
box -2 -3 18 103
use OR2X2  OR2X2_46
timestamp 1693479267
transform 1 0 164 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_386
timestamp 1693479267
transform -1 0 220 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_831
timestamp 1693479267
transform -1 0 252 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_832
timestamp 1693479267
transform 1 0 252 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_183
timestamp 1693479267
transform -1 0 316 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_168
timestamp 1693479267
transform 1 0 316 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_21
timestamp 1693479267
transform -1 0 380 0 1 305
box -2 -3 34 103
use NOR3X1  NOR3X1_65
timestamp 1693479267
transform 1 0 380 0 1 305
box -2 -3 66 103
use NOR2X1  NOR2X1_384
timestamp 1693479267
transform 1 0 444 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_825
timestamp 1693479267
transform -1 0 500 0 1 305
box -2 -3 34 103
use FILL  FILL_3_0_0
timestamp 1693479267
transform -1 0 508 0 1 305
box -2 -3 10 103
use FILL  FILL_3_0_1
timestamp 1693479267
transform -1 0 516 0 1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_824
timestamp 1693479267
transform -1 0 548 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_382
timestamp 1693479267
transform -1 0 572 0 1 305
box -2 -3 26 103
use NAND3X1  NAND3X1_180
timestamp 1693479267
transform -1 0 604 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_447
timestamp 1693479267
transform -1 0 700 0 1 305
box -2 -3 98 103
use INVX1  INVX1_471
timestamp 1693479267
transform 1 0 700 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_820
timestamp 1693479267
transform 1 0 716 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_648
timestamp 1693479267
transform -1 0 772 0 1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_651
timestamp 1693479267
transform 1 0 772 0 1 305
box -2 -3 26 103
use CLKBUF1  CLKBUF1_33
timestamp 1693479267
transform -1 0 868 0 1 305
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_477
timestamp 1693479267
transform -1 0 964 0 1 305
box -2 -3 98 103
use FILL  FILL_3_1_0
timestamp 1693479267
transform 1 0 964 0 1 305
box -2 -3 10 103
use FILL  FILL_3_1_1
timestamp 1693479267
transform 1 0 972 0 1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_166
timestamp 1693479267
transform 1 0 980 0 1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_261
timestamp 1693479267
transform 1 0 1076 0 1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_165
timestamp 1693479267
transform 1 0 1172 0 1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_162
timestamp 1693479267
transform 1 0 1268 0 1 305
box -2 -3 98 103
use XNOR2X1  XNOR2X1_32
timestamp 1693479267
transform 1 0 1364 0 1 305
box -2 -3 58 103
use NOR2X1  NOR2X1_47
timestamp 1693479267
transform 1 0 1420 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_21
timestamp 1693479267
transform 1 0 1444 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_149
timestamp 1693479267
transform -1 0 1500 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_22
timestamp 1693479267
transform 1 0 1500 0 1 305
box -2 -3 34 103
use FILL  FILL_3_2_0
timestamp 1693479267
transform 1 0 1532 0 1 305
box -2 -3 10 103
use FILL  FILL_3_2_1
timestamp 1693479267
transform 1 0 1540 0 1 305
box -2 -3 10 103
use INVX2  INVX2_12
timestamp 1693479267
transform 1 0 1548 0 1 305
box -2 -3 18 103
use NOR2X1  NOR2X1_37
timestamp 1693479267
transform 1 0 1564 0 1 305
box -2 -3 26 103
use XNOR2X1  XNOR2X1_31
timestamp 1693479267
transform -1 0 1644 0 1 305
box -2 -3 58 103
use XNOR2X1  XNOR2X1_33
timestamp 1693479267
transform -1 0 1700 0 1 305
box -2 -3 58 103
use NAND2X1  NAND2X1_261
timestamp 1693479267
transform 1 0 1700 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_314
timestamp 1693479267
transform 1 0 1724 0 1 305
box -2 -3 34 103
use INVX1  INVX1_326
timestamp 1693479267
transform 1 0 1756 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_696
timestamp 1693479267
transform -1 0 1804 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_302
timestamp 1693479267
transform -1 0 1836 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_609
timestamp 1693479267
transform 1 0 1836 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_148
timestamp 1693479267
transform -1 0 1900 0 1 305
box -2 -3 34 103
use INVX1  INVX1_401
timestamp 1693479267
transform -1 0 1916 0 1 305
box -2 -3 18 103
use INVX2  INVX2_67
timestamp 1693479267
transform 1 0 1916 0 1 305
box -2 -3 18 103
use INVX2  INVX2_68
timestamp 1693479267
transform -1 0 1948 0 1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_238
timestamp 1693479267
transform 1 0 1948 0 1 305
box -2 -3 26 103
use AOI22X1  AOI22X1_101
timestamp 1693479267
transform 1 0 1972 0 1 305
box -2 -3 42 103
use OAI21X1  OAI21X1_641
timestamp 1693479267
transform -1 0 2044 0 1 305
box -2 -3 34 103
use FILL  FILL_3_3_0
timestamp 1693479267
transform -1 0 2052 0 1 305
box -2 -3 10 103
use FILL  FILL_3_3_1
timestamp 1693479267
transform -1 0 2060 0 1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_617
timestamp 1693479267
transform -1 0 2092 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_103
timestamp 1693479267
transform -1 0 2116 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_494
timestamp 1693479267
transform -1 0 2148 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_117
timestamp 1693479267
transform 1 0 2148 0 1 305
box -2 -3 34 103
use AOI22X1  AOI22X1_85
timestamp 1693479267
transform -1 0 2220 0 1 305
box -2 -3 42 103
use NOR2X1  NOR2X1_232
timestamp 1693479267
transform 1 0 2220 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_492
timestamp 1693479267
transform -1 0 2276 0 1 305
box -2 -3 34 103
use AOI22X1  AOI22X1_86
timestamp 1693479267
transform 1 0 2276 0 1 305
box -2 -3 42 103
use INVX2  INVX2_57
timestamp 1693479267
transform 1 0 2316 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_500
timestamp 1693479267
transform -1 0 2364 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_228
timestamp 1693479267
transform 1 0 2364 0 1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_460
timestamp 1693479267
transform -1 0 2412 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_490
timestamp 1693479267
transform 1 0 2412 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_486
timestamp 1693479267
transform -1 0 2476 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_501
timestamp 1693479267
transform 1 0 2476 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_470
timestamp 1693479267
transform -1 0 2532 0 1 305
box -2 -3 26 103
use FILL  FILL_3_4_0
timestamp 1693479267
transform 1 0 2532 0 1 305
box -2 -3 10 103
use FILL  FILL_3_4_1
timestamp 1693479267
transform 1 0 2540 0 1 305
box -2 -3 10 103
use AOI22X1  AOI22X1_88
timestamp 1693479267
transform 1 0 2548 0 1 305
box -2 -3 42 103
use OAI21X1  OAI21X1_325
timestamp 1693479267
transform -1 0 2620 0 1 305
box -2 -3 34 103
use INVX2  INVX2_47
timestamp 1693479267
transform -1 0 2636 0 1 305
box -2 -3 18 103
use NOR2X1  NOR2X1_152
timestamp 1693479267
transform 1 0 2636 0 1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_296
timestamp 1693479267
transform -1 0 2684 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_503
timestamp 1693479267
transform 1 0 2684 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_112
timestamp 1693479267
transform -1 0 2748 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_469
timestamp 1693479267
transform -1 0 2780 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_43
timestamp 1693479267
transform 1 0 2780 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_146
timestamp 1693479267
transform 1 0 2812 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_394
timestamp 1693479267
transform -1 0 2876 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_398
timestamp 1693479267
transform 1 0 2876 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_384
timestamp 1693479267
transform -1 0 2932 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_419
timestamp 1693479267
transform 1 0 2932 0 1 305
box -2 -3 34 103
use INVX1  INVX1_386
timestamp 1693479267
transform 1 0 2964 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_505
timestamp 1693479267
transform 1 0 2980 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_481
timestamp 1693479267
transform -1 0 3044 0 1 305
box -2 -3 34 103
use FILL  FILL_3_5_0
timestamp 1693479267
transform -1 0 3052 0 1 305
box -2 -3 10 103
use FILL  FILL_3_5_1
timestamp 1693479267
transform -1 0 3060 0 1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_416
timestamp 1693479267
transform -1 0 3092 0 1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_27
timestamp 1693479267
transform 1 0 3092 0 1 305
box -2 -3 50 103
use MUX2X1  MUX2X1_41
timestamp 1693479267
transform 1 0 3140 0 1 305
box -2 -3 50 103
use NAND2X1  NAND2X1_331
timestamp 1693479267
transform -1 0 3212 0 1 305
box -2 -3 26 103
use BUFX4  BUFX4_227
timestamp 1693479267
transform -1 0 3244 0 1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_39
timestamp 1693479267
transform 1 0 3244 0 1 305
box -2 -3 50 103
use OAI21X1  OAI21X1_404
timestamp 1693479267
transform 1 0 3292 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_389
timestamp 1693479267
transform -1 0 3348 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_405
timestamp 1693479267
transform -1 0 3380 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_537
timestamp 1693479267
transform 1 0 3380 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_532
timestamp 1693479267
transform 1 0 3404 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_612
timestamp 1693479267
transform -1 0 3468 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_229
timestamp 1693479267
transform -1 0 3500 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_333
timestamp 1693479267
transform 1 0 3500 0 1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_332
timestamp 1693479267
transform -1 0 3548 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_108
timestamp 1693479267
transform 1 0 3548 0 1 305
box -2 -3 34 103
use FILL  FILL_3_6_0
timestamp 1693479267
transform 1 0 3580 0 1 305
box -2 -3 10 103
use FILL  FILL_3_6_1
timestamp 1693479267
transform 1 0 3588 0 1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_542
timestamp 1693479267
transform 1 0 3596 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_385
timestamp 1693479267
transform -1 0 3652 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_594
timestamp 1693479267
transform -1 0 3684 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_108
timestamp 1693479267
transform 1 0 3684 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_551
timestamp 1693479267
transform 1 0 3708 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_552
timestamp 1693479267
transform -1 0 3772 0 1 305
box -2 -3 34 103
use OR2X2  OR2X2_32
timestamp 1693479267
transform 1 0 3772 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_132
timestamp 1693479267
transform 1 0 3804 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_565
timestamp 1693479267
transform -1 0 3868 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_275
timestamp 1693479267
transform 1 0 3868 0 1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_276
timestamp 1693479267
transform -1 0 3916 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_555
timestamp 1693479267
transform -1 0 3948 0 1 305
box -2 -3 34 103
use INVX2  INVX2_61
timestamp 1693479267
transform -1 0 3964 0 1 305
box -2 -3 18 103
use AOI22X1  AOI22X1_97
timestamp 1693479267
transform 1 0 3964 0 1 305
box -2 -3 42 103
use NAND2X1  NAND2X1_308
timestamp 1693479267
transform -1 0 4028 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_560
timestamp 1693479267
transform 1 0 4028 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_134
timestamp 1693479267
transform 1 0 4060 0 1 305
box -2 -3 34 103
use FILL  FILL_3_7_0
timestamp 1693479267
transform 1 0 4092 0 1 305
box -2 -3 10 103
use FILL  FILL_3_7_1
timestamp 1693479267
transform 1 0 4100 0 1 305
box -2 -3 10 103
use NAND3X1  NAND3X1_140
timestamp 1693479267
transform 1 0 4108 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_119
timestamp 1693479267
transform -1 0 4164 0 1 305
box -2 -3 26 103
use OAI22X1  OAI22X1_36
timestamp 1693479267
transform 1 0 4164 0 1 305
box -2 -3 42 103
use AOI21X1  AOI21X1_127
timestamp 1693479267
transform -1 0 4236 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_144
timestamp 1693479267
transform 1 0 4236 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_304
timestamp 1693479267
transform 1 0 4268 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_125
timestamp 1693479267
transform -1 0 4324 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_582
timestamp 1693479267
transform -1 0 4356 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_294
timestamp 1693479267
transform 1 0 4356 0 1 305
box -2 -3 26 103
use AND2X2  AND2X2_47
timestamp 1693479267
transform 1 0 4380 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_574
timestamp 1693479267
transform 1 0 4412 0 1 305
box -2 -3 34 103
use OR2X2  OR2X2_34
timestamp 1693479267
transform 1 0 4444 0 1 305
box -2 -3 34 103
use INVX2  INVX2_63
timestamp 1693479267
transform 1 0 4476 0 1 305
box -2 -3 18 103
use NOR2X1  NOR2X1_286
timestamp 1693479267
transform 1 0 4492 0 1 305
box -2 -3 26 103
use AND2X2  AND2X2_46
timestamp 1693479267
transform -1 0 4548 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_572
timestamp 1693479267
transform 1 0 4548 0 1 305
box -2 -3 34 103
use FILL  FILL_4_1
timestamp 1693479267
transform 1 0 4580 0 1 305
box -2 -3 10 103
use FILL  FILL_4_2
timestamp 1693479267
transform 1 0 4588 0 1 305
box -2 -3 10 103
use FILL  FILL_4_3
timestamp 1693479267
transform 1 0 4596 0 1 305
box -2 -3 10 103
use BUFX2  BUFX2_50
timestamp 1693479267
transform -1 0 28 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_451
timestamp 1693479267
transform 1 0 28 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_483
timestamp 1693479267
transform -1 0 220 0 -1 505
box -2 -3 98 103
use NAND3X1  NAND3X1_29
timestamp 1693479267
transform 1 0 220 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_172
timestamp 1693479267
transform -1 0 284 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_28
timestamp 1693479267
transform 1 0 284 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_75
timestamp 1693479267
transform -1 0 348 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_20
timestamp 1693479267
transform -1 0 380 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_479
timestamp 1693479267
transform 1 0 380 0 -1 505
box -2 -3 98 103
use INVX1  INVX1_472
timestamp 1693479267
transform 1 0 476 0 -1 505
box -2 -3 18 103
use FILL  FILL_4_0_0
timestamp 1693479267
transform -1 0 500 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_0_1
timestamp 1693479267
transform -1 0 508 0 -1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_823
timestamp 1693479267
transform -1 0 540 0 -1 505
box -2 -3 34 103
use INVX2  INVX2_72
timestamp 1693479267
transform -1 0 556 0 -1 505
box -2 -3 18 103
use AND2X2  AND2X2_77
timestamp 1693479267
transform 1 0 556 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_181
timestamp 1693479267
transform -1 0 620 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_645
timestamp 1693479267
transform -1 0 644 0 -1 505
box -2 -3 26 103
use AND2X2  AND2X2_76
timestamp 1693479267
transform -1 0 676 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_179
timestamp 1693479267
transform -1 0 708 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_643
timestamp 1693479267
transform -1 0 732 0 -1 505
box -2 -3 26 103
use INVX1  INVX1_470
timestamp 1693479267
transform 1 0 732 0 -1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_821
timestamp 1693479267
transform 1 0 748 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_476
timestamp 1693479267
transform -1 0 876 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_166
timestamp 1693479267
transform -1 0 908 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_17
timestamp 1693479267
transform -1 0 940 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_16
timestamp 1693479267
transform -1 0 972 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_1_0
timestamp 1693479267
transform 1 0 972 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_1_1
timestamp 1693479267
transform 1 0 980 0 -1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_445
timestamp 1693479267
transform 1 0 988 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_259
timestamp 1693479267
transform 1 0 1084 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_265
timestamp 1693479267
transform 1 0 1180 0 -1 505
box -2 -3 98 103
use XNOR2X1  XNOR2X1_29
timestamp 1693479267
transform 1 0 1276 0 -1 505
box -2 -3 58 103
use XNOR2X1  XNOR2X1_30
timestamp 1693479267
transform 1 0 1332 0 -1 505
box -2 -3 58 103
use OAI21X1  OAI21X1_252
timestamp 1693479267
transform 1 0 1388 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_176
timestamp 1693479267
transform 1 0 1420 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_249
timestamp 1693479267
transform -1 0 1476 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_253
timestamp 1693479267
transform 1 0 1476 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_46
timestamp 1693479267
transform -1 0 1532 0 -1 505
box -2 -3 26 103
use FILL  FILL_4_2_0
timestamp 1693479267
transform -1 0 1540 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_2_1
timestamp 1693479267
transform -1 0 1548 0 -1 505
box -2 -3 10 103
use XNOR2X1  XNOR2X1_43
timestamp 1693479267
transform -1 0 1604 0 -1 505
box -2 -3 58 103
use AOI22X1  AOI22X1_48
timestamp 1693479267
transform 1 0 1604 0 -1 505
box -2 -3 42 103
use AOI22X1  AOI22X1_47
timestamp 1693479267
transform -1 0 1684 0 -1 505
box -2 -3 42 103
use OAI21X1  OAI21X1_299
timestamp 1693479267
transform 1 0 1684 0 -1 505
box -2 -3 34 103
use INVX1  INVX1_337
timestamp 1693479267
transform 1 0 1716 0 -1 505
box -2 -3 18 103
use MUX2X1  MUX2X1_10
timestamp 1693479267
transform -1 0 1780 0 -1 505
box -2 -3 50 103
use INVX1  INVX1_345
timestamp 1693479267
transform 1 0 1780 0 -1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_610
timestamp 1693479267
transform -1 0 1828 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_309
timestamp 1693479267
transform -1 0 1852 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_611
timestamp 1693479267
transform -1 0 1884 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_605
timestamp 1693479267
transform 1 0 1884 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_307
timestamp 1693479267
transform 1 0 1916 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_604
timestamp 1693479267
transform 1 0 1940 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_535
timestamp 1693479267
transform -1 0 1996 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_600
timestamp 1693479267
transform -1 0 2028 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_3_0
timestamp 1693479267
transform 1 0 2028 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_3_1
timestamp 1693479267
transform 1 0 2036 0 -1 505
box -2 -3 10 103
use NAND2X1  NAND2X1_531
timestamp 1693479267
transform 1 0 2044 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_450
timestamp 1693479267
transform 1 0 2068 0 -1 505
box -2 -3 26 103
use INVX1  INVX1_344
timestamp 1693479267
transform 1 0 2092 0 -1 505
box -2 -3 18 103
use INVX1  INVX1_399
timestamp 1693479267
transform -1 0 2124 0 -1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_322
timestamp 1693479267
transform 1 0 2124 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_283
timestamp 1693479267
transform -1 0 2180 0 -1 505
box -2 -3 26 103
use INVX1  INVX1_380
timestamp 1693479267
transform 1 0 2180 0 -1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_451
timestamp 1693479267
transform -1 0 2220 0 -1 505
box -2 -3 26 103
use OAI22X1  OAI22X1_18
timestamp 1693479267
transform -1 0 2260 0 -1 505
box -2 -3 42 103
use OAI21X1  OAI21X1_515
timestamp 1693479267
transform 1 0 2260 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_87
timestamp 1693479267
transform -1 0 2324 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_479
timestamp 1693479267
transform -1 0 2356 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_224
timestamp 1693479267
transform -1 0 2380 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_221
timestamp 1693479267
transform -1 0 2404 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_88
timestamp 1693479267
transform -1 0 2436 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_295
timestamp 1693479267
transform -1 0 2460 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_149
timestamp 1693479267
transform -1 0 2484 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_81
timestamp 1693479267
transform -1 0 2516 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_468
timestamp 1693479267
transform -1 0 2548 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_4_0
timestamp 1693479267
transform -1 0 2556 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_4_1
timestamp 1693479267
transform -1 0 2564 0 -1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_467
timestamp 1693479267
transform -1 0 2596 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_510
timestamp 1693479267
transform 1 0 2596 0 -1 505
box -2 -3 34 103
use OAI22X1  OAI22X1_12
timestamp 1693479267
transform -1 0 2668 0 -1 505
box -2 -3 42 103
use AOI21X1  AOI21X1_86
timestamp 1693479267
transform -1 0 2700 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_148
timestamp 1693479267
transform 1 0 2700 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_284
timestamp 1693479267
transform 1 0 2724 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_339
timestamp 1693479267
transform -1 0 2780 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_153
timestamp 1693479267
transform 1 0 2780 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_285
timestamp 1693479267
transform -1 0 2828 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_286
timestamp 1693479267
transform -1 0 2852 0 -1 505
box -2 -3 26 103
use OAI22X1  OAI22X1_15
timestamp 1693479267
transform -1 0 2892 0 -1 505
box -2 -3 42 103
use AOI21X1  AOI21X1_82
timestamp 1693479267
transform -1 0 2924 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_417
timestamp 1693479267
transform -1 0 2956 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_345
timestamp 1693479267
transform -1 0 2988 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_327
timestamp 1693479267
transform -1 0 3012 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_457
timestamp 1693479267
transform -1 0 3036 0 -1 505
box -2 -3 26 103
use INVX1  INVX1_375
timestamp 1693479267
transform 1 0 3036 0 -1 505
box -2 -3 18 103
use FILL  FILL_4_5_0
timestamp 1693479267
transform -1 0 3060 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_5_1
timestamp 1693479267
transform -1 0 3068 0 -1 505
box -2 -3 10 103
use NOR2X1  NOR2X1_225
timestamp 1693479267
transform -1 0 3092 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_435
timestamp 1693479267
transform 1 0 3092 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_451
timestamp 1693479267
transform 1 0 3124 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_429
timestamp 1693479267
transform -1 0 3180 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_353
timestamp 1693479267
transform -1 0 3212 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_427
timestamp 1693479267
transform -1 0 3236 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_67
timestamp 1693479267
transform -1 0 3268 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_548
timestamp 1693479267
transform -1 0 3292 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_434
timestamp 1693479267
transform -1 0 3324 0 -1 505
box -2 -3 34 103
use MUX2X1  MUX2X1_23
timestamp 1693479267
transform 1 0 3324 0 -1 505
box -2 -3 50 103
use NAND2X1  NAND2X1_502
timestamp 1693479267
transform -1 0 3396 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_556
timestamp 1693479267
transform -1 0 3428 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_226
timestamp 1693479267
transform -1 0 3460 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_495
timestamp 1693479267
transform 1 0 3460 0 -1 505
box -2 -3 34 103
use MUX2X1  MUX2X1_8
timestamp 1693479267
transform 1 0 3492 0 -1 505
box -2 -3 50 103
use NAND2X1  NAND2X1_255
timestamp 1693479267
transform -1 0 3564 0 -1 505
box -2 -3 26 103
use FILL  FILL_4_6_0
timestamp 1693479267
transform -1 0 3572 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_6_1
timestamp 1693479267
transform -1 0 3580 0 -1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_312
timestamp 1693479267
transform -1 0 3612 0 -1 505
box -2 -3 34 103
use INVX1  INVX1_335
timestamp 1693479267
transform -1 0 3628 0 -1 505
box -2 -3 18 103
use MUX2X1  MUX2X1_35
timestamp 1693479267
transform -1 0 3676 0 -1 505
box -2 -3 50 103
use NAND2X1  NAND2X1_258
timestamp 1693479267
transform 1 0 3676 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_313
timestamp 1693479267
transform -1 0 3732 0 -1 505
box -2 -3 34 103
use INVX1  INVX1_336
timestamp 1693479267
transform -1 0 3748 0 -1 505
box -2 -3 18 103
use MUX2X1  MUX2X1_9
timestamp 1693479267
transform 1 0 3748 0 -1 505
box -2 -3 50 103
use NOR2X1  NOR2X1_171
timestamp 1693479267
transform -1 0 3820 0 -1 505
box -2 -3 26 103
use NAND3X1  NAND3X1_98
timestamp 1693479267
transform 1 0 3820 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_167
timestamp 1693479267
transform -1 0 3876 0 -1 505
box -2 -3 26 103
use INVX2  INVX2_42
timestamp 1693479267
transform -1 0 3892 0 -1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_299
timestamp 1693479267
transform -1 0 3916 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_264
timestamp 1693479267
transform 1 0 3916 0 -1 505
box -2 -3 26 103
use NAND3X1  NAND3X1_93
timestamp 1693479267
transform 1 0 3940 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_253
timestamp 1693479267
transform -1 0 3996 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_298
timestamp 1693479267
transform -1 0 4020 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_329
timestamp 1693479267
transform -1 0 4052 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_130
timestamp 1693479267
transform -1 0 4084 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_7_0
timestamp 1693479267
transform 1 0 4084 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_7_1
timestamp 1693479267
transform 1 0 4092 0 -1 505
box -2 -3 10 103
use NOR2X1  NOR2X1_296
timestamp 1693479267
transform 1 0 4100 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_590
timestamp 1693479267
transform -1 0 4156 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_554
timestamp 1693479267
transform -1 0 4188 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_603
timestamp 1693479267
transform 1 0 4188 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_601
timestamp 1693479267
transform -1 0 4252 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_534
timestamp 1693479267
transform -1 0 4276 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_242
timestamp 1693479267
transform -1 0 4300 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_262
timestamp 1693479267
transform 1 0 4300 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_168
timestamp 1693479267
transform -1 0 4348 0 -1 505
box -2 -3 26 103
use INVX2  INVX2_45
timestamp 1693479267
transform 1 0 4348 0 -1 505
box -2 -3 18 103
use NOR2X1  NOR2X1_125
timestamp 1693479267
transform -1 0 4388 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_480
timestamp 1693479267
transform -1 0 4412 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_263
timestamp 1693479267
transform 1 0 4412 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_485
timestamp 1693479267
transform -1 0 4460 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_305
timestamp 1693479267
transform 1 0 4460 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_141
timestamp 1693479267
transform 1 0 4484 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_260
timestamp 1693479267
transform -1 0 4540 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_297
timestamp 1693479267
transform -1 0 4564 0 -1 505
box -2 -3 26 103
use INVX2  INVX2_44
timestamp 1693479267
transform -1 0 4580 0 -1 505
box -2 -3 18 103
use FILL  FILL_5_1
timestamp 1693479267
transform -1 0 4588 0 -1 505
box -2 -3 10 103
use FILL  FILL_5_2
timestamp 1693479267
transform -1 0 4596 0 -1 505
box -2 -3 10 103
use FILL  FILL_5_3
timestamp 1693479267
transform -1 0 4604 0 -1 505
box -2 -3 10 103
use BUFX2  BUFX2_56
timestamp 1693479267
transform -1 0 28 0 1 505
box -2 -3 26 103
use BUFX2  BUFX2_12
timestamp 1693479267
transform -1 0 52 0 1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_169
timestamp 1693479267
transform -1 0 148 0 1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_457
timestamp 1693479267
transform 1 0 148 0 1 505
box -2 -3 98 103
use NAND3X1  NAND3X1_40
timestamp 1693479267
transform 1 0 244 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_657
timestamp 1693479267
transform -1 0 300 0 1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_271
timestamp 1693479267
transform 1 0 300 0 1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_478
timestamp 1693479267
transform 1 0 396 0 1 505
box -2 -3 98 103
use FILL  FILL_5_0_0
timestamp 1693479267
transform -1 0 500 0 1 505
box -2 -3 10 103
use FILL  FILL_5_0_1
timestamp 1693479267
transform -1 0 508 0 1 505
box -2 -3 10 103
use XNOR2X1  XNOR2X1_50
timestamp 1693479267
transform -1 0 564 0 1 505
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_446
timestamp 1693479267
transform 1 0 564 0 1 505
box -2 -3 98 103
use AND2X2  AND2X2_75
timestamp 1693479267
transform -1 0 692 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_381
timestamp 1693479267
transform -1 0 716 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_819
timestamp 1693479267
transform 1 0 716 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_15
timestamp 1693479267
transform 1 0 748 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_165
timestamp 1693479267
transform -1 0 812 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_74
timestamp 1693479267
transform 1 0 812 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_15
timestamp 1693479267
transform -1 0 876 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_14
timestamp 1693479267
transform -1 0 908 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_444
timestamp 1693479267
transform 1 0 908 0 1 505
box -2 -3 98 103
use FILL  FILL_5_1_0
timestamp 1693479267
transform 1 0 1004 0 1 505
box -2 -3 10 103
use FILL  FILL_5_1_1
timestamp 1693479267
transform 1 0 1012 0 1 505
box -2 -3 10 103
use BUFX2  BUFX2_20
timestamp 1693479267
transform 1 0 1020 0 1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_260
timestamp 1693479267
transform 1 0 1044 0 1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_644
timestamp 1693479267
transform 1 0 1140 0 1 505
box -2 -3 26 103
use CLKBUF1  CLKBUF1_54
timestamp 1693479267
transform 1 0 1164 0 1 505
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_258
timestamp 1693479267
transform 1 0 1236 0 1 505
box -2 -3 98 103
use NOR2X1  NOR2X1_36
timestamp 1693479267
transform 1 0 1332 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_248
timestamp 1693479267
transform 1 0 1356 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_39
timestamp 1693479267
transform -1 0 1412 0 1 505
box -2 -3 26 103
use XNOR2X1  XNOR2X1_28
timestamp 1693479267
transform -1 0 1468 0 1 505
box -2 -3 58 103
use NAND3X1  NAND3X1_83
timestamp 1693479267
transform -1 0 1500 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_147
timestamp 1693479267
transform -1 0 1524 0 1 505
box -2 -3 26 103
use FILL  FILL_5_2_0
timestamp 1693479267
transform 1 0 1524 0 1 505
box -2 -3 10 103
use FILL  FILL_5_2_1
timestamp 1693479267
transform 1 0 1532 0 1 505
box -2 -3 10 103
use INVX1  INVX1_254
timestamp 1693479267
transform 1 0 1540 0 1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_148
timestamp 1693479267
transform 1 0 1556 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_251
timestamp 1693479267
transform -1 0 1612 0 1 505
box -2 -3 34 103
use INVX2  INVX2_11
timestamp 1693479267
transform -1 0 1628 0 1 505
box -2 -3 18 103
use INVX1  INVX1_257
timestamp 1693479267
transform -1 0 1644 0 1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_233
timestamp 1693479267
transform 1 0 1644 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_301
timestamp 1693479267
transform -1 0 1700 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_231
timestamp 1693479267
transform -1 0 1724 0 1 505
box -2 -3 26 103
use MUX2X1  MUX2X1_18
timestamp 1693479267
transform 1 0 1724 0 1 505
box -2 -3 50 103
use NAND2X1  NAND2X1_287
timestamp 1693479267
transform -1 0 1796 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_323
timestamp 1693479267
transform 1 0 1796 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_308
timestamp 1693479267
transform -1 0 1852 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_619
timestamp 1693479267
transform 1 0 1852 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_144
timestamp 1693479267
transform -1 0 1916 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_545
timestamp 1693479267
transform 1 0 1916 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_316
timestamp 1693479267
transform 1 0 1940 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_628
timestamp 1693479267
transform 1 0 1964 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_306
timestamp 1693479267
transform -1 0 2028 0 1 505
box -2 -3 34 103
use FILL  FILL_5_3_0
timestamp 1693479267
transform 1 0 2028 0 1 505
box -2 -3 10 103
use FILL  FILL_5_3_1
timestamp 1693479267
transform 1 0 2036 0 1 505
box -2 -3 10 103
use NOR2X1  NOR2X1_306
timestamp 1693479267
transform 1 0 2044 0 1 505
box -2 -3 26 103
use INVX1  INVX1_329
timestamp 1693479267
transform -1 0 2084 0 1 505
box -2 -3 18 103
use AOI22X1  AOI22X1_100
timestamp 1693479267
transform 1 0 2084 0 1 505
box -2 -3 42 103
use NAND3X1  NAND3X1_120
timestamp 1693479267
transform -1 0 2156 0 1 505
box -2 -3 34 103
use MUX2X1  MUX2X1_17
timestamp 1693479267
transform -1 0 2204 0 1 505
box -2 -3 50 103
use AOI21X1  AOI21X1_85
timestamp 1693479267
transform 1 0 2204 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_480
timestamp 1693479267
transform -1 0 2268 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_246
timestamp 1693479267
transform -1 0 2292 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_99
timestamp 1693479267
transform -1 0 2324 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_478
timestamp 1693479267
transform -1 0 2356 0 1 505
box -2 -3 34 103
use OAI22X1  OAI22X1_17
timestamp 1693479267
transform 1 0 2356 0 1 505
box -2 -3 42 103
use AND2X2  AND2X2_34
timestamp 1693479267
transform 1 0 2396 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_465
timestamp 1693479267
transform 1 0 2428 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_477
timestamp 1693479267
transform 1 0 2460 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_288
timestamp 1693479267
transform 1 0 2492 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_445
timestamp 1693479267
transform -1 0 2540 0 1 505
box -2 -3 26 103
use FILL  FILL_5_4_0
timestamp 1693479267
transform 1 0 2540 0 1 505
box -2 -3 10 103
use FILL  FILL_5_4_1
timestamp 1693479267
transform 1 0 2548 0 1 505
box -2 -3 10 103
use NOR2X1  NOR2X1_151
timestamp 1693479267
transform 1 0 2556 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_150
timestamp 1693479267
transform 1 0 2580 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_460
timestamp 1693479267
transform 1 0 2604 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_289
timestamp 1693479267
transform 1 0 2636 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_290
timestamp 1693479267
transform -1 0 2684 0 1 505
box -2 -3 26 103
use INVX1  INVX1_378
timestamp 1693479267
transform 1 0 2684 0 1 505
box -2 -3 18 103
use AOI22X1  AOI22X1_82
timestamp 1693479267
transform -1 0 2740 0 1 505
box -2 -3 42 103
use NAND2X1  NAND2X1_325
timestamp 1693479267
transform -1 0 2764 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_393
timestamp 1693479267
transform 1 0 2764 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_344
timestamp 1693479267
transform 1 0 2796 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_39
timestamp 1693479267
transform 1 0 2828 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_406
timestamp 1693479267
transform 1 0 2860 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_390
timestamp 1693479267
transform 1 0 2892 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_403
timestamp 1693479267
transform -1 0 2940 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_89
timestamp 1693479267
transform -1 0 2972 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_114
timestamp 1693479267
transform -1 0 3004 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_444
timestamp 1693479267
transform -1 0 3028 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_475
timestamp 1693479267
transform 1 0 3028 0 1 505
box -2 -3 34 103
use FILL  FILL_5_5_0
timestamp 1693479267
transform 1 0 3060 0 1 505
box -2 -3 10 103
use FILL  FILL_5_5_1
timestamp 1693479267
transform 1 0 3068 0 1 505
box -2 -3 10 103
use NAND2X1  NAND2X1_443
timestamp 1693479267
transform 1 0 3076 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_499
timestamp 1693479267
transform 1 0 3100 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_223
timestamp 1693479267
transform -1 0 3164 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_474
timestamp 1693479267
transform -1 0 3196 0 1 505
box -2 -3 34 103
use MUX2X1  MUX2X1_40
timestamp 1693479267
transform 1 0 3196 0 1 505
box -2 -3 50 103
use NAND2X1  NAND2X1_520
timestamp 1693479267
transform 1 0 3244 0 1 505
box -2 -3 26 103
use INVX1  INVX1_383
timestamp 1693479267
transform 1 0 3268 0 1 505
box -2 -3 18 103
use INVX1  INVX1_398
timestamp 1693479267
transform -1 0 3300 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_575
timestamp 1693479267
transform -1 0 3332 0 1 505
box -2 -3 34 103
use INVX1  INVX1_396
timestamp 1693479267
transform -1 0 3348 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_557
timestamp 1693479267
transform 1 0 3348 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_470
timestamp 1693479267
transform -1 0 3412 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_527
timestamp 1693479267
transform 1 0 3412 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_585
timestamp 1693479267
transform -1 0 3468 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_497
timestamp 1693479267
transform 1 0 3468 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_479
timestamp 1693479267
transform 1 0 3492 0 1 505
box -2 -3 26 103
use INVX1  INVX1_395
timestamp 1693479267
transform 1 0 3516 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_569
timestamp 1693479267
transform 1 0 3532 0 1 505
box -2 -3 34 103
use FILL  FILL_5_6_0
timestamp 1693479267
transform -1 0 3572 0 1 505
box -2 -3 10 103
use FILL  FILL_5_6_1
timestamp 1693479267
transform -1 0 3580 0 1 505
box -2 -3 10 103
use NAND2X1  NAND2X1_514
timestamp 1693479267
transform -1 0 3604 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_252
timestamp 1693479267
transform 1 0 3604 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_311
timestamp 1693479267
transform -1 0 3660 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_256
timestamp 1693479267
transform -1 0 3684 0 1 505
box -2 -3 26 103
use NAND3X1  NAND3X1_136
timestamp 1693479267
transform -1 0 3716 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_301
timestamp 1693479267
transform -1 0 3740 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_257
timestamp 1693479267
transform 1 0 3740 0 1 505
box -2 -3 26 103
use AOI22X1  AOI22X1_71
timestamp 1693479267
transform -1 0 3804 0 1 505
box -2 -3 42 103
use AOI21X1  AOI21X1_113
timestamp 1693479267
transform 1 0 3804 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_254
timestamp 1693479267
transform -1 0 3860 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_550
timestamp 1693479267
transform -1 0 3892 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_274
timestamp 1693479267
transform 1 0 3892 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_120
timestamp 1693479267
transform 1 0 3916 0 1 505
box -2 -3 26 103
use OAI22X1  OAI22X1_37
timestamp 1693479267
transform -1 0 3980 0 1 505
box -2 -3 42 103
use NOR2X1  NOR2X1_297
timestamp 1693479267
transform 1 0 3980 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_121
timestamp 1693479267
transform -1 0 4028 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_132
timestamp 1693479267
transform -1 0 4060 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_592
timestamp 1693479267
transform -1 0 4092 0 1 505
box -2 -3 34 103
use FILL  FILL_5_7_0
timestamp 1693479267
transform -1 0 4100 0 1 505
box -2 -3 10 103
use FILL  FILL_5_7_1
timestamp 1693479267
transform -1 0 4108 0 1 505
box -2 -3 10 103
use NOR2X1  NOR2X1_126
timestamp 1693479267
transform -1 0 4132 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_553
timestamp 1693479267
transform -1 0 4164 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_114
timestamp 1693479267
transform -1 0 4196 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_142
timestamp 1693479267
transform 1 0 4196 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_513
timestamp 1693479267
transform -1 0 4260 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_302
timestamp 1693479267
transform -1 0 4284 0 1 505
box -2 -3 26 103
use OAI22X1  OAI22X1_24
timestamp 1693479267
transform -1 0 4324 0 1 505
box -2 -3 42 103
use NOR2X1  NOR2X1_252
timestamp 1693479267
transform -1 0 4348 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_104
timestamp 1693479267
transform -1 0 4380 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_327
timestamp 1693479267
transform 1 0 4380 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_481
timestamp 1693479267
transform 1 0 4412 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_549
timestamp 1693479267
transform -1 0 4468 0 1 505
box -2 -3 34 103
use AOI22X1  AOI22X1_72
timestamp 1693479267
transform -1 0 4508 0 1 505
box -2 -3 42 103
use NOR2X1  NOR2X1_124
timestamp 1693479267
transform -1 0 4532 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_248
timestamp 1693479267
transform -1 0 4556 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_527
timestamp 1693479267
transform -1 0 4588 0 1 505
box -2 -3 34 103
use FILL  FILL_6_1
timestamp 1693479267
transform 1 0 4588 0 1 505
box -2 -3 10 103
use FILL  FILL_6_2
timestamp 1693479267
transform 1 0 4596 0 1 505
box -2 -3 10 103
use BUFX2  BUFX2_55
timestamp 1693479267
transform -1 0 28 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_489
timestamp 1693479267
transform -1 0 124 0 -1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_667
timestamp 1693479267
transform 1 0 124 0 -1 705
box -2 -3 26 103
use NAND3X1  NAND3X1_41
timestamp 1693479267
transform -1 0 180 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_178
timestamp 1693479267
transform -1 0 212 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_843
timestamp 1693479267
transform 1 0 212 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_14
timestamp 1693479267
transform -1 0 276 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_138
timestamp 1693479267
transform -1 0 308 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_72
timestamp 1693479267
transform -1 0 340 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_18
timestamp 1693479267
transform -1 0 372 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_19
timestamp 1693479267
transform -1 0 404 0 -1 705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_10
timestamp 1693479267
transform 1 0 404 0 -1 705
box -2 -3 74 103
use BUFX4  BUFX4_110
timestamp 1693479267
transform -1 0 508 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_0_0
timestamp 1693479267
transform -1 0 516 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_0_1
timestamp 1693479267
transform -1 0 524 0 -1 705
box -2 -3 10 103
use NAND3X1  NAND3X1_13
timestamp 1693479267
transform -1 0 556 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_475
timestamp 1693479267
transform 1 0 556 0 -1 705
box -2 -3 98 103
use NOR2X1  NOR2X1_380
timestamp 1693479267
transform 1 0 652 0 -1 705
box -2 -3 26 103
use BUFX4  BUFX4_111
timestamp 1693479267
transform 1 0 676 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_139
timestamp 1693479267
transform 1 0 708 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_12
timestamp 1693479267
transform -1 0 772 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_443
timestamp 1693479267
transform -1 0 868 0 -1 705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_257
timestamp 1693479267
transform 1 0 868 0 -1 705
box -2 -3 98 103
use XNOR2X1  XNOR2X1_25
timestamp 1693479267
transform 1 0 964 0 -1 705
box -2 -3 58 103
use FILL  FILL_6_1_0
timestamp 1693479267
transform 1 0 1020 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_1_1
timestamp 1693479267
transform 1 0 1028 0 -1 705
box -2 -3 10 103
use AOI21X1  AOI21X1_17
timestamp 1693479267
transform 1 0 1036 0 -1 705
box -2 -3 34 103
use XNOR2X1  XNOR2X1_22
timestamp 1693479267
transform 1 0 1068 0 -1 705
box -2 -3 58 103
use XNOR2X1  XNOR2X1_21
timestamp 1693479267
transform 1 0 1124 0 -1 705
box -2 -3 58 103
use NOR2X1  NOR2X1_31
timestamp 1693479267
transform 1 0 1180 0 -1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_18
timestamp 1693479267
transform 1 0 1204 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_32
timestamp 1693479267
transform -1 0 1260 0 -1 705
box -2 -3 26 103
use XNOR2X1  XNOR2X1_27
timestamp 1693479267
transform -1 0 1316 0 -1 705
box -2 -3 58 103
use NOR2X1  NOR2X1_34
timestamp 1693479267
transform -1 0 1340 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_35
timestamp 1693479267
transform -1 0 1364 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_145
timestamp 1693479267
transform 1 0 1364 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_48
timestamp 1693479267
transform 1 0 1388 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_33
timestamp 1693479267
transform -1 0 1436 0 -1 705
box -2 -3 26 103
use XNOR2X1  XNOR2X1_26
timestamp 1693479267
transform -1 0 1492 0 -1 705
box -2 -3 58 103
use OAI21X1  OAI21X1_250
timestamp 1693479267
transform 1 0 1492 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_2_0
timestamp 1693479267
transform 1 0 1524 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_2_1
timestamp 1693479267
transform 1 0 1532 0 -1 705
box -2 -3 10 103
use NOR3X1  NOR3X1_53
timestamp 1693479267
transform 1 0 1540 0 -1 705
box -2 -3 66 103
use AOI22X1  AOI22X1_49
timestamp 1693479267
transform 1 0 1604 0 -1 705
box -2 -3 42 103
use INVX1  INVX1_325
timestamp 1693479267
transform 1 0 1644 0 -1 705
box -2 -3 18 103
use INVX2  INVX2_34
timestamp 1693479267
transform -1 0 1676 0 -1 705
box -2 -3 18 103
use NOR2X1  NOR2X1_320
timestamp 1693479267
transform 1 0 1676 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_640
timestamp 1693479267
transform -1 0 1732 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_639
timestamp 1693479267
transform 1 0 1732 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_148
timestamp 1693479267
transform -1 0 1796 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_630
timestamp 1693479267
transform 1 0 1796 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_629
timestamp 1693479267
transform -1 0 1860 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_147
timestamp 1693479267
transform -1 0 1892 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_228
timestamp 1693479267
transform 1 0 1892 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_229
timestamp 1693479267
transform 1 0 1916 0 -1 705
box -2 -3 26 103
use NAND3X1  NAND3X1_146
timestamp 1693479267
transform 1 0 1940 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_403
timestamp 1693479267
transform 1 0 1972 0 -1 705
box -2 -3 18 103
use NOR2X1  NOR2X1_321
timestamp 1693479267
transform -1 0 2012 0 -1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_155
timestamp 1693479267
transform 1 0 2012 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_3_0
timestamp 1693479267
transform -1 0 2052 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_3_1
timestamp 1693479267
transform -1 0 2060 0 -1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_642
timestamp 1693479267
transform -1 0 2092 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_598
timestamp 1693479267
transform 1 0 2092 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_131
timestamp 1693479267
transform -1 0 2156 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_169
timestamp 1693479267
transform 1 0 2156 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_226
timestamp 1693479267
transform -1 0 2204 0 -1 705
box -2 -3 26 103
use OAI22X1  OAI22X1_39
timestamp 1693479267
transform -1 0 2244 0 -1 705
box -2 -3 42 103
use BUFX4  BUFX4_190
timestamp 1693479267
transform -1 0 2276 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_266
timestamp 1693479267
transform 1 0 2276 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_315
timestamp 1693479267
transform -1 0 2332 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_338
timestamp 1693479267
transform -1 0 2348 0 -1 705
box -2 -3 18 103
use MUX2X1  MUX2X1_11
timestamp 1693479267
transform 1 0 2348 0 -1 705
box -2 -3 50 103
use INVX1  INVX1_350
timestamp 1693479267
transform 1 0 2396 0 -1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_320
timestamp 1693479267
transform -1 0 2436 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_267
timestamp 1693479267
transform 1 0 2436 0 -1 705
box -2 -3 26 103
use BUFX4  BUFX4_275
timestamp 1693479267
transform -1 0 2492 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_462
timestamp 1693479267
transform -1 0 2516 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_230
timestamp 1693479267
transform 1 0 2516 0 -1 705
box -2 -3 26 103
use FILL  FILL_6_4_0
timestamp 1693479267
transform -1 0 2548 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_4_1
timestamp 1693479267
transform -1 0 2556 0 -1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_342
timestamp 1693479267
transform -1 0 2588 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_425
timestamp 1693479267
transform -1 0 2612 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_220
timestamp 1693479267
transform -1 0 2636 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_219
timestamp 1693479267
transform -1 0 2660 0 -1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_84
timestamp 1693479267
transform 1 0 2660 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_79
timestamp 1693479267
transform 1 0 2692 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_80
timestamp 1693479267
transform 1 0 2724 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_463
timestamp 1693479267
transform -1 0 2788 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_379
timestamp 1693479267
transform -1 0 2812 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_452
timestamp 1693479267
transform -1 0 2844 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_189
timestamp 1693479267
transform -1 0 2876 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_346
timestamp 1693479267
transform 1 0 2876 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_343
timestamp 1693479267
transform 1 0 2908 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_385
timestamp 1693479267
transform 1 0 2940 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_52
timestamp 1693479267
transform -1 0 3004 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_484
timestamp 1693479267
transform 1 0 3004 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_430
timestamp 1693479267
transform -1 0 3060 0 -1 705
box -2 -3 26 103
use FILL  FILL_6_5_0
timestamp 1693479267
transform 1 0 3060 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_5_1
timestamp 1693479267
transform 1 0 3068 0 -1 705
box -2 -3 10 103
use NAND2X1  NAND2X1_472
timestamp 1693479267
transform 1 0 3076 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_365
timestamp 1693479267
transform 1 0 3100 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_215
timestamp 1693479267
transform -1 0 3164 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_473
timestamp 1693479267
transform 1 0 3164 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_370
timestamp 1693479267
transform 1 0 3188 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_450
timestamp 1693479267
transform 1 0 3212 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_632
timestamp 1693479267
transform 1 0 3244 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_596
timestamp 1693479267
transform 1 0 3276 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_532
timestamp 1693479267
transform -1 0 3332 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_551
timestamp 1693479267
transform -1 0 3356 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_482
timestamp 1693479267
transform 1 0 3356 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_489
timestamp 1693479267
transform 1 0 3380 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_533
timestamp 1693479267
transform -1 0 3436 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_521
timestamp 1693479267
transform 1 0 3436 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_576
timestamp 1693479267
transform -1 0 3492 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_547
timestamp 1693479267
transform -1 0 3516 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_519
timestamp 1693479267
transform -1 0 3548 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_438
timestamp 1693479267
transform -1 0 3572 0 -1 705
box -2 -3 26 103
use FILL  FILL_6_6_0
timestamp 1693479267
transform 1 0 3572 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_6_1
timestamp 1693479267
transform 1 0 3580 0 -1 705
box -2 -3 10 103
use NAND2X1  NAND2X1_465
timestamp 1693479267
transform 1 0 3588 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_543
timestamp 1693479267
transform -1 0 3644 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_334
timestamp 1693479267
transform -1 0 3660 0 -1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_538
timestamp 1693479267
transform 1 0 3660 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_613
timestamp 1693479267
transform -1 0 3716 0 -1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_7
timestamp 1693479267
transform -1 0 3764 0 -1 705
box -2 -3 50 103
use BUFX4  BUFX4_214
timestamp 1693479267
transform -1 0 3796 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_123
timestamp 1693479267
transform 1 0 3796 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_556
timestamp 1693479267
transform -1 0 3844 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_487
timestamp 1693479267
transform -1 0 3868 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_270
timestamp 1693479267
transform -1 0 3892 0 -1 705
box -2 -3 26 103
use INVX2  INVX2_43
timestamp 1693479267
transform 1 0 3892 0 -1 705
box -2 -3 18 103
use NOR2X1  NOR2X1_122
timestamp 1693479267
transform 1 0 3908 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_268
timestamp 1693479267
transform -1 0 3956 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_301
timestamp 1693479267
transform 1 0 3956 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_488
timestamp 1693479267
transform 1 0 3980 0 -1 705
box -2 -3 26 103
use AOI22X1  AOI22X1_96
timestamp 1693479267
transform -1 0 4044 0 -1 705
box -2 -3 42 103
use OAI21X1  OAI21X1_328
timestamp 1693479267
transform -1 0 4076 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_7_0
timestamp 1693479267
transform 1 0 4076 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_7_1
timestamp 1693479267
transform 1 0 4084 0 -1 705
box -2 -3 10 103
use NAND2X1  NAND2X1_300
timestamp 1693479267
transform 1 0 4092 0 -1 705
box -2 -3 26 103
use OAI22X1  OAI22X1_9
timestamp 1693479267
transform -1 0 4156 0 -1 705
box -2 -3 42 103
use OAI22X1  OAI22X1_26
timestamp 1693479267
transform -1 0 4196 0 -1 705
box -2 -3 42 103
use AOI21X1  AOI21X1_109
timestamp 1693479267
transform -1 0 4228 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_94
timestamp 1693479267
transform 1 0 4228 0 -1 705
box -2 -3 34 103
use OAI22X1  OAI22X1_20
timestamp 1693479267
transform 1 0 4260 0 -1 705
box -2 -3 42 103
use NOR2X1  NOR2X1_253
timestamp 1693479267
transform 1 0 4300 0 -1 705
box -2 -3 26 103
use NAND3X1  NAND3X1_133
timestamp 1693479267
transform -1 0 4356 0 -1 705
box -2 -3 34 103
use INVX4  INVX4_8
timestamp 1693479267
transform 1 0 4356 0 -1 705
box -2 -3 26 103
use AND2X2  AND2X2_36
timestamp 1693479267
transform -1 0 4412 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_529
timestamp 1693479267
transform -1 0 4444 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_486
timestamp 1693479267
transform 1 0 4444 0 -1 705
box -2 -3 26 103
use NAND3X1  NAND3X1_123
timestamp 1693479267
transform -1 0 4500 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_526
timestamp 1693479267
transform 1 0 4500 0 -1 705
box -2 -3 34 103
use INVX2  INVX2_58
timestamp 1693479267
transform 1 0 4532 0 -1 705
box -2 -3 18 103
use AOI21X1  AOI21X1_101
timestamp 1693479267
transform 1 0 4548 0 -1 705
box -2 -3 34 103
use FILL  FILL_7_1
timestamp 1693479267
transform -1 0 4588 0 -1 705
box -2 -3 10 103
use FILL  FILL_7_2
timestamp 1693479267
transform -1 0 4596 0 -1 705
box -2 -3 10 103
use FILL  FILL_7_3
timestamp 1693479267
transform -1 0 4604 0 -1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_488
timestamp 1693479267
transform -1 0 100 0 1 705
box -2 -3 98 103
use INVX1  INVX1_479
timestamp 1693479267
transform 1 0 100 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_841
timestamp 1693479267
transform -1 0 148 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_842
timestamp 1693479267
transform -1 0 180 0 1 705
box -2 -3 34 103
use INVX1  INVX1_478
timestamp 1693479267
transform 1 0 180 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_839
timestamp 1693479267
transform 1 0 196 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_388
timestamp 1693479267
transform 1 0 228 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_840
timestamp 1693479267
transform 1 0 252 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_177
timestamp 1693479267
transform -1 0 316 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_39
timestamp 1693479267
transform -1 0 348 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_167
timestamp 1693479267
transform 1 0 348 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_822
timestamp 1693479267
transform -1 0 412 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_197
timestamp 1693479267
transform -1 0 444 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_243
timestamp 1693479267
transform -1 0 476 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_12
timestamp 1693479267
transform 1 0 476 0 1 705
box -2 -3 34 103
use FILL  FILL_7_0_0
timestamp 1693479267
transform 1 0 508 0 1 705
box -2 -3 10 103
use FILL  FILL_7_0_1
timestamp 1693479267
transform 1 0 516 0 1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_164
timestamp 1693479267
transform 1 0 524 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_666
timestamp 1693479267
transform 1 0 556 0 1 705
box -2 -3 26 103
use OR2X2  OR2X2_45
timestamp 1693479267
transform 1 0 580 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_818
timestamp 1693479267
transform 1 0 612 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_200
timestamp 1693479267
transform 1 0 644 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_642
timestamp 1693479267
transform -1 0 700 0 1 705
box -2 -3 26 103
use BUFX4  BUFX4_245
timestamp 1693479267
transform 1 0 700 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_668
timestamp 1693479267
transform 1 0 732 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_646
timestamp 1693479267
transform 1 0 756 0 1 705
box -2 -3 26 103
use BUFX2  BUFX2_18
timestamp 1693479267
transform -1 0 804 0 1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_175
timestamp 1693479267
transform -1 0 900 0 1 705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_177
timestamp 1693479267
transform 1 0 900 0 1 705
box -2 -3 98 103
use FILL  FILL_7_1_0
timestamp 1693479267
transform 1 0 996 0 1 705
box -2 -3 10 103
use FILL  FILL_7_1_1
timestamp 1693479267
transform 1 0 1004 0 1 705
box -2 -3 10 103
use XNOR2X1  XNOR2X1_23
timestamp 1693479267
transform 1 0 1012 0 1 705
box -2 -3 58 103
use NAND2X1  NAND2X1_144
timestamp 1693479267
transform 1 0 1068 0 1 705
box -2 -3 26 103
use XNOR2X1  XNOR2X1_24
timestamp 1693479267
transform -1 0 1148 0 1 705
box -2 -3 58 103
use INVX2  INVX2_9
timestamp 1693479267
transform 1 0 1148 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_246
timestamp 1693479267
transform 1 0 1164 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_247
timestamp 1693479267
transform 1 0 1196 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_38
timestamp 1693479267
transform 1 0 1228 0 1 705
box -2 -3 26 103
use INVX2  INVX2_10
timestamp 1693479267
transform 1 0 1252 0 1 705
box -2 -3 18 103
use XNOR2X1  XNOR2X1_18
timestamp 1693479267
transform 1 0 1268 0 1 705
box -2 -3 58 103
use NAND2X1  NAND2X1_143
timestamp 1693479267
transform 1 0 1324 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_142
timestamp 1693479267
transform 1 0 1348 0 1 705
box -2 -3 26 103
use XNOR2X1  XNOR2X1_19
timestamp 1693479267
transform 1 0 1372 0 1 705
box -2 -3 58 103
use NAND2X1  NAND2X1_141
timestamp 1693479267
transform -1 0 1452 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_245
timestamp 1693479267
transform -1 0 1484 0 1 705
box -2 -3 34 103
use INVX1  INVX1_258
timestamp 1693479267
transform 1 0 1484 0 1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_146
timestamp 1693479267
transform 1 0 1500 0 1 705
box -2 -3 26 103
use FILL  FILL_7_2_0
timestamp 1693479267
transform -1 0 1532 0 1 705
box -2 -3 10 103
use FILL  FILL_7_2_1
timestamp 1693479267
transform -1 0 1540 0 1 705
box -2 -3 10 103
use AOI21X1  AOI21X1_20
timestamp 1693479267
transform -1 0 1572 0 1 705
box -2 -3 34 103
use NOR3X1  NOR3X1_54
timestamp 1693479267
transform -1 0 1636 0 1 705
box -2 -3 66 103
use NAND2X1  NAND2X1_225
timestamp 1693479267
transform 1 0 1636 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_94
timestamp 1693479267
transform 1 0 1660 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_644
timestamp 1693479267
transform 1 0 1684 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_317
timestamp 1693479267
transform -1 0 1740 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_319
timestamp 1693479267
transform 1 0 1740 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_37
timestamp 1693479267
transform -1 0 1796 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_303
timestamp 1693479267
transform -1 0 1828 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_95
timestamp 1693479267
transform -1 0 1852 0 1 705
box -2 -3 26 103
use INVX2  INVX2_35
timestamp 1693479267
transform 1 0 1852 0 1 705
box -2 -3 18 103
use NAND3X1  NAND3X1_149
timestamp 1693479267
transform 1 0 1868 0 1 705
box -2 -3 34 103
use AND2X2  AND2X2_48
timestamp 1693479267
transform -1 0 1932 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_620
timestamp 1693479267
transform 1 0 1932 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_313
timestamp 1693479267
transform -1 0 1988 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_230
timestamp 1693479267
transform -1 0 2012 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_227
timestamp 1693479267
transform -1 0 2036 0 1 705
box -2 -3 26 103
use FILL  FILL_7_3_0
timestamp 1693479267
transform 1 0 2036 0 1 705
box -2 -3 10 103
use FILL  FILL_7_3_1
timestamp 1693479267
transform 1 0 2044 0 1 705
box -2 -3 10 103
use NAND2X1  NAND2X1_224
timestamp 1693479267
transform 1 0 2052 0 1 705
box -2 -3 26 103
use INVX1  INVX1_402
timestamp 1693479267
transform 1 0 2076 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_591
timestamp 1693479267
transform 1 0 2092 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_595
timestamp 1693479267
transform 1 0 2124 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_135
timestamp 1693479267
transform -1 0 2188 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_625
timestamp 1693479267
transform 1 0 2188 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_153
timestamp 1693479267
transform 1 0 2220 0 1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_42
timestamp 1693479267
transform 1 0 2252 0 1 705
box -2 -3 50 103
use NAND2X1  NAND2X1_270
timestamp 1693479267
transform 1 0 2300 0 1 705
box -2 -3 26 103
use OR2X2  OR2X2_18
timestamp 1693479267
transform 1 0 2324 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_76
timestamp 1693479267
transform 1 0 2356 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_47
timestamp 1693479267
transform 1 0 2388 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_459
timestamp 1693479267
transform 1 0 2420 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_74
timestamp 1693479267
transform -1 0 2484 0 1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_24
timestamp 1693479267
transform 1 0 2484 0 1 705
box -2 -3 50 103
use NAND2X1  NAND2X1_324
timestamp 1693479267
transform -1 0 2556 0 1 705
box -2 -3 26 103
use FILL  FILL_7_4_0
timestamp 1693479267
transform 1 0 2556 0 1 705
box -2 -3 10 103
use FILL  FILL_7_4_1
timestamp 1693479267
transform 1 0 2564 0 1 705
box -2 -3 10 103
use NAND3X1  NAND3X1_115
timestamp 1693479267
transform 1 0 2572 0 1 705
box -2 -3 34 103
use OR2X2  OR2X2_28
timestamp 1693479267
transform 1 0 2604 0 1 705
box -2 -3 34 103
use AOI22X1  AOI22X1_84
timestamp 1693479267
transform 1 0 2636 0 1 705
box -2 -3 42 103
use NAND2X1  NAND2X1_461
timestamp 1693479267
transform 1 0 2676 0 1 705
box -2 -3 26 103
use AOI22X1  AOI22X1_83
timestamp 1693479267
transform -1 0 2740 0 1 705
box -2 -3 42 103
use NAND2X1  NAND2X1_436
timestamp 1693479267
transform 1 0 2740 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_75
timestamp 1693479267
transform -1 0 2796 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_368
timestamp 1693479267
transform 1 0 2796 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_354
timestamp 1693479267
transform 1 0 2820 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_50
timestamp 1693479267
transform 1 0 2852 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_384
timestamp 1693479267
transform 1 0 2884 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_631
timestamp 1693479267
transform -1 0 2948 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_369
timestamp 1693479267
transform 1 0 2948 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_441
timestamp 1693479267
transform 1 0 2972 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_83
timestamp 1693479267
transform -1 0 3028 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_90
timestamp 1693479267
transform -1 0 3060 0 1 705
box -2 -3 34 103
use FILL  FILL_7_5_0
timestamp 1693479267
transform 1 0 3060 0 1 705
box -2 -3 10 103
use FILL  FILL_7_5_1
timestamp 1693479267
transform 1 0 3068 0 1 705
box -2 -3 10 103
use INVX1  INVX1_362
timestamp 1693479267
transform 1 0 3076 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_461
timestamp 1693479267
transform 1 0 3092 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_434
timestamp 1693479267
transform 1 0 3124 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_469
timestamp 1693479267
transform 1 0 3148 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_442
timestamp 1693479267
transform -1 0 3196 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_386
timestamp 1693479267
transform -1 0 3228 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_342
timestamp 1693479267
transform -1 0 3252 0 1 705
box -2 -3 26 103
use INVX1  INVX1_384
timestamp 1693479267
transform -1 0 3268 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_498
timestamp 1693479267
transform 1 0 3268 0 1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_43
timestamp 1693479267
transform 1 0 3300 0 1 705
box -2 -3 50 103
use BUFX4  BUFX4_217
timestamp 1693479267
transform 1 0 3348 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_437
timestamp 1693479267
transform -1 0 3404 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_234
timestamp 1693479267
transform 1 0 3404 0 1 705
box -2 -3 26 103
use MUX2X1  MUX2X1_25
timestamp 1693479267
transform 1 0 3428 0 1 705
box -2 -3 50 103
use OAI21X1  OAI21X1_621
timestamp 1693479267
transform 1 0 3476 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_541
timestamp 1693479267
transform -1 0 3532 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_633
timestamp 1693479267
transform -1 0 3564 0 1 705
box -2 -3 34 103
use FILL  FILL_7_6_0
timestamp 1693479267
transform -1 0 3572 0 1 705
box -2 -3 10 103
use FILL  FILL_7_6_1
timestamp 1693479267
transform -1 0 3580 0 1 705
box -2 -3 10 103
use INVX1  INVX1_404
timestamp 1693479267
transform -1 0 3596 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_496
timestamp 1693479267
transform -1 0 3628 0 1 705
box -2 -3 34 103
use AND2X2  AND2X2_32
timestamp 1693479267
transform 1 0 3628 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_216
timestamp 1693479267
transform -1 0 3692 0 1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_38
timestamp 1693479267
transform -1 0 3740 0 1 705
box -2 -3 50 103
use NAND2X1  NAND2X1_374
timestamp 1693479267
transform 1 0 3740 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_390
timestamp 1693479267
transform -1 0 3796 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_91
timestamp 1693479267
transform -1 0 3828 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_135
timestamp 1693479267
transform 1 0 3828 0 1 705
box -2 -3 34 103
use INVX1  INVX1_365
timestamp 1693479267
transform 1 0 3860 0 1 705
box -2 -3 18 103
use INVX8  INVX8_4
timestamp 1693479267
transform -1 0 3916 0 1 705
box -2 -3 42 103
use BUFX4  BUFX4_274
timestamp 1693479267
transform -1 0 3948 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_92
timestamp 1693479267
transform 1 0 3948 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_122
timestamp 1693479267
transform -1 0 4012 0 1 705
box -2 -3 34 103
use AOI22X1  AOI22X1_90
timestamp 1693479267
transform -1 0 4052 0 1 705
box -2 -3 42 103
use AOI21X1  AOI21X1_100
timestamp 1693479267
transform -1 0 4084 0 1 705
box -2 -3 34 103
use FILL  FILL_7_7_0
timestamp 1693479267
transform 1 0 4084 0 1 705
box -2 -3 10 103
use FILL  FILL_7_7_1
timestamp 1693479267
transform 1 0 4092 0 1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_504
timestamp 1693479267
transform 1 0 4100 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_92
timestamp 1693479267
transform -1 0 4164 0 1 705
box -2 -3 34 103
use INVX1  INVX1_393
timestamp 1693479267
transform 1 0 4164 0 1 705
box -2 -3 18 103
use NAND3X1  NAND3X1_129
timestamp 1693479267
transform 1 0 4180 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_130
timestamp 1693479267
transform 1 0 4212 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_540
timestamp 1693479267
transform -1 0 4276 0 1 705
box -2 -3 34 103
use INVX1  INVX1_392
timestamp 1693479267
transform -1 0 4292 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_539
timestamp 1693479267
transform -1 0 4324 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_139
timestamp 1693479267
transform -1 0 4356 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_254
timestamp 1693479267
transform -1 0 4380 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_103
timestamp 1693479267
transform -1 0 4412 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_528
timestamp 1693479267
transform -1 0 4444 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_525
timestamp 1693479267
transform 1 0 4444 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_102
timestamp 1693479267
transform 1 0 4476 0 1 705
box -2 -3 34 103
use AOI22X1  AOI22X1_92
timestamp 1693479267
transform -1 0 4548 0 1 705
box -2 -3 42 103
use XNOR2X1  XNOR2X1_49
timestamp 1693479267
transform 1 0 4548 0 1 705
box -2 -3 58 103
use BUFX2  BUFX2_57
timestamp 1693479267
transform -1 0 28 0 -1 905
box -2 -3 26 103
use BUFX2  BUFX2_6
timestamp 1693479267
transform -1 0 52 0 -1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_163
timestamp 1693479267
transform -1 0 148 0 -1 905
box -2 -3 98 103
use CLKBUF1  CLKBUF1_35
timestamp 1693479267
transform -1 0 220 0 -1 905
box -2 -3 74 103
use NAND2X1  NAND2X1_669
timestamp 1693479267
transform 1 0 220 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_217
timestamp 1693479267
transform 1 0 244 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_456
timestamp 1693479267
transform 1 0 276 0 -1 905
box -2 -3 98 103
use CLKBUF1  CLKBUF1_45
timestamp 1693479267
transform -1 0 444 0 -1 905
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_490
timestamp 1693479267
transform -1 0 540 0 -1 905
box -2 -3 98 103
use FILL  FILL_8_0_0
timestamp 1693479267
transform 1 0 540 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_0_1
timestamp 1693479267
transform 1 0 548 0 -1 905
box -2 -3 10 103
use NAND3X1  NAND3X1_43
timestamp 1693479267
transform 1 0 556 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_458
timestamp 1693479267
transform 1 0 588 0 -1 905
box -2 -3 98 103
use NAND3X1  NAND3X1_42
timestamp 1693479267
transform 1 0 684 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_38
timestamp 1693479267
transform 1 0 716 0 -1 905
box -2 -3 34 103
use INVX8  INVX8_2
timestamp 1693479267
transform 1 0 748 0 -1 905
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_270
timestamp 1693479267
transform 1 0 788 0 -1 905
box -2 -3 98 103
use XOR2X1  XOR2X1_3
timestamp 1693479267
transform -1 0 940 0 -1 905
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_272
timestamp 1693479267
transform 1 0 940 0 -1 905
box -2 -3 98 103
use FILL  FILL_8_1_0
timestamp 1693479267
transform -1 0 1044 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_1_1
timestamp 1693479267
transform -1 0 1052 0 -1 905
box -2 -3 10 103
use XNOR2X1  XNOR2X1_36
timestamp 1693479267
transform -1 0 1108 0 -1 905
box -2 -3 58 103
use NAND2X1  NAND2X1_152
timestamp 1693479267
transform 1 0 1108 0 -1 905
box -2 -3 26 103
use INVX1  INVX1_259
timestamp 1693479267
transform -1 0 1148 0 -1 905
box -2 -3 18 103
use AOI21X1  AOI21X1_24
timestamp 1693479267
transform -1 0 1180 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_154
timestamp 1693479267
transform -1 0 1204 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_23
timestamp 1693479267
transform -1 0 1236 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_150
timestamp 1693479267
transform 1 0 1236 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_157
timestamp 1693479267
transform -1 0 1284 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_267
timestamp 1693479267
transform 1 0 1284 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_242
timestamp 1693479267
transform 1 0 1316 0 -1 905
box -2 -3 34 103
use XNOR2X1  XNOR2X1_20
timestamp 1693479267
transform -1 0 1404 0 -1 905
box -2 -3 58 103
use OAI21X1  OAI21X1_243
timestamp 1693479267
transform -1 0 1436 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_244
timestamp 1693479267
transform -1 0 1468 0 -1 905
box -2 -3 34 103
use INVX2  INVX2_8
timestamp 1693479267
transform -1 0 1484 0 -1 905
box -2 -3 18 103
use XNOR2X1  XNOR2X1_17
timestamp 1693479267
transform -1 0 1540 0 -1 905
box -2 -3 58 103
use FILL  FILL_8_2_0
timestamp 1693479267
transform -1 0 1548 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_2_1
timestamp 1693479267
transform -1 0 1556 0 -1 905
box -2 -3 10 103
use AOI21X1  AOI21X1_15
timestamp 1693479267
transform -1 0 1588 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_255
timestamp 1693479267
transform -1 0 1604 0 -1 905
box -2 -3 18 103
use AOI22X1  AOI22X1_54
timestamp 1693479267
transform 1 0 1604 0 -1 905
box -2 -3 42 103
use BUFX4  BUFX4_235
timestamp 1693479267
transform -1 0 1676 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_327
timestamp 1693479267
transform 1 0 1676 0 -1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_300
timestamp 1693479267
transform 1 0 1692 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_645
timestamp 1693479267
transform -1 0 1756 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_178
timestamp 1693479267
transform -1 0 1788 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_415
timestamp 1693479267
transform -1 0 1804 0 -1 905
box -2 -3 18 103
use MUX2X1  MUX2X1_2
timestamp 1693479267
transform -1 0 1852 0 -1 905
box -2 -3 50 103
use INVX1  INVX1_407
timestamp 1693479267
transform 1 0 1852 0 -1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_646
timestamp 1693479267
transform -1 0 1900 0 -1 905
box -2 -3 34 103
use OR2X2  OR2X2_39
timestamp 1693479267
transform 1 0 1900 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_337
timestamp 1693479267
transform 1 0 1932 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_158
timestamp 1693479267
transform -1 0 1988 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_104
timestamp 1693479267
transform -1 0 2012 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_577
timestamp 1693479267
transform -1 0 2036 0 -1 905
box -2 -3 26 103
use FILL  FILL_8_3_0
timestamp 1693479267
transform 1 0 2036 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_3_1
timestamp 1693479267
transform 1 0 2044 0 -1 905
box -2 -3 10 103
use AND2X2  AND2X2_52
timestamp 1693479267
transform 1 0 2052 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_544
timestamp 1693479267
transform 1 0 2084 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_316
timestamp 1693479267
transform 1 0 2108 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_180
timestamp 1693479267
transform -1 0 2172 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_70
timestamp 1693479267
transform -1 0 2204 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_71
timestamp 1693479267
transform 1 0 2204 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_373
timestamp 1693479267
transform -1 0 2252 0 -1 905
box -2 -3 18 103
use AOI21X1  AOI21X1_72
timestamp 1693479267
transform 1 0 2252 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_447
timestamp 1693479267
transform -1 0 2316 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_514
timestamp 1693479267
transform 1 0 2316 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_448
timestamp 1693479267
transform 1 0 2348 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_410
timestamp 1693479267
transform -1 0 2404 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_268
timestamp 1693479267
transform 1 0 2404 0 -1 905
box -2 -3 26 103
use AOI22X1  AOI22X1_73
timestamp 1693479267
transform -1 0 2468 0 -1 905
box -2 -3 42 103
use AOI21X1  AOI21X1_97
timestamp 1693479267
transform -1 0 2500 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_464
timestamp 1693479267
transform 1 0 2500 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_276
timestamp 1693479267
transform -1 0 2556 0 -1 905
box -2 -3 26 103
use FILL  FILL_8_4_0
timestamp 1693479267
transform -1 0 2564 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_4_1
timestamp 1693479267
transform -1 0 2572 0 -1 905
box -2 -3 10 103
use AOI22X1  AOI22X1_81
timestamp 1693479267
transform -1 0 2612 0 -1 905
box -2 -3 42 103
use NAND2X1  NAND2X1_265
timestamp 1693479267
transform -1 0 2636 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_426
timestamp 1693479267
transform -1 0 2660 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_275
timestamp 1693479267
transform -1 0 2684 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_140
timestamp 1693479267
transform 1 0 2684 0 -1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_111
timestamp 1693479267
transform -1 0 2740 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_449
timestamp 1693479267
transform 1 0 2740 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_392
timestamp 1693479267
transform 1 0 2772 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_378
timestamp 1693479267
transform 1 0 2804 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_73
timestamp 1693479267
transform -1 0 2860 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_323
timestamp 1693479267
transform -1 0 2884 0 -1 905
box -2 -3 26 103
use BUFX4  BUFX4_77
timestamp 1693479267
transform -1 0 2916 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_58
timestamp 1693479267
transform 1 0 2916 0 -1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_21
timestamp 1693479267
transform 1 0 2948 0 -1 905
box -2 -3 50 103
use NAND3X1  NAND3X1_119
timestamp 1693479267
transform 1 0 2996 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_374
timestamp 1693479267
transform -1 0 3044 0 -1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_540
timestamp 1693479267
transform 1 0 3044 0 -1 905
box -2 -3 26 103
use FILL  FILL_8_5_0
timestamp 1693479267
transform 1 0 3068 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_5_1
timestamp 1693479267
transform 1 0 3076 0 -1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_445
timestamp 1693479267
transform 1 0 3084 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_363
timestamp 1693479267
transform -1 0 3148 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_339
timestamp 1693479267
transform -1 0 3172 0 -1 905
box -2 -3 26 103
use BUFX4  BUFX4_79
timestamp 1693479267
transform 1 0 3172 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_453
timestamp 1693479267
transform -1 0 3236 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_507
timestamp 1693479267
transform 1 0 3236 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_648
timestamp 1693479267
transform 1 0 3268 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_454
timestamp 1693479267
transform 1 0 3300 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_455
timestamp 1693479267
transform -1 0 3364 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_506
timestamp 1693479267
transform -1 0 3396 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_420
timestamp 1693479267
transform -1 0 3420 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_485
timestamp 1693479267
transform -1 0 3452 0 -1 905
box -2 -3 34 103
use BUFX4  BUFX4_213
timestamp 1693479267
transform -1 0 3484 0 -1 905
box -2 -3 34 103
use BUFX4  BUFX4_228
timestamp 1693479267
transform -1 0 3516 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_136
timestamp 1693479267
transform -1 0 3548 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_550
timestamp 1693479267
transform -1 0 3572 0 -1 905
box -2 -3 26 103
use FILL  FILL_8_6_0
timestamp 1693479267
transform 1 0 3572 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_6_1
timestamp 1693479267
transform 1 0 3580 0 -1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_649
timestamp 1693479267
transform 1 0 3588 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_650
timestamp 1693479267
transform -1 0 3652 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_187
timestamp 1693479267
transform -1 0 3676 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_362
timestamp 1693479267
transform 1 0 3676 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_471
timestamp 1693479267
transform 1 0 3700 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_238
timestamp 1693479267
transform -1 0 3756 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_222
timestamp 1693479267
transform -1 0 3780 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_424
timestamp 1693479267
transform -1 0 3804 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_546
timestamp 1693479267
transform -1 0 3828 0 -1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_34
timestamp 1693479267
transform 1 0 3828 0 -1 905
box -2 -3 50 103
use OAI21X1  OAI21X1_614
timestamp 1693479267
transform 1 0 3876 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_539
timestamp 1693479267
transform -1 0 3932 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_126
timestamp 1693479267
transform 1 0 3932 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_477
timestamp 1693479267
transform -1 0 3988 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_375
timestamp 1693479267
transform -1 0 4012 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_522
timestamp 1693479267
transform 1 0 4012 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_520
timestamp 1693479267
transform 1 0 4044 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_7_0
timestamp 1693479267
transform -1 0 4084 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_7_1
timestamp 1693479267
transform -1 0 4092 0 -1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_570
timestamp 1693479267
transform -1 0 4124 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_118
timestamp 1693479267
transform 1 0 4124 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_95
timestamp 1693479267
transform 1 0 4156 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_509
timestamp 1693479267
transform 1 0 4188 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_241
timestamp 1693479267
transform -1 0 4244 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_568
timestamp 1693479267
transform -1 0 4276 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_284
timestamp 1693479267
transform 1 0 4276 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_295
timestamp 1693479267
transform 1 0 4300 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_128
timestamp 1693479267
transform 1 0 4324 0 -1 905
box -2 -3 34 103
use OR2X2  OR2X2_35
timestamp 1693479267
transform -1 0 4388 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_587
timestamp 1693479267
transform -1 0 4420 0 -1 905
box -2 -3 34 103
use INVX2  INVX2_59
timestamp 1693479267
transform 1 0 4420 0 -1 905
box -2 -3 18 103
use INVX2  INVX2_60
timestamp 1693479267
transform 1 0 4436 0 -1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_541
timestamp 1693479267
transform 1 0 4452 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_107
timestamp 1693479267
transform -1 0 4516 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_269
timestamp 1693479267
transform 1 0 4516 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_255
timestamp 1693479267
transform -1 0 4564 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_530
timestamp 1693479267
transform 1 0 4564 0 -1 905
box -2 -3 34 103
use FILL  FILL_9_1
timestamp 1693479267
transform -1 0 4604 0 -1 905
box -2 -3 10 103
use BUFX2  BUFX2_7
timestamp 1693479267
transform -1 0 28 0 1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_164
timestamp 1693479267
transform -1 0 124 0 1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_671
timestamp 1693479267
transform 1 0 124 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_390
timestamp 1693479267
transform -1 0 172 0 1 905
box -2 -3 26 103
use INVX1  INVX1_480
timestamp 1693479267
transform 1 0 172 0 1 905
box -2 -3 18 103
use INVX1  INVX1_481
timestamp 1693479267
transform 1 0 188 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_844
timestamp 1693479267
transform -1 0 236 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_846
timestamp 1693479267
transform 1 0 236 0 1 905
box -2 -3 34 103
use INVX1  INVX1_482
timestamp 1693479267
transform -1 0 284 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_845
timestamp 1693479267
transform 1 0 284 0 1 905
box -2 -3 34 103
use INVX8  INVX8_13
timestamp 1693479267
transform 1 0 316 0 1 905
box -2 -3 42 103
use OAI21X1  OAI21X1_179
timestamp 1693479267
transform -1 0 388 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_647
timestamp 1693479267
transform -1 0 412 0 1 905
box -2 -3 26 103
use BUFX4  BUFX4_247
timestamp 1693479267
transform -1 0 444 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_163
timestamp 1693479267
transform 1 0 444 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_11
timestamp 1693479267
transform -1 0 508 0 1 905
box -2 -3 34 103
use FILL  FILL_9_0_0
timestamp 1693479267
transform 1 0 508 0 1 905
box -2 -3 10 103
use FILL  FILL_9_0_1
timestamp 1693479267
transform 1 0 516 0 1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_474
timestamp 1693479267
transform 1 0 524 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_817
timestamp 1693479267
transform 1 0 620 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_10
timestamp 1693479267
transform -1 0 684 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_442
timestamp 1693479267
transform -1 0 780 0 1 905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_256
timestamp 1693479267
transform 1 0 780 0 1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_155
timestamp 1693479267
transform 1 0 876 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_43
timestamp 1693479267
transform 1 0 900 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_255
timestamp 1693479267
transform -1 0 956 0 1 905
box -2 -3 34 103
use INVX1  INVX1_260
timestamp 1693479267
transform -1 0 972 0 1 905
box -2 -3 18 103
use NOR2X1  NOR2X1_41
timestamp 1693479267
transform -1 0 996 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_151
timestamp 1693479267
transform 1 0 996 0 1 905
box -2 -3 26 103
use FILL  FILL_9_1_0
timestamp 1693479267
transform 1 0 1020 0 1 905
box -2 -3 10 103
use FILL  FILL_9_1_1
timestamp 1693479267
transform 1 0 1028 0 1 905
box -2 -3 10 103
use INVX1  INVX1_263
timestamp 1693479267
transform 1 0 1036 0 1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_158
timestamp 1693479267
transform 1 0 1052 0 1 905
box -2 -3 26 103
use XNOR2X1  XNOR2X1_13
timestamp 1693479267
transform 1 0 1076 0 1 905
box -2 -3 58 103
use OAI21X1  OAI21X1_254
timestamp 1693479267
transform -1 0 1164 0 1 905
box -2 -3 34 103
use XNOR2X1  XNOR2X1_15
timestamp 1693479267
transform 1 0 1164 0 1 905
box -2 -3 58 103
use NOR2X1  NOR2X1_30
timestamp 1693479267
transform 1 0 1220 0 1 905
box -2 -3 26 103
use INVX1  INVX1_253
timestamp 1693479267
transform 1 0 1244 0 1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_140
timestamp 1693479267
transform 1 0 1260 0 1 905
box -2 -3 26 103
use INVX1  INVX1_247
timestamp 1693479267
transform 1 0 1284 0 1 905
box -2 -3 18 103
use NOR3X1  NOR3X1_51
timestamp 1693479267
transform -1 0 1364 0 1 905
box -2 -3 66 103
use AOI21X1  AOI21X1_19
timestamp 1693479267
transform 1 0 1364 0 1 905
box -2 -3 34 103
use INVX1  INVX1_256
timestamp 1693479267
transform -1 0 1412 0 1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_133
timestamp 1693479267
transform 1 0 1412 0 1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_16
timestamp 1693479267
transform 1 0 1436 0 1 905
box -2 -3 34 103
use AOI22X1  AOI22X1_53
timestamp 1693479267
transform 1 0 1468 0 1 905
box -2 -3 42 103
use NAND2X1  NAND2X1_232
timestamp 1693479267
transform -1 0 1532 0 1 905
box -2 -3 26 103
use FILL  FILL_9_2_0
timestamp 1693479267
transform 1 0 1532 0 1 905
box -2 -3 10 103
use FILL  FILL_9_2_1
timestamp 1693479267
transform 1 0 1540 0 1 905
box -2 -3 10 103
use NAND2X1  NAND2X1_223
timestamp 1693479267
transform 1 0 1548 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_298
timestamp 1693479267
transform -1 0 1604 0 1 905
box -2 -3 34 103
use INVX1  INVX1_324
timestamp 1693479267
transform -1 0 1620 0 1 905
box -2 -3 18 103
use BUFX4  BUFX4_151
timestamp 1693479267
transform 1 0 1620 0 1 905
box -2 -3 34 103
use INVX2  INVX2_33
timestamp 1693479267
transform 1 0 1652 0 1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_240
timestamp 1693479267
transform -1 0 1692 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_697
timestamp 1693479267
transform -1 0 1724 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_186
timestamp 1693479267
transform 1 0 1724 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_712
timestamp 1693479267
transform -1 0 1788 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_39
timestamp 1693479267
transform 1 0 1788 0 1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_12
timestamp 1693479267
transform 1 0 1820 0 1 905
box -2 -3 50 103
use NAND3X1  NAND3X1_142
timestamp 1693479267
transform -1 0 1900 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_269
timestamp 1693479267
transform -1 0 1924 0 1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_145
timestamp 1693479267
transform -1 0 1956 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_87
timestamp 1693479267
transform -1 0 1988 0 1 905
box -2 -3 34 103
use INVX1  INVX1_339
timestamp 1693479267
transform 1 0 1988 0 1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_423
timestamp 1693479267
transform -1 0 2028 0 1 905
box -2 -3 26 103
use FILL  FILL_9_3_0
timestamp 1693479267
transform -1 0 2036 0 1 905
box -2 -3 10 103
use FILL  FILL_9_3_1
timestamp 1693479267
transform -1 0 2044 0 1 905
box -2 -3 10 103
use NAND3X1  NAND3X1_141
timestamp 1693479267
transform -1 0 2076 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_143
timestamp 1693479267
transform 1 0 2076 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_214
timestamp 1693479267
transform -1 0 2132 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_446
timestamp 1693479267
transform -1 0 2164 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_64
timestamp 1693479267
transform -1 0 2196 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_141
timestamp 1693479267
transform -1 0 2220 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_411
timestamp 1693479267
transform -1 0 2244 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_211
timestamp 1693479267
transform -1 0 2268 0 1 905
box -2 -3 26 103
use OAI22X1  OAI22X1_10
timestamp 1693479267
transform -1 0 2308 0 1 905
box -2 -3 42 103
use OAI22X1  OAI22X1_21
timestamp 1693479267
transform -1 0 2348 0 1 905
box -2 -3 42 103
use AOI21X1  AOI21X1_78
timestamp 1693479267
transform 1 0 2348 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_319
timestamp 1693479267
transform 1 0 2380 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_110
timestamp 1693479267
transform -1 0 2436 0 1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_40
timestamp 1693479267
transform -1 0 2468 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_77
timestamp 1693479267
transform 1 0 2468 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_109
timestamp 1693479267
transform 1 0 2500 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_466
timestamp 1693479267
transform -1 0 2556 0 1 905
box -2 -3 34 103
use FILL  FILL_9_4_0
timestamp 1693479267
transform -1 0 2564 0 1 905
box -2 -3 10 103
use FILL  FILL_9_4_1
timestamp 1693479267
transform -1 0 2572 0 1 905
box -2 -3 10 103
use INVX2  INVX2_52
timestamp 1693479267
transform -1 0 2588 0 1 905
box -2 -3 18 103
use AOI21X1  AOI21X1_147
timestamp 1693479267
transform -1 0 2620 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_332
timestamp 1693479267
transform -1 0 2652 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_198
timestamp 1693479267
transform 1 0 2652 0 1 905
box -2 -3 26 103
use BUFX4  BUFX4_86
timestamp 1693479267
transform 1 0 2676 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_153
timestamp 1693479267
transform 1 0 2708 0 1 905
box -2 -3 34 103
use AOI22X1  AOI22X1_80
timestamp 1693479267
transform 1 0 2740 0 1 905
box -2 -3 42 103
use NOR2X1  NOR2X1_188
timestamp 1693479267
transform 1 0 2780 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_533
timestamp 1693479267
transform 1 0 2804 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_299
timestamp 1693479267
transform -1 0 2852 0 1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_137
timestamp 1693479267
transform -1 0 2884 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_300
timestamp 1693479267
transform 1 0 2884 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_408
timestamp 1693479267
transform -1 0 2932 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_423
timestamp 1693479267
transform -1 0 2964 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_140
timestamp 1693479267
transform -1 0 2996 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_599
timestamp 1693479267
transform -1 0 3028 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_139
timestamp 1693479267
transform -1 0 3060 0 1 905
box -2 -3 34 103
use FILL  FILL_9_5_0
timestamp 1693479267
transform -1 0 3068 0 1 905
box -2 -3 10 103
use FILL  FILL_9_5_1
timestamp 1693479267
transform -1 0 3076 0 1 905
box -2 -3 10 103
use AND2X2  AND2X2_31
timestamp 1693479267
transform -1 0 3108 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_68
timestamp 1693479267
transform -1 0 3140 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_444
timestamp 1693479267
transform -1 0 3172 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_597
timestamp 1693479267
transform -1 0 3204 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_215
timestamp 1693479267
transform 1 0 3204 0 1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_138
timestamp 1693479267
transform -1 0 3260 0 1 905
box -2 -3 34 103
use INVX2  INVX2_66
timestamp 1693479267
transform -1 0 3276 0 1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_458
timestamp 1693479267
transform -1 0 3300 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_468
timestamp 1693479267
transform 1 0 3300 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_638
timestamp 1693479267
transform -1 0 3356 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_54
timestamp 1693479267
transform -1 0 3388 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_437
timestamp 1693479267
transform 1 0 3388 0 1 905
box -2 -3 34 103
use AND2X2  AND2X2_55
timestamp 1693479267
transform 1 0 3420 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_665
timestamp 1693479267
transform -1 0 3484 0 1 905
box -2 -3 34 103
use OR2X2  OR2X2_37
timestamp 1693479267
transform 1 0 3484 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_154
timestamp 1693479267
transform -1 0 3548 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_637
timestamp 1693479267
transform 1 0 3548 0 1 905
box -2 -3 34 103
use FILL  FILL_9_6_0
timestamp 1693479267
transform -1 0 3588 0 1 905
box -2 -3 10 103
use FILL  FILL_9_6_1
timestamp 1693479267
transform -1 0 3596 0 1 905
box -2 -3 10 103
use NOR2X1  NOR2X1_318
timestamp 1693479267
transform -1 0 3620 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_635
timestamp 1693479267
transform 1 0 3620 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_685
timestamp 1693479267
transform 1 0 3652 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_549
timestamp 1693479267
transform 1 0 3684 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_634
timestamp 1693479267
transform 1 0 3708 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_636
timestamp 1693479267
transform 1 0 3740 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_438
timestamp 1693479267
transform 1 0 3772 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_152
timestamp 1693479267
transform -1 0 3836 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_164
timestamp 1693479267
transform 1 0 3836 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_664
timestamp 1693479267
transform -1 0 3900 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_443
timestamp 1693479267
transform 1 0 3900 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_422
timestamp 1693479267
transform -1 0 3956 0 1 905
box -2 -3 26 103
use BUFX4  BUFX4_51
timestamp 1693479267
transform -1 0 3988 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_391
timestamp 1693479267
transform -1 0 4020 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_271
timestamp 1693479267
transform -1 0 4044 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_545
timestamp 1693479267
transform 1 0 4044 0 1 905
box -2 -3 34 103
use FILL  FILL_9_7_0
timestamp 1693479267
transform -1 0 4084 0 1 905
box -2 -3 10 103
use FILL  FILL_9_7_1
timestamp 1693479267
transform -1 0 4092 0 1 905
box -2 -3 10 103
use NAND2X1  NAND2X1_515
timestamp 1693479267
transform -1 0 4116 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_566
timestamp 1693479267
transform 1 0 4116 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_52
timestamp 1693479267
transform -1 0 4180 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_116
timestamp 1693479267
transform 1 0 4180 0 1 905
box -2 -3 34 103
use INVX4  INVX4_6
timestamp 1693479267
transform -1 0 4236 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_546
timestamp 1693479267
transform 1 0 4236 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_498
timestamp 1693479267
transform 1 0 4268 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_547
timestamp 1693479267
transform -1 0 4324 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_273
timestamp 1693479267
transform 1 0 4324 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_567
timestamp 1693479267
transform 1 0 4348 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_131
timestamp 1693479267
transform 1 0 4380 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_110
timestamp 1693479267
transform -1 0 4444 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_124
timestamp 1693479267
transform 1 0 4444 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_544
timestamp 1693479267
transform -1 0 4508 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_247
timestamp 1693479267
transform -1 0 4532 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_250
timestamp 1693479267
transform -1 0 4556 0 1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_137
timestamp 1693479267
transform 1 0 4556 0 1 905
box -2 -3 34 103
use FILL  FILL_10_1
timestamp 1693479267
transform 1 0 4588 0 1 905
box -2 -3 10 103
use FILL  FILL_10_2
timestamp 1693479267
transform 1 0 4596 0 1 905
box -2 -3 10 103
use BUFX2  BUFX2_22
timestamp 1693479267
transform -1 0 28 0 -1 1105
box -2 -3 26 103
use BUFX2  BUFX2_59
timestamp 1693479267
transform -1 0 52 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_179
timestamp 1693479267
transform -1 0 148 0 -1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_492
timestamp 1693479267
transform -1 0 244 0 -1 1105
box -2 -3 98 103
use AOI21X1  AOI21X1_218
timestamp 1693479267
transform 1 0 244 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_848
timestamp 1693479267
transform -1 0 308 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_849
timestamp 1693479267
transform 1 0 308 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_181
timestamp 1693479267
transform -1 0 372 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_47
timestamp 1693479267
transform -1 0 404 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_673
timestamp 1693479267
transform -1 0 428 0 -1 1105
box -2 -3 26 103
use BUFX4  BUFX4_199
timestamp 1693479267
transform 1 0 428 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_483
timestamp 1693479267
transform 1 0 460 0 -1 1105
box -2 -3 18 103
use FILL  FILL_10_0_0
timestamp 1693479267
transform 1 0 476 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_0_1
timestamp 1693479267
transform 1 0 484 0 -1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_460
timestamp 1693479267
transform 1 0 492 0 -1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_459
timestamp 1693479267
transform 1 0 588 0 -1 1105
box -2 -3 98 103
use NAND3X1  NAND3X1_46
timestamp 1693479267
transform 1 0 684 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_274
timestamp 1693479267
transform 1 0 716 0 -1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_273
timestamp 1693479267
transform 1 0 812 0 -1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_153
timestamp 1693479267
transform 1 0 908 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_256
timestamp 1693479267
transform -1 0 964 0 -1 1105
box -2 -3 34 103
use BUFX4  BUFX4_3
timestamp 1693479267
transform -1 0 996 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_1_0
timestamp 1693479267
transform 1 0 996 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_1_1
timestamp 1693479267
transform 1 0 1004 0 -1 1105
box -2 -3 10 103
use AND2X2  AND2X2_18
timestamp 1693479267
transform 1 0 1012 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_177
timestamp 1693479267
transform -1 0 1068 0 -1 1105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_14
timestamp 1693479267
transform 1 0 1068 0 -1 1105
box -2 -3 58 103
use AOI21X1  AOI21X1_29
timestamp 1693479267
transform -1 0 1156 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_248
timestamp 1693479267
transform 1 0 1156 0 -1 1105
box -2 -3 18 103
use INVX1  INVX1_261
timestamp 1693479267
transform 1 0 1172 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_238
timestamp 1693479267
transform 1 0 1188 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_241
timestamp 1693479267
transform 1 0 1220 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_252
timestamp 1693479267
transform -1 0 1268 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_240
timestamp 1693479267
transform 1 0 1268 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_134
timestamp 1693479267
transform -1 0 1324 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_13
timestamp 1693479267
transform -1 0 1356 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_245
timestamp 1693479267
transform 1 0 1356 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_236
timestamp 1693479267
transform -1 0 1404 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_237
timestamp 1693479267
transform 1 0 1404 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_81
timestamp 1693479267
transform 1 0 1436 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_11
timestamp 1693479267
transform 1 0 1468 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_246
timestamp 1693479267
transform -1 0 1516 0 -1 1105
box -2 -3 18 103
use FILL  FILL_10_2_0
timestamp 1693479267
transform 1 0 1516 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_2_1
timestamp 1693479267
transform 1 0 1524 0 -1 1105
box -2 -3 10 103
use AOI22X1  AOI22X1_43
timestamp 1693479267
transform 1 0 1532 0 -1 1105
box -2 -3 42 103
use BUFX4  BUFX4_150
timestamp 1693479267
transform -1 0 1604 0 -1 1105
box -2 -3 34 103
use AOI22X1  AOI22X1_44
timestamp 1693479267
transform 1 0 1604 0 -1 1105
box -2 -3 42 103
use MUX2X1  MUX2X1_1
timestamp 1693479267
transform -1 0 1692 0 -1 1105
box -2 -3 50 103
use AND2X2  AND2X2_62
timestamp 1693479267
transform -1 0 1724 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_571
timestamp 1693479267
transform -1 0 1748 0 -1 1105
box -2 -3 26 103
use INVX1  INVX1_413
timestamp 1693479267
transform 1 0 1748 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_711
timestamp 1693479267
transform -1 0 1796 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_409
timestamp 1693479267
transform 1 0 1796 0 -1 1105
box -2 -3 18 103
use NOR2X1  NOR2X1_324
timestamp 1693479267
transform 1 0 1812 0 -1 1105
box -2 -3 26 103
use NAND3X1  NAND3X1_89
timestamp 1693479267
transform -1 0 1868 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_351
timestamp 1693479267
transform 1 0 1868 0 -1 1105
box -2 -3 18 103
use AOI21X1  AOI21X1_156
timestamp 1693479267
transform 1 0 1884 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_405
timestamp 1693479267
transform -1 0 1932 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_708
timestamp 1693479267
transform 1 0 1932 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_185
timestamp 1693479267
transform -1 0 1996 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_342
timestamp 1693479267
transform -1 0 2020 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_321
timestamp 1693479267
transform 1 0 2020 0 -1 1105
box -2 -3 26 103
use FILL  FILL_10_3_0
timestamp 1693479267
transform -1 0 2052 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_3_1
timestamp 1693479267
transform -1 0 2060 0 -1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_626
timestamp 1693479267
transform -1 0 2092 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_322
timestamp 1693479267
transform -1 0 2116 0 -1 1105
box -2 -3 26 103
use BUFX4  BUFX4_154
timestamp 1693479267
transform -1 0 2148 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_62
timestamp 1693479267
transform 1 0 2148 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_48
timestamp 1693479267
transform 1 0 2180 0 -1 1105
box -2 -3 34 103
use AOI22X1  AOI22X1_79
timestamp 1693479267
transform -1 0 2252 0 -1 1105
box -2 -3 42 103
use OAI21X1  OAI21X1_427
timestamp 1693479267
transform 1 0 2252 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_425
timestamp 1693479267
transform 1 0 2284 0 -1 1105
box -2 -3 34 103
use AOI22X1  AOI22X1_78
timestamp 1693479267
transform 1 0 2316 0 -1 1105
box -2 -3 42 103
use NOR2X1  NOR2X1_210
timestamp 1693479267
transform 1 0 2356 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_429
timestamp 1693479267
transform 1 0 2380 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_318
timestamp 1693479267
transform 1 0 2412 0 -1 1105
box -2 -3 34 103
use NOR3X1  NOR3X1_57
timestamp 1693479267
transform -1 0 2508 0 -1 1105
box -2 -3 66 103
use NAND2X1  NAND2X1_392
timestamp 1693479267
transform -1 0 2532 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_376
timestamp 1693479267
transform 1 0 2532 0 -1 1105
box -2 -3 26 103
use FILL  FILL_10_4_0
timestamp 1693479267
transform 1 0 2556 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_4_1
timestamp 1693479267
transform 1 0 2564 0 -1 1105
box -2 -3 10 103
use NAND2X1  NAND2X1_363
timestamp 1693479267
transform 1 0 2572 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_618
timestamp 1693479267
transform -1 0 2628 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_400
timestamp 1693479267
transform -1 0 2644 0 -1 1105
box -2 -3 18 103
use AOI21X1  AOI21X1_66
timestamp 1693479267
transform 1 0 2644 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_414
timestamp 1693479267
transform 1 0 2676 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_394
timestamp 1693479267
transform -1 0 2724 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_310
timestamp 1693479267
transform -1 0 2748 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_615
timestamp 1693479267
transform -1 0 2780 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_543
timestamp 1693479267
transform 1 0 2780 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_209
timestamp 1693479267
transform 1 0 2804 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_182
timestamp 1693479267
transform 1 0 2828 0 -1 1105
box -2 -3 26 103
use NAND3X1  NAND3X1_105
timestamp 1693479267
transform -1 0 2884 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_409
timestamp 1693479267
transform 1 0 2884 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_165
timestamp 1693479267
transform -1 0 2940 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_382
timestamp 1693479267
transform -1 0 2956 0 -1 1105
box -2 -3 18 103
use NAND3X1  NAND3X1_118
timestamp 1693479267
transform -1 0 2988 0 -1 1105
box -2 -3 34 103
use AOI22X1  AOI22X1_87
timestamp 1693479267
transform 1 0 2988 0 -1 1105
box -2 -3 42 103
use INVX2  INVX2_65
timestamp 1693479267
transform 1 0 3028 0 -1 1105
box -2 -3 18 103
use FILL  FILL_10_5_0
timestamp 1693479267
transform 1 0 3044 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_5_1
timestamp 1693479267
transform 1 0 3052 0 -1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_482
timestamp 1693479267
transform 1 0 3060 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_239
timestamp 1693479267
transform -1 0 3116 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_411
timestamp 1693479267
transform 1 0 3116 0 -1 1105
box -2 -3 34 103
use OAI22X1  OAI22X1_14
timestamp 1693479267
transform 1 0 3148 0 -1 1105
box -2 -3 42 103
use OAI21X1  OAI21X1_367
timestamp 1693479267
transform 1 0 3188 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_366
timestamp 1693479267
transform -1 0 3252 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_567
timestamp 1693479267
transform 1 0 3252 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_237
timestamp 1693479267
transform 1 0 3276 0 -1 1105
box -2 -3 26 103
use INVX1  INVX1_385
timestamp 1693479267
transform -1 0 3316 0 -1 1105
box -2 -3 18 103
use NAND3X1  NAND3X1_152
timestamp 1693479267
transform -1 0 3348 0 -1 1105
box -2 -3 34 103
use AND2X2  AND2X2_60
timestamp 1693479267
transform 1 0 3348 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_687
timestamp 1693479267
transform 1 0 3380 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_227
timestamp 1693479267
transform 1 0 3412 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_459
timestamp 1693479267
transform 1 0 3436 0 -1 1105
box -2 -3 26 103
use BUFX4  BUFX4_176
timestamp 1693479267
transform -1 0 3492 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_379
timestamp 1693479267
transform -1 0 3508 0 -1 1105
box -2 -3 18 103
use NOR2X1  NOR2X1_272
timestamp 1693479267
transform -1 0 3532 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_149
timestamp 1693479267
transform 1 0 3532 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_6_0
timestamp 1693479267
transform -1 0 3572 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_6_1
timestamp 1693479267
transform -1 0 3580 0 -1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_663
timestamp 1693479267
transform -1 0 3612 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_327
timestamp 1693479267
transform 1 0 3612 0 -1 1105
box -2 -3 26 103
use OAI22X1  OAI22X1_16
timestamp 1693479267
transform 1 0 3636 0 -1 1105
box -2 -3 42 103
use NAND2X1  NAND2X1_572
timestamp 1693479267
transform -1 0 3700 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_446
timestamp 1693479267
transform -1 0 3724 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_240
timestamp 1693479267
transform 1 0 3724 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_516
timestamp 1693479267
transform 1 0 3748 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_686
timestamp 1693479267
transform 1 0 3780 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_172
timestamp 1693479267
transform -1 0 3844 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_428
timestamp 1693479267
transform -1 0 3868 0 -1 1105
box -2 -3 26 103
use OAI22X1  OAI22X1_28
timestamp 1693479267
transform -1 0 3908 0 -1 1105
box -2 -3 42 103
use OAI21X1  OAI21X1_558
timestamp 1693479267
transform 1 0 3908 0 -1 1105
box -2 -3 34 103
use INVX2  INVX2_55
timestamp 1693479267
transform -1 0 3956 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_702
timestamp 1693479267
transform 1 0 3956 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_338
timestamp 1693479267
transform 1 0 3988 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_703
timestamp 1693479267
transform 1 0 4012 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_340
timestamp 1693479267
transform -1 0 4068 0 -1 1105
box -2 -3 26 103
use FILL  FILL_10_7_0
timestamp 1693479267
transform -1 0 4076 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_7_1
timestamp 1693479267
transform -1 0 4084 0 -1 1105
box -2 -3 10 103
use AOI21X1  AOI21X1_182
timestamp 1693479267
transform -1 0 4116 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_561
timestamp 1693479267
transform -1 0 4140 0 -1 1105
box -2 -3 26 103
use INVX1  INVX1_387
timestamp 1693479267
transform 1 0 4140 0 -1 1105
box -2 -3 18 103
use OR2X2  OR2X2_29
timestamp 1693479267
transform 1 0 4156 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_121
timestamp 1693479267
transform -1 0 4220 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_476
timestamp 1693479267
transform 1 0 4220 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_343
timestamp 1693479267
transform -1 0 4268 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_115
timestamp 1693479267
transform 1 0 4268 0 -1 1105
box -2 -3 34 103
use OAI22X1  OAI22X1_35
timestamp 1693479267
transform 1 0 4300 0 -1 1105
box -2 -3 42 103
use AND2X2  AND2X2_45
timestamp 1693479267
transform 1 0 4340 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_134
timestamp 1693479267
transform -1 0 4404 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_278
timestamp 1693479267
transform -1 0 4428 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_559
timestamp 1693479267
transform -1 0 4460 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_279
timestamp 1693479267
transform -1 0 4484 0 -1 1105
box -2 -3 26 103
use OAI22X1  OAI22X1_30
timestamp 1693479267
transform 1 0 4484 0 -1 1105
box -2 -3 42 103
use NAND2X1  NAND2X1_516
timestamp 1693479267
transform -1 0 4548 0 -1 1105
box -2 -3 26 103
use INVX4  INVX4_9
timestamp 1693479267
transform 1 0 4548 0 -1 1105
box -2 -3 26 103
use AND2X2  AND2X2_72
timestamp 1693479267
transform -1 0 4604 0 -1 1105
box -2 -3 34 103
use BUFX2  BUFX2_58
timestamp 1693479267
transform -1 0 28 0 1 1105
box -2 -3 26 103
use BUFX2  BUFX2_19
timestamp 1693479267
transform -1 0 52 0 1 1105
box -2 -3 26 103
use BUFX2  BUFX2_60
timestamp 1693479267
transform -1 0 76 0 1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_176
timestamp 1693479267
transform -1 0 172 0 1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_493
timestamp 1693479267
transform -1 0 268 0 1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_676
timestamp 1693479267
transform 1 0 268 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_670
timestamp 1693479267
transform -1 0 316 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_675
timestamp 1693479267
transform 1 0 316 0 1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_491
timestamp 1693479267
transform -1 0 436 0 1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_851
timestamp 1693479267
transform 1 0 436 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_850
timestamp 1693479267
transform 1 0 468 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_0_0
timestamp 1693479267
transform -1 0 508 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_0_1
timestamp 1693479267
transform -1 0 516 0 1 1105
box -2 -3 10 103
use INVX1  INVX1_484
timestamp 1693479267
transform -1 0 532 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_182
timestamp 1693479267
transform 1 0 532 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_852
timestamp 1693479267
transform 1 0 564 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_677
timestamp 1693479267
transform -1 0 620 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_847
timestamp 1693479267
transform 1 0 620 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_641
timestamp 1693479267
transform -1 0 676 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_674
timestamp 1693479267
transform 1 0 676 0 1 1105
box -2 -3 26 103
use NAND3X1  NAND3X1_44
timestamp 1693479267
transform 1 0 700 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_48
timestamp 1693479267
transform -1 0 764 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_113
timestamp 1693479267
transform -1 0 796 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_461
timestamp 1693479267
transform 1 0 796 0 1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_275
timestamp 1693479267
transform 1 0 892 0 1 1105
box -2 -3 98 103
use AND2X2  AND2X2_14
timestamp 1693479267
transform -1 0 1020 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_1_0
timestamp 1693479267
transform -1 0 1028 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_1_1
timestamp 1693479267
transform -1 0 1036 0 1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_263
timestamp 1693479267
transform -1 0 1068 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_259
timestamp 1693479267
transform -1 0 1100 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_159
timestamp 1693479267
transform -1 0 1124 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_276
timestamp 1693479267
transform -1 0 1156 0 1 1105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_39
timestamp 1693479267
transform 1 0 1156 0 1 1105
box -2 -3 58 103
use AOI21X1  AOI21X1_26
timestamp 1693479267
transform -1 0 1244 0 1 1105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_12
timestamp 1693479267
transform 1 0 1244 0 1 1105
box -2 -3 58 103
use AOI21X1  AOI21X1_25
timestamp 1693479267
transform -1 0 1332 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_138
timestamp 1693479267
transform 1 0 1332 0 1 1105
box -2 -3 26 103
use INVX1  INVX1_244
timestamp 1693479267
transform 1 0 1356 0 1 1105
box -2 -3 18 103
use AOI21X1  AOI21X1_10
timestamp 1693479267
transform -1 0 1404 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_240
timestamp 1693479267
transform 1 0 1404 0 1 1105
box -2 -3 18 103
use NOR2X1  NOR2X1_29
timestamp 1693479267
transform -1 0 1444 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_233
timestamp 1693479267
transform 1 0 1444 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_131
timestamp 1693479267
transform -1 0 1500 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_137
timestamp 1693479267
transform -1 0 1524 0 1 1105
box -2 -3 26 103
use FILL  FILL_11_2_0
timestamp 1693479267
transform 1 0 1524 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_2_1
timestamp 1693479267
transform 1 0 1532 0 1 1105
box -2 -3 10 103
use NAND2X1  NAND2X1_130
timestamp 1693479267
transform 1 0 1540 0 1 1105
box -2 -3 26 103
use NOR3X1  NOR3X1_50
timestamp 1693479267
transform -1 0 1628 0 1 1105
box -2 -3 66 103
use INVX1  INVX1_242
timestamp 1693479267
transform -1 0 1644 0 1 1105
box -2 -3 18 103
use NAND2X1  NAND2X1_132
timestamp 1693479267
transform -1 0 1668 0 1 1105
box -2 -3 26 103
use AOI22X1  AOI22X1_56
timestamp 1693479267
transform -1 0 1708 0 1 1105
box -2 -3 42 103
use BUFX4  BUFX4_147
timestamp 1693479267
transform -1 0 1740 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_231
timestamp 1693479267
transform 1 0 1740 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_222
timestamp 1693479267
transform -1 0 1796 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_297
timestamp 1693479267
transform -1 0 1828 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_323
timestamp 1693479267
transform -1 0 1844 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_305
timestamp 1693479267
transform 1 0 1844 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_328
timestamp 1693479267
transform -1 0 1892 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_659
timestamp 1693479267
transform -1 0 1924 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_661
timestamp 1693479267
transform 1 0 1924 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_166
timestamp 1693479267
transform 1 0 1956 0 1 1105
box -2 -3 34 103
use INVX4  INVX4_10
timestamp 1693479267
transform 1 0 1988 0 1 1105
box -2 -3 26 103
use NAND3X1  NAND3X1_160
timestamp 1693479267
transform 1 0 2012 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_3_0
timestamp 1693479267
transform 1 0 2044 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_3_1
timestamp 1693479267
transform 1 0 2052 0 1 1105
box -2 -3 10 103
use NOR2X1  NOR2X1_326
timestamp 1693479267
transform 1 0 2060 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_325
timestamp 1693479267
transform -1 0 2108 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_680
timestamp 1693479267
transform 1 0 2108 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_216
timestamp 1693479267
transform 1 0 2140 0 1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_176
timestamp 1693479267
transform -1 0 2196 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_570
timestamp 1693479267
transform 1 0 2196 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_660
timestamp 1693479267
transform -1 0 2252 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_410
timestamp 1693479267
transform 1 0 2252 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_694
timestamp 1693479267
transform -1 0 2300 0 1 1105
box -2 -3 34 103
use AOI22X1  AOI22X1_102
timestamp 1693479267
transform 1 0 2300 0 1 1105
box -2 -3 42 103
use OAI21X1  OAI21X1_666
timestamp 1693479267
transform 1 0 2340 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_428
timestamp 1693479267
transform 1 0 2372 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_155
timestamp 1693479267
transform -1 0 2436 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_274
timestamp 1693479267
transform -1 0 2460 0 1 1105
box -2 -3 26 103
use NAND3X1  NAND3X1_116
timestamp 1693479267
transform 1 0 2460 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_231
timestamp 1693479267
transform -1 0 2516 0 1 1105
box -2 -3 26 103
use INVX1  INVX1_370
timestamp 1693479267
transform -1 0 2532 0 1 1105
box -2 -3 18 103
use FILL  FILL_11_4_0
timestamp 1693479267
transform 1 0 2532 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_4_1
timestamp 1693479267
transform 1 0 2540 0 1 1105
box -2 -3 10 103
use AOI21X1  AOI21X1_63
timestamp 1693479267
transform 1 0 2548 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_213
timestamp 1693479267
transform -1 0 2604 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_311
timestamp 1693479267
transform -1 0 2628 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_271
timestamp 1693479267
transform -1 0 2652 0 1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_65
timestamp 1693479267
transform -1 0 2684 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_372
timestamp 1693479267
transform -1 0 2700 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_616
timestamp 1693479267
transform 1 0 2700 0 1 1105
box -2 -3 34 103
use OR2X2  OR2X2_36
timestamp 1693479267
transform -1 0 2764 0 1 1105
box -2 -3 34 103
use NOR3X1  NOR3X1_58
timestamp 1693479267
transform 1 0 2764 0 1 1105
box -2 -3 66 103
use AND2X2  AND2X2_49
timestamp 1693479267
transform -1 0 2860 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_623
timestamp 1693479267
transform -1 0 2892 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_357
timestamp 1693479267
transform -1 0 2908 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_368
timestamp 1693479267
transform -1 0 2940 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_173
timestamp 1693479267
transform -1 0 2964 0 1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_150
timestamp 1693479267
transform 1 0 2964 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_456
timestamp 1693479267
transform 1 0 2996 0 1 1105
box -2 -3 26 103
use NAND3X1  NAND3X1_112
timestamp 1693479267
transform -1 0 3052 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_5_0
timestamp 1693479267
transform 1 0 3052 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_5_1
timestamp 1693479267
transform 1 0 3060 0 1 1105
box -2 -3 10 103
use INVX2  INVX2_54
timestamp 1693479267
transform 1 0 3068 0 1 1105
box -2 -3 18 103
use OAI22X1  OAI22X1_19
timestamp 1693479267
transform 1 0 3084 0 1 1105
box -2 -3 42 103
use BUFX4  BUFX4_126
timestamp 1693479267
transform -1 0 3156 0 1 1105
box -2 -3 34 103
use INVX4  INVX4_5
timestamp 1693479267
transform 1 0 3156 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_467
timestamp 1693479267
transform -1 0 3204 0 1 1105
box -2 -3 26 103
use BUFX4  BUFX4_82
timestamp 1693479267
transform -1 0 3236 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_397
timestamp 1693479267
transform -1 0 3260 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_489
timestamp 1693479267
transform -1 0 3292 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_690
timestamp 1693479267
transform -1 0 3324 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_173
timestamp 1693479267
transform -1 0 3356 0 1 1105
box -2 -3 34 103
use NOR3X1  NOR3X1_61
timestamp 1693479267
transform 1 0 3356 0 1 1105
box -2 -3 66 103
use OAI21X1  OAI21X1_483
timestamp 1693479267
transform -1 0 3452 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_488
timestamp 1693479267
transform -1 0 3484 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_124
timestamp 1693479267
transform -1 0 3516 0 1 1105
box -2 -3 34 103
use OR2X2  OR2X2_27
timestamp 1693479267
transform -1 0 3548 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_624
timestamp 1693479267
transform -1 0 3580 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_6_0
timestamp 1693479267
transform -1 0 3588 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_6_1
timestamp 1693479267
transform -1 0 3596 0 1 1105
box -2 -3 10 103
use OR2X2  OR2X2_26
timestamp 1693479267
transform -1 0 3628 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_389
timestamp 1693479267
transform 1 0 3628 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_534
timestamp 1693479267
transform 1 0 3644 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_337
timestamp 1693479267
transform -1 0 3700 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_491
timestamp 1693479267
transform -1 0 3724 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_701
timestamp 1693479267
transform 1 0 3724 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_57
timestamp 1693479267
transform -1 0 3788 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_622
timestamp 1693479267
transform -1 0 3820 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_315
timestamp 1693479267
transform 1 0 3820 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_559
timestamp 1693479267
transform 1 0 3844 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_334
timestamp 1693479267
transform -1 0 3892 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_688
timestamp 1693479267
transform 1 0 3892 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_508
timestamp 1693479267
transform -1 0 3948 0 1 1105
box -2 -3 26 103
use AND2X2  AND2X2_61
timestamp 1693479267
transform -1 0 3980 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_125
timestamp 1693479267
transform -1 0 4012 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_339
timestamp 1693479267
transform -1 0 4036 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_704
timestamp 1693479267
transform 1 0 4036 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_7_0
timestamp 1693479267
transform -1 0 4076 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_7_1
timestamp 1693479267
transform -1 0 4084 0 1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_705
timestamp 1693479267
transform -1 0 4116 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_163
timestamp 1693479267
transform 1 0 4116 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_447
timestamp 1693479267
transform -1 0 4172 0 1 1105
box -2 -3 26 103
use OAI22X1  OAI22X1_27
timestamp 1693479267
transform 1 0 4172 0 1 1105
box -2 -3 42 103
use NAND2X1  NAND2X1_475
timestamp 1693479267
transform -1 0 4236 0 1 1105
box -2 -3 26 103
use INVX1  INVX1_388
timestamp 1693479267
transform 1 0 4236 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_524
timestamp 1693479267
transform 1 0 4252 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_523
timestamp 1693479267
transform 1 0 4284 0 1 1105
box -2 -3 34 103
use AOI22X1  AOI22X1_91
timestamp 1693479267
transform -1 0 4356 0 1 1105
box -2 -3 42 103
use BUFX4  BUFX4_53
timestamp 1693479267
transform 1 0 4356 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_529
timestamp 1693479267
transform -1 0 4412 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_517
timestamp 1693479267
transform 1 0 4412 0 1 1105
box -2 -3 26 103
use OAI22X1  OAI22X1_33
timestamp 1693479267
transform -1 0 4476 0 1 1105
box -2 -3 42 103
use NAND2X1  NAND2X1_361
timestamp 1693479267
transform -1 0 4500 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_779
timestamp 1693479267
transform 1 0 4500 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_368
timestamp 1693479267
transform -1 0 4556 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_778
timestamp 1693479267
transform -1 0 4588 0 1 1105
box -2 -3 34 103
use FILL  FILL_12_1
timestamp 1693479267
transform 1 0 4588 0 1 1105
box -2 -3 10 103
use FILL  FILL_12_2
timestamp 1693479267
transform 1 0 4596 0 1 1105
box -2 -3 10 103
use BUFX2  BUFX2_4
timestamp 1693479267
transform -1 0 28 0 -1 1305
box -2 -3 26 103
use BUFX2  BUFX2_21
timestamp 1693479267
transform -1 0 52 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_178
timestamp 1693479267
transform -1 0 148 0 -1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_681
timestamp 1693479267
transform 1 0 148 0 -1 1305
box -2 -3 26 103
use AND2X2  AND2X2_78
timestamp 1693479267
transform 1 0 172 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_393
timestamp 1693479267
transform -1 0 228 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_672
timestamp 1693479267
transform 1 0 228 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_391
timestamp 1693479267
transform -1 0 276 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_219
timestamp 1693479267
transform 1 0 276 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_392
timestamp 1693479267
transform -1 0 332 0 -1 1305
box -2 -3 26 103
use OR2X2  OR2X2_48
timestamp 1693479267
transform 1 0 332 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_485
timestamp 1693479267
transform 1 0 364 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_853
timestamp 1693479267
transform 1 0 380 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_854
timestamp 1693479267
transform 1 0 412 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_16
timestamp 1693479267
transform 1 0 444 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_198
timestamp 1693479267
transform 1 0 476 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_0_0
timestamp 1693479267
transform -1 0 516 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_0_1
timestamp 1693479267
transform -1 0 524 0 -1 1305
box -2 -3 10 103
use NAND3X1  NAND3X1_49
timestamp 1693479267
transform -1 0 556 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_45
timestamp 1693479267
transform 1 0 556 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_180
timestamp 1693479267
transform 1 0 588 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_161
timestamp 1693479267
transform -1 0 716 0 -1 1305
box -2 -3 98 103
use CLKBUF1  CLKBUF1_52
timestamp 1693479267
transform -1 0 788 0 -1 1305
box -2 -3 74 103
use XNOR2X1  XNOR2X1_40
timestamp 1693479267
transform 1 0 788 0 -1 1305
box -2 -3 58 103
use AOI21X1  AOI21X1_28
timestamp 1693479267
transform 1 0 844 0 -1 1305
box -2 -3 34 103
use AND2X2  AND2X2_15
timestamp 1693479267
transform -1 0 908 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_166
timestamp 1693479267
transform -1 0 932 0 -1 1305
box -2 -3 26 103
use INVX1  INVX1_270
timestamp 1693479267
transform -1 0 948 0 -1 1305
box -2 -3 18 103
use XOR2X1  XOR2X1_4
timestamp 1693479267
transform 1 0 948 0 -1 1305
box -2 -3 58 103
use FILL  FILL_12_1_0
timestamp 1693479267
transform -1 0 1012 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_1_1
timestamp 1693479267
transform -1 0 1020 0 -1 1305
box -2 -3 10 103
use NOR2X1  NOR2X1_44
timestamp 1693479267
transform -1 0 1044 0 -1 1305
box -2 -3 26 103
use OR2X2  OR2X2_11
timestamp 1693479267
transform 1 0 1044 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_27
timestamp 1693479267
transform -1 0 1108 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_265
timestamp 1693479267
transform -1 0 1124 0 -1 1305
box -2 -3 18 103
use XNOR2X1  XNOR2X1_16
timestamp 1693479267
transform -1 0 1180 0 -1 1305
box -2 -3 58 103
use NAND2X1  NAND2X1_139
timestamp 1693479267
transform -1 0 1204 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_129
timestamp 1693479267
transform 1 0 1204 0 -1 1305
box -2 -3 26 103
use XNOR2X1  XNOR2X1_38
timestamp 1693479267
transform 1 0 1228 0 -1 1305
box -2 -3 58 103
use INVX1  INVX1_243
timestamp 1693479267
transform 1 0 1284 0 -1 1305
box -2 -3 18 103
use NAND3X1  NAND3X1_80
timestamp 1693479267
transform 1 0 1300 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_14
timestamp 1693479267
transform -1 0 1364 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_235
timestamp 1693479267
transform 1 0 1364 0 -1 1305
box -2 -3 34 103
use AOI22X1  AOI22X1_45
timestamp 1693479267
transform 1 0 1396 0 -1 1305
box -2 -3 42 103
use NAND2X1  NAND2X1_128
timestamp 1693479267
transform -1 0 1460 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_136
timestamp 1693479267
transform 1 0 1460 0 -1 1305
box -2 -3 26 103
use INVX1  INVX1_249
timestamp 1693479267
transform 1 0 1484 0 -1 1305
box -2 -3 18 103
use NAND3X1  NAND3X1_82
timestamp 1693479267
transform 1 0 1500 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_2_0
timestamp 1693479267
transform -1 0 1540 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_2_1
timestamp 1693479267
transform -1 0 1548 0 -1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_234
timestamp 1693479267
transform -1 0 1580 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_135
timestamp 1693479267
transform -1 0 1604 0 -1 1305
box -2 -3 26 103
use AOI22X1  AOI22X1_46
timestamp 1693479267
transform -1 0 1644 0 -1 1305
box -2 -3 42 103
use OAI21X1  OAI21X1_667
timestamp 1693479267
transform -1 0 1676 0 -1 1305
box -2 -3 34 103
use AND2X2  AND2X2_54
timestamp 1693479267
transform -1 0 1708 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_658
timestamp 1693479267
transform 1 0 1708 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_679
timestamp 1693479267
transform -1 0 1772 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_304
timestamp 1693479267
transform 1 0 1772 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_411
timestamp 1693479267
transform 1 0 1804 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_647
timestamp 1693479267
transform -1 0 1852 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_159
timestamp 1693479267
transform 1 0 1852 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_657
timestamp 1693479267
transform 1 0 1884 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_221
timestamp 1693479267
transform 1 0 1916 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_220
timestamp 1693479267
transform 1 0 1940 0 -1 1305
box -2 -3 26 103
use AND2X2  AND2X2_51
timestamp 1693479267
transform 1 0 1964 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_417
timestamp 1693479267
transform -1 0 2012 0 -1 1305
box -2 -3 18 103
use AOI21X1  AOI21X1_184
timestamp 1693479267
transform 1 0 2012 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_3_0
timestamp 1693479267
transform -1 0 2052 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_3_1
timestamp 1693479267
transform -1 0 2060 0 -1 1305
box -2 -3 10 103
use INVX1  INVX1_418
timestamp 1693479267
transform -1 0 2076 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_655
timestamp 1693479267
transform -1 0 2108 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_408
timestamp 1693479267
transform 1 0 2108 0 -1 1305
box -2 -3 18 103
use INVX2  INVX2_69
timestamp 1693479267
transform 1 0 2124 0 -1 1305
box -2 -3 18 103
use AOI21X1  AOI21X1_167
timestamp 1693479267
transform -1 0 2172 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_554
timestamp 1693479267
transform 1 0 2172 0 -1 1305
box -2 -3 26 103
use NAND3X1  NAND3X1_150
timestamp 1693479267
transform 1 0 2196 0 -1 1305
box -2 -3 34 103
use AND2X2  AND2X2_22
timestamp 1693479267
transform -1 0 2260 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_393
timestamp 1693479267
transform -1 0 2284 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_212
timestamp 1693479267
transform 1 0 2284 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_426
timestamp 1693479267
transform 1 0 2308 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_142
timestamp 1693479267
transform 1 0 2340 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_356
timestamp 1693479267
transform 1 0 2364 0 -1 1305
box -2 -3 26 103
use INVX1  INVX1_369
timestamp 1693479267
transform 1 0 2388 0 -1 1305
box -2 -3 18 103
use NOR2X1  NOR2X1_195
timestamp 1693479267
transform -1 0 2428 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_196
timestamp 1693479267
transform -1 0 2452 0 -1 1305
box -2 -3 26 103
use AOI22X1  AOI22X1_76
timestamp 1693479267
transform 1 0 2452 0 -1 1305
box -2 -3 42 103
use NAND2X1  NAND2X1_377
timestamp 1693479267
transform 1 0 2492 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_391
timestamp 1693479267
transform -1 0 2540 0 -1 1305
box -2 -3 26 103
use FILL  FILL_12_4_0
timestamp 1693479267
transform 1 0 2540 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_4_1
timestamp 1693479267
transform 1 0 2548 0 -1 1305
box -2 -3 10 103
use NAND2X1  NAND2X1_357
timestamp 1693479267
transform 1 0 2556 0 -1 1305
box -2 -3 26 103
use INVX8  INVX8_6
timestamp 1693479267
transform -1 0 2620 0 -1 1305
box -2 -3 42 103
use AOI21X1  AOI21X1_162
timestamp 1693479267
transform -1 0 2652 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_78
timestamp 1693479267
transform 1 0 2652 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_194
timestamp 1693479267
transform 1 0 2684 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_407
timestamp 1693479267
transform -1 0 2740 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_59
timestamp 1693479267
transform 1 0 2740 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_54
timestamp 1693479267
transform -1 0 2804 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_370
timestamp 1693479267
transform 1 0 2804 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_57
timestamp 1693479267
transform 1 0 2836 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_433
timestamp 1693479267
transform 1 0 2868 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_369
timestamp 1693479267
transform 1 0 2892 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_678
timestamp 1693479267
transform -1 0 2956 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_80
timestamp 1693479267
transform 1 0 2956 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_453
timestamp 1693479267
transform -1 0 3012 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_204
timestamp 1693479267
transform 1 0 3012 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_458
timestamp 1693479267
transform -1 0 3068 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_5_0
timestamp 1693479267
transform -1 0 3076 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_5_1
timestamp 1693479267
transform -1 0 3084 0 -1 1305
box -2 -3 10 103
use AND2X2  AND2X2_53
timestamp 1693479267
transform -1 0 3116 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_509
timestamp 1693479267
transform 1 0 3116 0 -1 1305
box -2 -3 26 103
use AND2X2  AND2X2_33
timestamp 1693479267
transform -1 0 3172 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_371
timestamp 1693479267
transform 1 0 3172 0 -1 1305
box -2 -3 18 103
use NOR3X1  NOR3X1_60
timestamp 1693479267
transform -1 0 3252 0 -1 1305
box -2 -3 66 103
use NAND2X1  NAND2X1_463
timestamp 1693479267
transform -1 0 3276 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_170
timestamp 1693479267
transform -1 0 3308 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_563
timestamp 1693479267
transform -1 0 3332 0 -1 1305
box -2 -3 26 103
use INVX8  INVX8_9
timestamp 1693479267
transform -1 0 3372 0 -1 1305
box -2 -3 42 103
use NOR2X1  NOR2X1_226
timestamp 1693479267
transform -1 0 3396 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_229
timestamp 1693479267
transform 1 0 3396 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_217
timestamp 1693479267
transform 1 0 3420 0 -1 1305
box -2 -3 26 103
use BUFX4  BUFX4_174
timestamp 1693479267
transform -1 0 3476 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_564
timestamp 1693479267
transform -1 0 3500 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_202
timestamp 1693479267
transform -1 0 3524 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_653
timestamp 1693479267
transform 1 0 3524 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_6_0
timestamp 1693479267
transform -1 0 3564 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_6_1
timestamp 1693479267
transform -1 0 3572 0 -1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_652
timestamp 1693479267
transform -1 0 3604 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_456
timestamp 1693479267
transform -1 0 3636 0 -1 1305
box -2 -3 34 103
use AND2X2  AND2X2_57
timestamp 1693479267
transform -1 0 3668 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_675
timestamp 1693479267
transform 1 0 3668 0 -1 1305
box -2 -3 34 103
use AND2X2  AND2X2_67
timestamp 1693479267
transform -1 0 3732 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_542
timestamp 1693479267
transform -1 0 3756 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_552
timestamp 1693479267
transform -1 0 3780 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_314
timestamp 1693479267
transform -1 0 3804 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_501
timestamp 1693479267
transform -1 0 3828 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_505
timestamp 1693479267
transform 1 0 3828 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_504
timestamp 1693479267
transform -1 0 3876 0 -1 1305
box -2 -3 26 103
use BUFX4  BUFX4_81
timestamp 1693479267
transform -1 0 3908 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_674
timestamp 1693479267
transform -1 0 3940 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_586
timestamp 1693479267
transform 1 0 3940 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_329
timestamp 1693479267
transform 1 0 3972 0 -1 1305
box -2 -3 26 103
use AND2X2  AND2X2_63
timestamp 1693479267
transform -1 0 4028 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_473
timestamp 1693479267
transform -1 0 4060 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_440
timestamp 1693479267
transform -1 0 4084 0 -1 1305
box -2 -3 26 103
use FILL  FILL_12_7_0
timestamp 1693479267
transform 1 0 4084 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_7_1
timestamp 1693479267
transform 1 0 4092 0 -1 1305
box -2 -3 10 103
use AND2X2  AND2X2_38
timestamp 1693479267
transform 1 0 4100 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_508
timestamp 1693479267
transform 1 0 4132 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_560
timestamp 1693479267
transform 1 0 4164 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_484
timestamp 1693479267
transform -1 0 4212 0 -1 1305
box -2 -3 26 103
use OR2X2  OR2X2_33
timestamp 1693479267
transform -1 0 4244 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_128
timestamp 1693479267
transform -1 0 4276 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_328
timestamp 1693479267
transform 1 0 4276 0 -1 1305
box -2 -3 26 103
use AOI22X1  AOI22X1_107
timestamp 1693479267
transform -1 0 4340 0 -1 1305
box -2 -3 42 103
use NAND2X1  NAND2X1_598
timestamp 1693479267
transform -1 0 4364 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_758
timestamp 1693479267
transform -1 0 4396 0 -1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_55
timestamp 1693479267
transform 1 0 4396 0 -1 1305
box -2 -3 50 103
use OAI21X1  OAI21X1_673
timestamp 1693479267
transform -1 0 4476 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_759
timestamp 1693479267
transform -1 0 4508 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_761
timestamp 1693479267
transform -1 0 4540 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_206
timestamp 1693479267
transform -1 0 4572 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_175
timestamp 1693479267
transform -1 0 4604 0 -1 1305
box -2 -3 34 103
use BUFX2  BUFX2_24
timestamp 1693479267
transform -1 0 28 0 1 1305
box -2 -3 26 103
use BUFX2  BUFX2_25
timestamp 1693479267
transform -1 0 52 0 1 1305
box -2 -3 26 103
use BUFX2  BUFX2_23
timestamp 1693479267
transform -1 0 76 0 1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_181
timestamp 1693479267
transform -1 0 172 0 1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_680
timestamp 1693479267
transform 1 0 172 0 1 1305
box -2 -3 26 103
use NAND3X1  NAND3X1_184
timestamp 1693479267
transform 1 0 196 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_182
timestamp 1693479267
transform -1 0 324 0 1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_855
timestamp 1693479267
transform 1 0 324 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_856
timestamp 1693479267
transform 1 0 356 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_679
timestamp 1693479267
transform -1 0 412 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_678
timestamp 1693479267
transform 1 0 412 0 1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_180
timestamp 1693479267
transform -1 0 532 0 1 1305
box -2 -3 98 103
use FILL  FILL_13_0_0
timestamp 1693479267
transform 1 0 532 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_0_1
timestamp 1693479267
transform 1 0 540 0 1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_184
timestamp 1693479267
transform 1 0 548 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_183
timestamp 1693479267
transform -1 0 612 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_494
timestamp 1693479267
transform -1 0 708 0 1 1305
box -2 -3 98 103
use NAND3X1  NAND3X1_51
timestamp 1693479267
transform -1 0 740 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_137
timestamp 1693479267
transform -1 0 772 0 1 1305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_27
timestamp 1693479267
transform 1 0 772 0 1 1305
box -2 -3 74 103
use XNOR2X1  XNOR2X1_41
timestamp 1693479267
transform 1 0 844 0 1 1305
box -2 -3 58 103
use INVX1  INVX1_272
timestamp 1693479267
transform 1 0 900 0 1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_264
timestamp 1693479267
transform 1 0 916 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_45
timestamp 1693479267
transform 1 0 948 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_178
timestamp 1693479267
transform -1 0 996 0 1 1305
box -2 -3 26 103
use FILL  FILL_13_1_0
timestamp 1693479267
transform 1 0 996 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_1_1
timestamp 1693479267
transform 1 0 1004 0 1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_265
timestamp 1693479267
transform 1 0 1012 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_33
timestamp 1693479267
transform -1 0 1076 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_262
timestamp 1693479267
transform 1 0 1076 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_50
timestamp 1693479267
transform -1 0 1132 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_268
timestamp 1693479267
transform -1 0 1164 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_269
timestamp 1693479267
transform -1 0 1180 0 1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_261
timestamp 1693479267
transform -1 0 1212 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_165
timestamp 1693479267
transform -1 0 1236 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_161
timestamp 1693479267
transform -1 0 1260 0 1 1305
box -2 -3 26 103
use OR2X2  OR2X2_10
timestamp 1693479267
transform -1 0 1292 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_160
timestamp 1693479267
transform -1 0 1316 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_42
timestamp 1693479267
transform 1 0 1316 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_156
timestamp 1693479267
transform -1 0 1364 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_122
timestamp 1693479267
transform 1 0 1364 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_127
timestamp 1693479267
transform -1 0 1412 0 1 1305
box -2 -3 26 103
use INVX1  INVX1_251
timestamp 1693479267
transform 1 0 1412 0 1 1305
box -2 -3 18 103
use NOR3X1  NOR3X1_52
timestamp 1693479267
transform 1 0 1428 0 1 1305
box -2 -3 66 103
use OAI21X1  OAI21X1_239
timestamp 1693479267
transform -1 0 1524 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_2_0
timestamp 1693479267
transform 1 0 1524 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_2_1
timestamp 1693479267
transform 1 0 1532 0 1 1305
box -2 -3 10 103
use AOI21X1  AOI21X1_9
timestamp 1693479267
transform 1 0 1540 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_241
timestamp 1693479267
transform -1 0 1588 0 1 1305
box -2 -3 18 103
use AOI21X1  AOI21X1_12
timestamp 1693479267
transform 1 0 1588 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_250
timestamp 1693479267
transform -1 0 1636 0 1 1305
box -2 -3 18 103
use BUFX4  BUFX4_232
timestamp 1693479267
transform -1 0 1668 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_296
timestamp 1693479267
transform 1 0 1668 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_219
timestamp 1693479267
transform 1 0 1700 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_555
timestamp 1693479267
transform 1 0 1724 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_102
timestamp 1693479267
transform 1 0 1748 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_101
timestamp 1693479267
transform -1 0 1796 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_235
timestamp 1693479267
transform -1 0 1820 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_668
timestamp 1693479267
transform 1 0 1820 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_151
timestamp 1693479267
transform -1 0 1884 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_643
timestamp 1693479267
transform 1 0 1884 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_406
timestamp 1693479267
transform 1 0 1916 0 1 1305
box -2 -3 18 103
use AOI21X1  AOI21X1_157
timestamp 1693479267
transform 1 0 1932 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_669
timestamp 1693479267
transform 1 0 1964 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_336
timestamp 1693479267
transform 1 0 1996 0 1 1305
box -2 -3 26 103
use FILL  FILL_13_3_0
timestamp 1693479267
transform 1 0 2020 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_3_1
timestamp 1693479267
transform 1 0 2028 0 1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_693
timestamp 1693479267
transform 1 0 2036 0 1 1305
box -2 -3 34 103
use INVX2  INVX2_31
timestamp 1693479267
transform -1 0 2084 0 1 1305
box -2 -3 18 103
use NAND2X1  NAND2X1_215
timestamp 1693479267
transform 1 0 2084 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_218
timestamp 1693479267
transform -1 0 2132 0 1 1305
box -2 -3 26 103
use INVX2  INVX2_32
timestamp 1693479267
transform -1 0 2148 0 1 1305
box -2 -3 18 103
use NAND3X1  NAND3X1_97
timestamp 1693479267
transform 1 0 2148 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_214
timestamp 1693479267
transform 1 0 2180 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_654
timestamp 1693479267
transform 1 0 2204 0 1 1305
box -2 -3 34 103
use AOI22X1  AOI22X1_77
timestamp 1693479267
transform 1 0 2236 0 1 1305
box -2 -3 42 103
use NOR2X1  NOR2X1_197
timestamp 1693479267
transform -1 0 2300 0 1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_69
timestamp 1693479267
transform -1 0 2332 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_273
timestamp 1693479267
transform -1 0 2356 0 1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_60
timestamp 1693479267
transform 1 0 2356 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_193
timestamp 1693479267
transform -1 0 2412 0 1 1305
box -2 -3 26 103
use OAI22X1  OAI22X1_13
timestamp 1693479267
transform -1 0 2452 0 1 1305
box -2 -3 42 103
use NAND3X1  NAND3X1_108
timestamp 1693479267
transform -1 0 2484 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_321
timestamp 1693479267
transform 1 0 2484 0 1 1305
box -2 -3 18 103
use NOR2X1  NOR2X1_184
timestamp 1693479267
transform -1 0 2524 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_161
timestamp 1693479267
transform -1 0 2548 0 1 1305
box -2 -3 26 103
use FILL  FILL_13_4_0
timestamp 1693479267
transform 1 0 2548 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_4_1
timestamp 1693479267
transform 1 0 2556 0 1 1305
box -2 -3 10 103
use NAND3X1  NAND3X1_109
timestamp 1693479267
transform 1 0 2564 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_200
timestamp 1693479267
transform 1 0 2596 0 1 1305
box -2 -3 26 103
use NAND3X1  NAND3X1_94
timestamp 1693479267
transform 1 0 2620 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_143
timestamp 1693479267
transform 1 0 2652 0 1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_171
timestamp 1693479267
transform -1 0 2708 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_298
timestamp 1693479267
transform -1 0 2732 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_359
timestamp 1693479267
transform -1 0 2756 0 1 1305
box -2 -3 26 103
use NAND3X1  NAND3X1_106
timestamp 1693479267
transform -1 0 2788 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_376
timestamp 1693479267
transform -1 0 2820 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_358
timestamp 1693479267
transform 1 0 2820 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_656
timestamp 1693479267
transform -1 0 2876 0 1 1305
box -2 -3 34 103
use NOR3X1  NOR3X1_59
timestamp 1693479267
transform -1 0 2940 0 1 1305
box -2 -3 66 103
use AOI21X1  AOI21X1_61
timestamp 1693479267
transform 1 0 2940 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_83
timestamp 1693479267
transform -1 0 3004 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_85
timestamp 1693479267
transform -1 0 3036 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_457
timestamp 1693479267
transform 1 0 3036 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_5_0
timestamp 1693479267
transform -1 0 3076 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_5_1
timestamp 1693479267
transform -1 0 3084 0 1 1305
box -2 -3 10 103
use BUFX4  BUFX4_124
timestamp 1693479267
transform -1 0 3116 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_113
timestamp 1693479267
transform 1 0 3116 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_360
timestamp 1693479267
transform 1 0 3148 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_203
timestamp 1693479267
transform 1 0 3172 0 1 1305
box -2 -3 26 103
use INVX1  INVX1_360
timestamp 1693479267
transform -1 0 3212 0 1 1305
box -2 -3 18 103
use NOR2X1  NOR2X1_160
timestamp 1693479267
transform 1 0 3212 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_201
timestamp 1693479267
transform 1 0 3236 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_431
timestamp 1693479267
transform -1 0 3284 0 1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_160
timestamp 1693479267
transform -1 0 3316 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_553
timestamp 1693479267
transform -1 0 3340 0 1 1305
box -2 -3 26 103
use AND2X2  AND2X2_50
timestamp 1693479267
transform -1 0 3372 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_557
timestamp 1693479267
transform -1 0 3396 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_662
timestamp 1693479267
transform 1 0 3396 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_265
timestamp 1693479267
transform -1 0 3452 0 1 1305
box -2 -3 26 103
use BUFX4  BUFX4_129
timestamp 1693479267
transform 1 0 3452 0 1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_45
timestamp 1693479267
transform -1 0 3532 0 1 1305
box -2 -3 50 103
use AOI21X1  AOI21X1_161
timestamp 1693479267
transform 1 0 3532 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_6_0
timestamp 1693479267
transform -1 0 3572 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_6_1
timestamp 1693479267
transform -1 0 3580 0 1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_651
timestamp 1693479267
transform -1 0 3612 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_432
timestamp 1693479267
transform -1 0 3636 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_323
timestamp 1693479267
transform -1 0 3660 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_566
timestamp 1693479267
transform 1 0 3660 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_322
timestamp 1693479267
transform 1 0 3684 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_730
timestamp 1693479267
transform -1 0 3740 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_558
timestamp 1693479267
transform 1 0 3740 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_419
timestamp 1693479267
transform 1 0 3764 0 1 1305
box -2 -3 26 103
use INVX1  INVX1_425
timestamp 1693479267
transform 1 0 3788 0 1 1305
box -2 -3 18 103
use AOI22X1  AOI22X1_106
timestamp 1693479267
transform -1 0 3844 0 1 1305
box -2 -3 42 103
use MUX2X1  MUX2X1_54
timestamp 1693479267
transform 1 0 3844 0 1 1305
box -2 -3 50 103
use BUFX4  BUFX4_84
timestamp 1693479267
transform 1 0 3892 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_330
timestamp 1693479267
transform -1 0 3948 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_359
timestamp 1693479267
transform -1 0 3972 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_575
timestamp 1693479267
transform 1 0 3972 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_576
timestamp 1693479267
transform 1 0 3996 0 1 1305
box -2 -3 26 103
use AND2X2  AND2X2_39
timestamp 1693479267
transform -1 0 4052 0 1 1305
box -2 -3 34 103
use AND2X2  AND2X2_40
timestamp 1693479267
transform 1 0 4052 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_7_0
timestamp 1693479267
transform 1 0 4084 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_7_1
timestamp 1693479267
transform 1 0 4092 0 1 1305
box -2 -3 10 103
use NOR2X1  NOR2X1_277
timestamp 1693479267
transform 1 0 4100 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_507
timestamp 1693479267
transform 1 0 4124 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_483
timestamp 1693479267
transform 1 0 4148 0 1 1305
box -2 -3 26 103
use MUX2X1  MUX2X1_53
timestamp 1693479267
transform 1 0 4172 0 1 1305
box -2 -3 50 103
use OAI21X1  OAI21X1_748
timestamp 1693479267
transform 1 0 4220 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_360
timestamp 1693479267
transform -1 0 4276 0 1 1305
box -2 -3 26 103
use AND2X2  AND2X2_74
timestamp 1693479267
transform 1 0 4276 0 1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_56
timestamp 1693479267
transform -1 0 4356 0 1 1305
box -2 -3 50 103
use BUFX4  BUFX4_55
timestamp 1693479267
transform 1 0 4356 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_672
timestamp 1693479267
transform 1 0 4388 0 1 1305
box -2 -3 34 103
use AND2X2  AND2X2_56
timestamp 1693479267
transform 1 0 4420 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_130
timestamp 1693479267
transform -1 0 4484 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_353
timestamp 1693479267
transform 1 0 4484 0 1 1305
box -2 -3 26 103
use MUX2X1  MUX2X1_52
timestamp 1693479267
transform 1 0 4508 0 1 1305
box -2 -3 50 103
use MUX2X1  MUX2X1_51
timestamp 1693479267
transform -1 0 4604 0 1 1305
box -2 -3 50 103
use BUFX2  BUFX2_31
timestamp 1693479267
transform -1 0 28 0 -1 1505
box -2 -3 26 103
use BUFX2  BUFX2_61
timestamp 1693479267
transform -1 0 52 0 -1 1505
box -2 -3 26 103
use CLKBUF1  CLKBUF1_6
timestamp 1693479267
transform -1 0 124 0 -1 1505
box -2 -3 74 103
use NOR3X1  NOR3X1_67
timestamp 1693479267
transform -1 0 188 0 -1 1505
box -2 -3 66 103
use INVX1  INVX1_487
timestamp 1693479267
transform -1 0 204 0 -1 1505
box -2 -3 18 103
use NOR2X1  NOR2X1_396
timestamp 1693479267
transform 1 0 204 0 -1 1505
box -2 -3 26 103
use INVX1  INVX1_486
timestamp 1693479267
transform 1 0 228 0 -1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_689
timestamp 1693479267
transform 1 0 244 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_695
timestamp 1693479267
transform -1 0 292 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_394
timestamp 1693479267
transform -1 0 316 0 -1 1505
box -2 -3 26 103
use BUFX4  BUFX4_241
timestamp 1693479267
transform 1 0 316 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_682
timestamp 1693479267
transform 1 0 348 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_395
timestamp 1693479267
transform -1 0 396 0 -1 1505
box -2 -3 26 103
use BUFX4  BUFX4_196
timestamp 1693479267
transform -1 0 428 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_684
timestamp 1693479267
transform 1 0 428 0 -1 1505
box -2 -3 26 103
use FILL  FILL_14_0_0
timestamp 1693479267
transform -1 0 460 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_0_1
timestamp 1693479267
transform -1 0 468 0 -1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_495
timestamp 1693479267
transform -1 0 564 0 -1 1505
box -2 -3 98 103
use NAND3X1  NAND3X1_53
timestamp 1693479267
transform -1 0 596 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_73
timestamp 1693479267
transform 1 0 596 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_462
timestamp 1693479267
transform 1 0 628 0 -1 1505
box -2 -3 98 103
use NAND3X1  NAND3X1_50
timestamp 1693479267
transform 1 0 724 0 -1 1505
box -2 -3 34 103
use XNOR2X1  XNOR2X1_42
timestamp 1693479267
transform 1 0 756 0 -1 1505
box -2 -3 58 103
use XOR2X1  XOR2X1_5
timestamp 1693479267
transform 1 0 812 0 -1 1505
box -2 -3 58 103
use OAI21X1  OAI21X1_266
timestamp 1693479267
transform 1 0 868 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_49
timestamp 1693479267
transform -1 0 924 0 -1 1505
box -2 -3 26 103
use INVX1  INVX1_277
timestamp 1693479267
transform 1 0 924 0 -1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_168
timestamp 1693479267
transform -1 0 964 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_269
timestamp 1693479267
transform -1 0 996 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_175
timestamp 1693479267
transform -1 0 1020 0 -1 1505
box -2 -3 26 103
use FILL  FILL_14_1_0
timestamp 1693479267
transform 1 0 1020 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_1_1
timestamp 1693479267
transform 1 0 1028 0 -1 1505
box -2 -3 10 103
use NAND3X1  NAND3X1_86
timestamp 1693479267
transform 1 0 1036 0 -1 1505
box -2 -3 34 103
use AND2X2  AND2X2_16
timestamp 1693479267
transform 1 0 1068 0 -1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_85
timestamp 1693479267
transform 1 0 1100 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_266
timestamp 1693479267
transform 1 0 1132 0 -1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_163
timestamp 1693479267
transform 1 0 1148 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_260
timestamp 1693479267
transform 1 0 1172 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_267
timestamp 1693479267
transform -1 0 1220 0 -1 1505
box -2 -3 18 103
use INVX1  INVX1_268
timestamp 1693479267
transform 1 0 1220 0 -1 1505
box -2 -3 18 103
use NAND3X1  NAND3X1_84
timestamp 1693479267
transform 1 0 1236 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_164
timestamp 1693479267
transform -1 0 1292 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_258
timestamp 1693479267
transform -1 0 1324 0 -1 1505
box -2 -3 34 103
use XNOR2X1  XNOR2X1_8
timestamp 1693479267
transform 1 0 1324 0 -1 1505
box -2 -3 58 103
use XNOR2X1  XNOR2X1_37
timestamp 1693479267
transform -1 0 1436 0 -1 1505
box -2 -3 58 103
use INVX1  INVX1_234
timestamp 1693479267
transform 1 0 1436 0 -1 1505
box -2 -3 18 103
use NAND3X1  NAND3X1_79
timestamp 1693479267
transform 1 0 1452 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_124
timestamp 1693479267
transform -1 0 1508 0 -1 1505
box -2 -3 26 103
use FILL  FILL_14_2_0
timestamp 1693479267
transform -1 0 1516 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_2_1
timestamp 1693479267
transform -1 0 1524 0 -1 1505
box -2 -3 10 103
use AOI22X1  AOI22X1_55
timestamp 1693479267
transform -1 0 1564 0 -1 1505
box -2 -3 42 103
use NAND2X1  NAND2X1_162
timestamp 1693479267
transform -1 0 1588 0 -1 1505
box -2 -3 26 103
use AOI22X1  AOI22X1_57
timestamp 1693479267
transform 1 0 1588 0 -1 1505
box -2 -3 42 103
use OAI21X1  OAI21X1_232
timestamp 1693479267
transform -1 0 1660 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_239
timestamp 1693479267
transform 1 0 1660 0 -1 1505
box -2 -3 18 103
use NOR3X1  NOR3X1_49
timestamp 1693479267
transform 1 0 1676 0 -1 1505
box -2 -3 66 103
use INVX1  INVX1_320
timestamp 1693479267
transform 1 0 1740 0 -1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_294
timestamp 1693479267
transform 1 0 1756 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_322
timestamp 1693479267
transform 1 0 1788 0 -1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_295
timestamp 1693479267
transform 1 0 1804 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_217
timestamp 1693479267
transform -1 0 1860 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_569
timestamp 1693479267
transform 1 0 1860 0 -1 1505
box -2 -3 26 103
use NAND3X1  NAND3X1_156
timestamp 1693479267
transform -1 0 1916 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_691
timestamp 1693479267
transform -1 0 1948 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_335
timestamp 1693479267
transform -1 0 1972 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_692
timestamp 1693479267
transform -1 0 2004 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_682
timestamp 1693479267
transform 1 0 2004 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_3_0
timestamp 1693479267
transform 1 0 2036 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_3_1
timestamp 1693479267
transform 1 0 2044 0 -1 1505
box -2 -3 10 103
use NOR2X1  NOR2X1_341
timestamp 1693479267
transform 1 0 2052 0 -1 1505
box -2 -3 26 103
use AND2X2  AND2X2_58
timestamp 1693479267
transform -1 0 2108 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_331
timestamp 1693479267
transform -1 0 2132 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_681
timestamp 1693479267
transform -1 0 2164 0 -1 1505
box -2 -3 34 103
use INVX2  INVX2_70
timestamp 1693479267
transform 1 0 2164 0 -1 1505
box -2 -3 18 103
use NAND3X1  NAND3X1_154
timestamp 1693479267
transform -1 0 2212 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_670
timestamp 1693479267
transform 1 0 2212 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_168
timestamp 1693479267
transform -1 0 2276 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_164
timestamp 1693479267
transform -1 0 2300 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_565
timestamp 1693479267
transform 1 0 2300 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_677
timestamp 1693479267
transform -1 0 2356 0 -1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_153
timestamp 1693479267
transform 1 0 2356 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_89
timestamp 1693479267
transform 1 0 2388 0 -1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_44
timestamp 1693479267
transform -1 0 2468 0 -1 1505
box -2 -3 50 103
use AND2X2  AND2X2_30
timestamp 1693479267
transform 1 0 2468 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_424
timestamp 1693479267
transform 1 0 2500 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_412
timestamp 1693479267
transform -1 0 2556 0 -1 1505
box -2 -3 26 103
use FILL  FILL_14_4_0
timestamp 1693479267
transform -1 0 2564 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_4_1
timestamp 1693479267
transform -1 0 2572 0 -1 1505
box -2 -3 10 103
use NAND2X1  NAND2X1_372
timestamp 1693479267
transform -1 0 2596 0 -1 1505
box -2 -3 26 103
use INVX8  INVX8_10
timestamp 1693479267
transform -1 0 2636 0 -1 1505
box -2 -3 42 103
use NAND3X1  NAND3X1_104
timestamp 1693479267
transform -1 0 2668 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_283
timestamp 1693479267
transform -1 0 2692 0 -1 1505
box -2 -3 26 103
use NAND3X1  NAND3X1_103
timestamp 1693479267
transform -1 0 2724 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_513
timestamp 1693479267
transform -1 0 2748 0 -1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_151
timestamp 1693479267
transform -1 0 2780 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_627
timestamp 1693479267
transform -1 0 2812 0 -1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_107
timestamp 1693479267
transform 1 0 2812 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_56
timestamp 1693479267
transform -1 0 2876 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_399
timestamp 1693479267
transform -1 0 2900 0 -1 1505
box -2 -3 26 103
use BUFX4  BUFX4_44
timestamp 1693479267
transform -1 0 2932 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_205
timestamp 1693479267
transform 1 0 2932 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_406
timestamp 1693479267
transform 1 0 2956 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_421
timestamp 1693479267
transform 1 0 2980 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_420
timestamp 1693479267
transform -1 0 3044 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_5_0
timestamp 1693479267
transform -1 0 3052 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_5_1
timestamp 1693479267
transform -1 0 3060 0 -1 1505
box -2 -3 10 103
use AOI21X1  AOI21X1_174
timestamp 1693479267
transform -1 0 3092 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_259
timestamp 1693479267
transform -1 0 3116 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_476
timestamp 1693479267
transform 1 0 3116 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_494
timestamp 1693479267
transform -1 0 3172 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_362
timestamp 1693479267
transform 1 0 3172 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_361
timestamp 1693479267
transform -1 0 3236 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_230
timestamp 1693479267
transform -1 0 3268 0 -1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_47
timestamp 1693479267
transform 1 0 3268 0 -1 1505
box -2 -3 50 103
use MUX2X1  MUX2X1_26
timestamp 1693479267
transform 1 0 3316 0 -1 1505
box -2 -3 50 103
use BUFX4  BUFX4_58
timestamp 1693479267
transform -1 0 3396 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_579
timestamp 1693479267
transform 1 0 3396 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_731
timestamp 1693479267
transform 1 0 3428 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_671
timestamp 1693479267
transform 1 0 3460 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_585
timestamp 1693479267
transform -1 0 3516 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_359
timestamp 1693479267
transform -1 0 3548 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_218
timestamp 1693479267
transform -1 0 3572 0 -1 1505
box -2 -3 26 103
use FILL  FILL_14_6_0
timestamp 1693479267
transform 1 0 3572 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_6_1
timestamp 1693479267
transform 1 0 3580 0 -1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_728
timestamp 1693479267
transform 1 0 3588 0 -1 1505
box -2 -3 34 103
use AND2X2  AND2X2_68
timestamp 1693479267
transform 1 0 3620 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_348
timestamp 1693479267
transform -1 0 3676 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_727
timestamp 1693479267
transform -1 0 3708 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_193
timestamp 1693479267
transform -1 0 3740 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_56
timestamp 1693479267
transform 1 0 3740 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_506
timestamp 1693479267
transform -1 0 3796 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_497
timestamp 1693479267
transform 1 0 3796 0 -1 1505
box -2 -3 34 103
use NOR3X1  NOR3X1_62
timestamp 1693479267
transform -1 0 3892 0 -1 1505
box -2 -3 66 103
use OAI21X1  OAI21X1_383
timestamp 1693479267
transform -1 0 3924 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_472
timestamp 1693479267
transform -1 0 3956 0 -1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_158
timestamp 1693479267
transform -1 0 3988 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_397
timestamp 1693479267
transform 1 0 3988 0 -1 1505
box -2 -3 18 103
use AOI21X1  AOI21X1_212
timestamp 1693479267
transform -1 0 4036 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_251
timestamp 1693479267
transform -1 0 4060 0 -1 1505
box -2 -3 26 103
use INVX8  INVX8_3
timestamp 1693479267
transform 1 0 4060 0 -1 1505
box -2 -3 42 103
use FILL  FILL_14_7_0
timestamp 1693479267
transform 1 0 4100 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_7_1
timestamp 1693479267
transform 1 0 4108 0 -1 1505
box -2 -3 10 103
use NAND2X1  NAND2X1_579
timestamp 1693479267
transform 1 0 4116 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_719
timestamp 1693479267
transform 1 0 4140 0 -1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_161
timestamp 1693479267
transform 1 0 4172 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_718
timestamp 1693479267
transform -1 0 4236 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_782
timestamp 1693479267
transform -1 0 4268 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_213
timestamp 1693479267
transform -1 0 4300 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_345
timestamp 1693479267
transform -1 0 4324 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_780
timestamp 1693479267
transform 1 0 4324 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_604
timestamp 1693479267
transform -1 0 4380 0 -1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_210
timestamp 1693479267
transform 1 0 4380 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_768
timestamp 1693479267
transform 1 0 4412 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_371
timestamp 1693479267
transform 1 0 4444 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_767
timestamp 1693479267
transform -1 0 4500 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_591
timestamp 1693479267
transform 1 0 4500 0 -1 1505
box -2 -3 26 103
use OAI22X1  OAI22X1_40
timestamp 1693479267
transform -1 0 4564 0 -1 1505
box -2 -3 42 103
use NAND2X1  NAND2X1_259
timestamp 1693479267
transform -1 0 4588 0 -1 1505
box -2 -3 26 103
use FILL  FILL_15_1
timestamp 1693479267
transform -1 0 4596 0 -1 1505
box -2 -3 10 103
use FILL  FILL_15_2
timestamp 1693479267
transform -1 0 4604 0 -1 1505
box -2 -3 10 103
use BUFX2  BUFX2_70
timestamp 1693479267
transform -1 0 28 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_188
timestamp 1693479267
transform -1 0 124 0 1 1505
box -2 -3 98 103
use BUFX2  BUFX2_32
timestamp 1693479267
transform -1 0 28 0 -1 1705
box -2 -3 26 103
use BUFX2  BUFX2_69
timestamp 1693479267
transform -1 0 52 0 -1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_189
timestamp 1693479267
transform -1 0 148 0 -1 1705
box -2 -3 98 103
use BUFX2  BUFX2_62
timestamp 1693479267
transform -1 0 148 0 1 1505
box -2 -3 26 103
use NOR3X1  NOR3X1_66
timestamp 1693479267
transform -1 0 212 0 1 1505
box -2 -3 66 103
use NAND2X1  NAND2X1_694
timestamp 1693479267
transform 1 0 148 0 -1 1705
box -2 -3 26 103
use INVX1  INVX1_492
timestamp 1693479267
transform 1 0 172 0 -1 1705
box -2 -3 18 103
use AOI21X1  AOI21X1_221
timestamp 1693479267
transform 1 0 188 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_686
timestamp 1693479267
transform 1 0 212 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_860
timestamp 1693479267
transform -1 0 268 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_866
timestamp 1693479267
transform 1 0 268 0 1 1505
box -2 -3 34 103
use NOR3X1  NOR3X1_68
timestamp 1693479267
transform -1 0 364 0 1 1505
box -2 -3 66 103
use INVX1  INVX1_491
timestamp 1693479267
transform 1 0 220 0 -1 1705
box -2 -3 18 103
use NAND3X1  NAND3X1_185
timestamp 1693479267
transform 1 0 236 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_490
timestamp 1693479267
transform 1 0 268 0 -1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_397
timestamp 1693479267
transform -1 0 308 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_867
timestamp 1693479267
transform 1 0 364 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_398
timestamp 1693479267
transform -1 0 420 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_863
timestamp 1693479267
transform -1 0 340 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_864
timestamp 1693479267
transform 1 0 340 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_494
timestamp 1693479267
transform -1 0 388 0 -1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_693
timestamp 1693479267
transform -1 0 412 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_868
timestamp 1693479267
transform 1 0 420 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_857
timestamp 1693479267
transform -1 0 484 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_683
timestamp 1693479267
transform -1 0 508 0 1 1505
box -2 -3 26 103
use FILL  FILL_15_0_0
timestamp 1693479267
transform -1 0 516 0 1 1505
box -2 -3 10 103
use NAND2X1  NAND2X1_696
timestamp 1693479267
transform 1 0 412 0 -1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_502
timestamp 1693479267
transform -1 0 532 0 -1 1705
box -2 -3 98 103
use FILL  FILL_15_0_1
timestamp 1693479267
transform -1 0 524 0 1 1505
box -2 -3 10 103
use INVX1  INVX1_493
timestamp 1693479267
transform -1 0 540 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_191
timestamp 1693479267
transform -1 0 572 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_192
timestamp 1693479267
transform -1 0 604 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_185
timestamp 1693479267
transform 1 0 604 0 1 1505
box -2 -3 34 103
use FILL  FILL_16_0_0
timestamp 1693479267
transform -1 0 540 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_0_1
timestamp 1693479267
transform -1 0 548 0 -1 1705
box -2 -3 10 103
use NAND3X1  NAND3X1_67
timestamp 1693479267
transform -1 0 580 0 -1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_470
timestamp 1693479267
transform 1 0 580 0 -1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_463
timestamp 1693479267
transform 1 0 636 0 1 1505
box -2 -3 98 103
use NAND3X1  NAND3X1_66
timestamp 1693479267
transform 1 0 676 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_52
timestamp 1693479267
transform 1 0 708 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_55
timestamp 1693479267
transform -1 0 764 0 1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_69
timestamp 1693479267
transform 1 0 764 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_503
timestamp 1693479267
transform 1 0 796 0 1 1505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_496
timestamp 1693479267
transform 1 0 740 0 -1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_471
timestamp 1693479267
transform 1 0 892 0 1 1505
box -2 -3 98 103
use NAND3X1  NAND3X1_54
timestamp 1693479267
transform -1 0 868 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_68
timestamp 1693479267
transform -1 0 900 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_5
timestamp 1693479267
transform -1 0 932 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_167
timestamp 1693479267
transform -1 0 1012 0 1 1505
box -2 -3 26 103
use FILL  FILL_15_1_0
timestamp 1693479267
transform -1 0 1020 0 1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_464
timestamp 1693479267
transform 1 0 932 0 -1 1705
box -2 -3 98 103
use FILL  FILL_15_1_1
timestamp 1693479267
transform -1 0 1028 0 1 1505
box -2 -3 10 103
use OR2X2  OR2X2_12
timestamp 1693479267
transform -1 0 1060 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_173
timestamp 1693479267
transform 1 0 1060 0 1 1505
box -2 -3 26 103
use INVX1  INVX1_276
timestamp 1693479267
transform 1 0 1084 0 1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_174
timestamp 1693479267
transform 1 0 1100 0 1 1505
box -2 -3 26 103
use FILL  FILL_16_1_0
timestamp 1693479267
transform 1 0 1028 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_1_1
timestamp 1693479267
transform 1 0 1036 0 -1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_276
timestamp 1693479267
transform 1 0 1044 0 -1 1705
box -2 -3 98 103
use INVX1  INVX1_275
timestamp 1693479267
transform -1 0 1140 0 1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_170
timestamp 1693479267
transform -1 0 1164 0 1 1505
box -2 -3 26 103
use OR2X2  OR2X2_13
timestamp 1693479267
transform -1 0 1196 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_169
timestamp 1693479267
transform -1 0 1220 0 1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_34
timestamp 1693479267
transform 1 0 1140 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_299
timestamp 1693479267
transform 1 0 1172 0 -1 1705
box -2 -3 18 103
use AOI21X1  AOI21X1_36
timestamp 1693479267
transform -1 0 1220 0 -1 1705
box -2 -3 34 103
use XNOR2X1  XNOR2X1_10
timestamp 1693479267
transform 1 0 1220 0 1 1505
box -2 -3 58 103
use NOR3X1  NOR3X1_55
timestamp 1693479267
transform -1 0 1340 0 1 1505
box -2 -3 66 103
use INVX1  INVX1_287
timestamp 1693479267
transform 1 0 1220 0 -1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_273
timestamp 1693479267
transform -1 0 1268 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_51
timestamp 1693479267
transform 1 0 1268 0 -1 1705
box -2 -3 26 103
use INVX1  INVX1_273
timestamp 1693479267
transform -1 0 1308 0 -1 1705
box -2 -3 18 103
use INVX1  INVX1_264
timestamp 1693479267
transform -1 0 1324 0 -1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_228
timestamp 1693479267
transform 1 0 1340 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_27
timestamp 1693479267
transform 1 0 1372 0 1 1505
box -2 -3 26 103
use INVX1  INVX1_233
timestamp 1693479267
transform 1 0 1396 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_257
timestamp 1693479267
transform 1 0 1412 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_172
timestamp 1693479267
transform -1 0 1348 0 -1 1705
box -2 -3 26 103
use INVX2  INVX2_6
timestamp 1693479267
transform 1 0 1348 0 -1 1705
box -2 -3 18 103
use XNOR2X1  XNOR2X1_7
timestamp 1693479267
transform 1 0 1364 0 -1 1705
box -2 -3 58 103
use INVX1  INVX1_262
timestamp 1693479267
transform -1 0 1460 0 1 1505
box -2 -3 18 103
use AOI21X1  AOI21X1_7
timestamp 1693479267
transform -1 0 1492 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_123
timestamp 1693479267
transform -1 0 1516 0 1 1505
box -2 -3 26 103
use FILL  FILL_15_2_0
timestamp 1693479267
transform 1 0 1516 0 1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_277
timestamp 1693479267
transform 1 0 1420 0 -1 1705
box -2 -3 98 103
use FILL  FILL_16_2_0
timestamp 1693479267
transform 1 0 1516 0 -1 1705
box -2 -3 10 103
use FILL  FILL_15_2_1
timestamp 1693479267
transform 1 0 1524 0 1 1505
box -2 -3 10 103
use NOR2X1  NOR2X1_28
timestamp 1693479267
transform 1 0 1532 0 1 1505
box -2 -3 26 103
use XNOR2X1  XNOR2X1_9
timestamp 1693479267
transform -1 0 1612 0 1 1505
box -2 -3 58 103
use BUFX4  BUFX4_146
timestamp 1693479267
transform 1 0 1612 0 1 1505
box -2 -3 34 103
use FILL  FILL_16_2_1
timestamp 1693479267
transform 1 0 1524 0 -1 1705
box -2 -3 10 103
use INVX2  INVX2_7
timestamp 1693479267
transform 1 0 1532 0 -1 1705
box -2 -3 18 103
use XNOR2X1  XNOR2X1_6
timestamp 1693479267
transform 1 0 1548 0 -1 1705
box -2 -3 58 103
use NAND3X1  NAND3X1_78
timestamp 1693479267
transform 1 0 1604 0 -1 1705
box -2 -3 34 103
use AOI22X1  AOI22X1_58
timestamp 1693479267
transform 1 0 1644 0 1 1505
box -2 -3 42 103
use BUFX4  BUFX4_234
timestamp 1693479267
transform -1 0 1716 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_235
timestamp 1693479267
transform 1 0 1716 0 1 1505
box -2 -3 18 103
use XNOR2X1  XNOR2X1_11
timestamp 1693479267
transform 1 0 1636 0 -1 1705
box -2 -3 58 103
use AOI22X1  AOI22X1_60
timestamp 1693479267
transform -1 0 1732 0 -1 1705
box -2 -3 42 103
use AOI21X1  AOI21X1_8
timestamp 1693479267
transform -1 0 1764 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_213
timestamp 1693479267
transform -1 0 1788 0 1 1505
box -2 -3 26 103
use INVX4  INVX4_4
timestamp 1693479267
transform 1 0 1788 0 1 1505
box -2 -3 26 103
use NAND3X1  NAND3X1_155
timestamp 1693479267
transform -1 0 1844 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_227
timestamp 1693479267
transform -1 0 1764 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_77
timestamp 1693479267
transform -1 0 1796 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_4
timestamp 1693479267
transform -1 0 1828 0 -1 1705
box -2 -3 34 103
use OR2X2  OR2X2_38
timestamp 1693479267
transform -1 0 1876 0 1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_157
timestamp 1693479267
transform 1 0 1876 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_179
timestamp 1693479267
transform -1 0 1940 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_117
timestamp 1693479267
transform -1 0 1852 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_231
timestamp 1693479267
transform 1 0 1852 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_118
timestamp 1693479267
transform -1 0 1908 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_210
timestamp 1693479267
transform -1 0 1932 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_684
timestamp 1693479267
transform -1 0 1972 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_38
timestamp 1693479267
transform -1 0 2004 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_100
timestamp 1693479267
transform -1 0 2028 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_293
timestamp 1693479267
transform -1 0 1964 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_319
timestamp 1693479267
transform -1 0 1980 0 -1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_208
timestamp 1693479267
transform 1 0 1980 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_291
timestamp 1693479267
transform 1 0 2004 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_206
timestamp 1693479267
transform 1 0 2052 0 -1 1705
box -2 -3 26 103
use FILL  FILL_16_3_1
timestamp 1693479267
transform 1 0 2044 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_3_0
timestamp 1693479267
transform 1 0 2036 0 -1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_683
timestamp 1693479267
transform -1 0 2076 0 1 1505
box -2 -3 34 103
use FILL  FILL_15_3_1
timestamp 1693479267
transform -1 0 2044 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_3_0
timestamp 1693479267
transform -1 0 2036 0 1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_292
timestamp 1693479267
transform -1 0 2108 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_333
timestamp 1693479267
transform -1 0 2100 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_99
timestamp 1693479267
transform -1 0 2148 0 -1 1705
box -2 -3 26 103
use INVX1  INVX1_318
timestamp 1693479267
transform -1 0 2124 0 -1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_211
timestamp 1693479267
transform 1 0 2116 0 1 1505
box -2 -3 26 103
use INVX2  INVX2_29
timestamp 1693479267
transform 1 0 2100 0 1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_562
timestamp 1693479267
transform -1 0 2164 0 1 1505
box -2 -3 26 103
use AOI22X1  AOI22X1_69
timestamp 1693479267
transform -1 0 2204 0 1 1505
box -2 -3 42 103
use NAND2X1  NAND2X1_234
timestamp 1693479267
transform -1 0 2228 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_332
timestamp 1693479267
transform -1 0 2172 0 -1 1705
box -2 -3 26 103
use INVX1  INVX1_317
timestamp 1693479267
transform -1 0 2188 0 -1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_207
timestamp 1693479267
transform 1 0 2188 0 -1 1705
box -2 -3 26 103
use AND2X2  AND2X2_59
timestamp 1693479267
transform 1 0 2212 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_175
timestamp 1693479267
transform 1 0 2228 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_414
timestamp 1693479267
transform 1 0 2260 0 1 1505
box -2 -3 18 103
use INVX1  INVX1_412
timestamp 1693479267
transform 1 0 2276 0 1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_212
timestamp 1693479267
transform -1 0 2316 0 1 1505
box -2 -3 26 103
use AOI22X1  AOI22X1_103
timestamp 1693479267
transform 1 0 2316 0 1 1505
box -2 -3 42 103
use NAND2X1  NAND2X1_209
timestamp 1693479267
transform -1 0 2268 0 -1 1705
box -2 -3 26 103
use MUX2X1  MUX2X1_14
timestamp 1693479267
transform -1 0 2316 0 -1 1705
box -2 -3 50 103
use INVX8  INVX8_11
timestamp 1693479267
transform -1 0 2356 0 -1 1705
box -2 -3 42 103
use OAI21X1  OAI21X1_676
timestamp 1693479267
transform 1 0 2356 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_689
timestamp 1693479267
transform 1 0 2388 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_568
timestamp 1693479267
transform 1 0 2420 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_272
timestamp 1693479267
transform -1 0 2380 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_317
timestamp 1693479267
transform -1 0 2412 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_340
timestamp 1693479267
transform -1 0 2428 0 -1 1705
box -2 -3 18 103
use BUFX4  BUFX4_187
timestamp 1693479267
transform -1 0 2476 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_373
timestamp 1693479267
transform -1 0 2508 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_413
timestamp 1693479267
transform -1 0 2532 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_181
timestamp 1693479267
transform -1 0 2452 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_352
timestamp 1693479267
transform -1 0 2476 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_179
timestamp 1693479267
transform -1 0 2500 0 -1 1705
box -2 -3 26 103
use OR2X2  OR2X2_22
timestamp 1693479267
transform 1 0 2500 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_4_1
timestamp 1693479267
transform 1 0 2564 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_4_0
timestamp 1693479267
transform 1 0 2556 0 -1 1705
box -2 -3 10 103
use NAND2X1  NAND2X1_353
timestamp 1693479267
transform 1 0 2532 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_388
timestamp 1693479267
transform 1 0 2564 0 1 1505
box -2 -3 34 103
use FILL  FILL_15_4_1
timestamp 1693479267
transform 1 0 2556 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_4_0
timestamp 1693479267
transform 1 0 2548 0 1 1505
box -2 -3 10 103
use INVX2  INVX2_30
timestamp 1693479267
transform -1 0 2548 0 1 1505
box -2 -3 18 103
use NOR2X1  NOR2X1_176
timestamp 1693479267
transform -1 0 2620 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_180
timestamp 1693479267
transform 1 0 2572 0 -1 1705
box -2 -3 26 103
use BUFX4  BUFX4_90
timestamp 1693479267
transform -1 0 2628 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_178
timestamp 1693479267
transform 1 0 2620 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_374
timestamp 1693479267
transform 1 0 2628 0 1 1505
box -2 -3 34 103
use AND2X2  AND2X2_27
timestamp 1693479267
transform 1 0 2660 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_277
timestamp 1693479267
transform -1 0 2724 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_394
timestamp 1693479267
transform 1 0 2724 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_375
timestamp 1693479267
transform 1 0 2644 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_258
timestamp 1693479267
transform 1 0 2676 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_345
timestamp 1693479267
transform -1 0 2724 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_346
timestamp 1693479267
transform -1 0 2748 0 -1 1705
box -2 -3 26 103
use NOR3X1  NOR3X1_56
timestamp 1693479267
transform 1 0 2740 0 1 1505
box -2 -3 66 103
use OAI21X1  OAI21X1_341
timestamp 1693479267
transform 1 0 2804 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_186
timestamp 1693479267
transform -1 0 2772 0 -1 1705
box -2 -3 26 103
use OR2X2  OR2X2_23
timestamp 1693479267
transform -1 0 2804 0 -1 1705
box -2 -3 34 103
use AND2X2  AND2X2_42
timestamp 1693479267
transform 1 0 2804 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_110
timestamp 1693479267
transform -1 0 2868 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_207
timestamp 1693479267
transform 1 0 2868 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_208
timestamp 1693479267
transform -1 0 2916 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_407
timestamp 1693479267
transform -1 0 2940 0 1 1505
box -2 -3 26 103
use BUFX4  BUFX4_152
timestamp 1693479267
transform 1 0 2836 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_377
timestamp 1693479267
transform -1 0 2900 0 -1 1705
box -2 -3 34 103
use OR2X2  OR2X2_24
timestamp 1693479267
transform -1 0 2932 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_316
timestamp 1693479267
transform 1 0 2932 0 -1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_422
timestamp 1693479267
transform -1 0 2972 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_206
timestamp 1693479267
transform -1 0 2996 0 1 1505
box -2 -3 26 103
use AND2X2  AND2X2_29
timestamp 1693479267
transform 1 0 2996 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_538
timestamp 1693479267
transform -1 0 3060 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_46
timestamp 1693479267
transform 1 0 2948 0 -1 1705
box -2 -3 34 103
use AOI22X1  AOI22X1_95
timestamp 1693479267
transform 1 0 2980 0 -1 1705
box -2 -3 42 103
use NOR2X1  NOR2X1_267
timestamp 1693479267
transform -1 0 3044 0 -1 1705
box -2 -3 26 103
use FILL  FILL_15_5_0
timestamp 1693479267
transform -1 0 3068 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_5_1
timestamp 1693479267
transform -1 0 3076 0 1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_536
timestamp 1693479267
transform -1 0 3108 0 1 1505
box -2 -3 34 103
use AND2X2  AND2X2_44
timestamp 1693479267
transform -1 0 3140 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_266
timestamp 1693479267
transform -1 0 3068 0 -1 1705
box -2 -3 26 103
use FILL  FILL_16_5_0
timestamp 1693479267
transform 1 0 3068 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_5_1
timestamp 1693479267
transform 1 0 3076 0 -1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_537
timestamp 1693479267
transform 1 0 3084 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_495
timestamp 1693479267
transform 1 0 3116 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_260
timestamp 1693479267
transform 1 0 3140 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_412
timestamp 1693479267
transform 1 0 3164 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_398
timestamp 1693479267
transform -1 0 3220 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_413
timestamp 1693479267
transform -1 0 3252 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_199
timestamp 1693479267
transform 1 0 3140 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_396
timestamp 1693479267
transform 1 0 3164 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_535
timestamp 1693479267
transform 1 0 3188 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_127
timestamp 1693479267
transform 1 0 3220 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_169
timestamp 1693479267
transform -1 0 3284 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_492
timestamp 1693479267
transform -1 0 3308 0 1 1505
box -2 -3 26 103
use INVX4  INVX4_7
timestamp 1693479267
transform 1 0 3308 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_256
timestamp 1693479267
transform 1 0 3332 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_263
timestamp 1693479267
transform -1 0 3276 0 -1 1705
box -2 -3 26 103
use MUX2X1  MUX2X1_46
timestamp 1693479267
transform -1 0 3324 0 -1 1705
box -2 -3 50 103
use NAND2X1  NAND2X1_371
timestamp 1693479267
transform -1 0 3348 0 -1 1705
box -2 -3 26 103
use MUX2X1  MUX2X1_29
timestamp 1693479267
transform -1 0 3404 0 1 1505
box -2 -3 50 103
use NAND2X1  NAND2X1_373
timestamp 1693479267
transform -1 0 3428 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_700
timestamp 1693479267
transform -1 0 3460 0 1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_28
timestamp 1693479267
transform 1 0 3348 0 -1 1705
box -2 -3 50 103
use OR2X2  OR2X2_40
timestamp 1693479267
transform 1 0 3396 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_389
timestamp 1693479267
transform -1 0 3460 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_225
timestamp 1693479267
transform -1 0 3492 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_336
timestamp 1693479267
transform -1 0 3516 0 1 1505
box -2 -3 26 103
use INVX8  INVX8_5
timestamp 1693479267
transform -1 0 3556 0 1 1505
box -2 -3 42 103
use NOR2X1  NOR2X1_261
timestamp 1693479267
transform 1 0 3460 0 -1 1705
box -2 -3 26 103
use MUX2X1  MUX2X1_20
timestamp 1693479267
transform -1 0 3532 0 -1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_19
timestamp 1693479267
transform 1 0 3532 0 -1 1705
box -2 -3 50 103
use NAND2X1  NAND2X1_595
timestamp 1693479267
transform 1 0 3556 0 1 1505
box -2 -3 26 103
use FILL  FILL_15_6_0
timestamp 1693479267
transform -1 0 3588 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_6_1
timestamp 1693479267
transform -1 0 3596 0 1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_747
timestamp 1693479267
transform -1 0 3628 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_726
timestamp 1693479267
transform -1 0 3660 0 1 1505
box -2 -3 34 103
use FILL  FILL_16_6_0
timestamp 1693479267
transform 1 0 3580 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_6_1
timestamp 1693479267
transform 1 0 3588 0 -1 1705
box -2 -3 10 103
use BUFX4  BUFX4_224
timestamp 1693479267
transform 1 0 3596 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_586
timestamp 1693479267
transform -1 0 3652 0 -1 1705
box -2 -3 26 103
use NOR3X1  NOR3X1_63
timestamp 1693479267
transform 1 0 3660 0 1 1505
box -2 -3 66 103
use AND2X2  AND2X2_66
timestamp 1693479267
transform 1 0 3724 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_580
timestamp 1693479267
transform -1 0 3676 0 -1 1705
box -2 -3 26 103
use NAND3X1  NAND3X1_164
timestamp 1693479267
transform 1 0 3676 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_364
timestamp 1693479267
transform 1 0 3708 0 -1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_715
timestamp 1693479267
transform -1 0 3756 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_211
timestamp 1693479267
transform -1 0 3788 0 1 1505
box -2 -3 34 103
use INVX2  INVX2_62
timestamp 1693479267
transform 1 0 3788 0 1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_466
timestamp 1693479267
transform 1 0 3804 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_236
timestamp 1693479267
transform 1 0 3828 0 1 1505
box -2 -3 26 103
use INVX1  INVX1_420
timestamp 1693479267
transform -1 0 3772 0 -1 1705
box -2 -3 18 103
use MUX2X1  MUX2X1_32
timestamp 1693479267
transform 1 0 3772 0 -1 1705
box -2 -3 50 103
use OAI21X1  OAI21X1_737
timestamp 1693479267
transform -1 0 3852 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_528
timestamp 1693479267
transform -1 0 3876 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_367
timestamp 1693479267
transform 1 0 3876 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_223
timestamp 1693479267
transform -1 0 3924 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_439
timestamp 1693479267
transform -1 0 3948 0 1 1505
box -2 -3 26 103
use INVX1  INVX1_381
timestamp 1693479267
transform 1 0 3852 0 -1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_441
timestamp 1693479267
transform 1 0 3868 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_442
timestamp 1693479267
transform 1 0 3900 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_775
timestamp 1693479267
transform -1 0 3964 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_212
timestamp 1693479267
transform 1 0 3948 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_289
timestamp 1693479267
transform -1 0 4004 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_738
timestamp 1693479267
transform 1 0 4004 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_209
timestamp 1693479267
transform 1 0 4036 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_776
timestamp 1693479267
transform 1 0 3964 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_777
timestamp 1693479267
transform -1 0 4028 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_590
timestamp 1693479267
transform -1 0 4052 0 -1 1705
box -2 -3 26 103
use FILL  FILL_15_7_0
timestamp 1693479267
transform 1 0 4068 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_7_1
timestamp 1693479267
transform 1 0 4076 0 1 1505
box -2 -3 10 103
use MUX2X1  MUX2X1_49
timestamp 1693479267
transform 1 0 4084 0 1 1505
box -2 -3 50 103
use AOI21X1  AOI21X1_188
timestamp 1693479267
transform -1 0 4164 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_757
timestamp 1693479267
transform 1 0 4052 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_7_0
timestamp 1693479267
transform 1 0 4084 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_7_1
timestamp 1693479267
transform 1 0 4092 0 -1 1705
box -2 -3 10 103
use OAI22X1  OAI22X1_42
timestamp 1693479267
transform 1 0 4100 0 -1 1705
box -2 -3 42 103
use NAND2X1  NAND2X1_581
timestamp 1693479267
transform 1 0 4140 0 -1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_189
timestamp 1693479267
transform -1 0 4196 0 1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_163
timestamp 1693479267
transform -1 0 4228 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_716
timestamp 1693479267
transform 1 0 4228 0 1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_162
timestamp 1693479267
transform 1 0 4164 0 -1 1705
box -2 -3 34 103
use OR2X2  OR2X2_20
timestamp 1693479267
transform 1 0 4196 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_165
timestamp 1693479267
transform -1 0 4252 0 -1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_201
timestamp 1693479267
transform 1 0 4260 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_717
timestamp 1693479267
transform -1 0 4324 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_344
timestamp 1693479267
transform -1 0 4348 0 1 1505
box -2 -3 26 103
use OR2X2  OR2X2_42
timestamp 1693479267
transform 1 0 4252 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_168
timestamp 1693479267
transform 1 0 4284 0 -1 1705
box -2 -3 34 103
use OR2X2  OR2X2_41
timestamp 1693479267
transform 1 0 4316 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_511
timestamp 1693479267
transform -1 0 4372 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_512
timestamp 1693479267
transform -1 0 4396 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_772
timestamp 1693479267
transform -1 0 4428 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_770
timestamp 1693479267
transform -1 0 4460 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_197
timestamp 1693479267
transform -1 0 4380 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_760
timestamp 1693479267
transform 1 0 4380 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_369
timestamp 1693479267
transform -1 0 4436 0 -1 1705
box -2 -3 26 103
use NOR3X1  NOR3X1_64
timestamp 1693479267
transform 1 0 4436 0 -1 1705
box -2 -3 66 103
use OAI21X1  OAI21X1_769
timestamp 1693479267
transform 1 0 4460 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_601
timestamp 1693479267
transform 1 0 4492 0 1 1505
box -2 -3 26 103
use AND2X2  AND2X2_71
timestamp 1693479267
transform 1 0 4516 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_198
timestamp 1693479267
transform 1 0 4548 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_739
timestamp 1693479267
transform 1 0 4500 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_347
timestamp 1693479267
transform -1 0 4556 0 -1 1705
box -2 -3 26 103
use FILL  FILL_16_1
timestamp 1693479267
transform 1 0 4580 0 1 1505
box -2 -3 10 103
use FILL  FILL_16_2
timestamp 1693479267
transform 1 0 4588 0 1 1505
box -2 -3 10 103
use FILL  FILL_16_3
timestamp 1693479267
transform 1 0 4596 0 1 1505
box -2 -3 10 103
use NOR2X1  NOR2X1_346
timestamp 1693479267
transform -1 0 4580 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_352
timestamp 1693479267
transform -1 0 4604 0 -1 1705
box -2 -3 26 103
use BUFX2  BUFX2_63
timestamp 1693479267
transform -1 0 28 0 1 1705
box -2 -3 26 103
use BUFX2  BUFX2_66
timestamp 1693479267
transform -1 0 52 0 1 1705
box -2 -3 26 103
use BUFX2  BUFX2_65
timestamp 1693479267
transform -1 0 76 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_467
timestamp 1693479267
transform 1 0 76 0 1 1705
box -2 -3 98 103
use XNOR2X1  XNOR2X1_53
timestamp 1693479267
transform 1 0 172 0 1 1705
box -2 -3 58 103
use NAND2X1  NAND2X1_690
timestamp 1693479267
transform 1 0 228 0 1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_220
timestamp 1693479267
transform 1 0 252 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_861
timestamp 1693479267
transform 1 0 284 0 1 1705
box -2 -3 34 103
use XNOR2X1  XNOR2X1_52
timestamp 1693479267
transform 1 0 316 0 1 1705
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_499
timestamp 1693479267
transform -1 0 468 0 1 1705
box -2 -3 98 103
use FILL  FILL_17_0_0
timestamp 1693479267
transform -1 0 476 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_0_1
timestamp 1693479267
transform -1 0 484 0 1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_498
timestamp 1693479267
transform -1 0 580 0 1 1705
box -2 -3 98 103
use NAND3X1  NAND3X1_59
timestamp 1693479267
transform 1 0 580 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_466
timestamp 1693479267
transform 1 0 612 0 1 1705
box -2 -3 98 103
use NAND3X1  NAND3X1_58
timestamp 1693479267
transform 1 0 708 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_136
timestamp 1693479267
transform 1 0 740 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_76
timestamp 1693479267
transform -1 0 804 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_114
timestamp 1693479267
transform 1 0 804 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_64
timestamp 1693479267
transform -1 0 868 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_280
timestamp 1693479267
transform 1 0 868 0 1 1705
box -2 -3 98 103
use NOR2X1  NOR2X1_67
timestamp 1693479267
transform 1 0 964 0 1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_66
timestamp 1693479267
transform -1 0 1012 0 1 1705
box -2 -3 26 103
use FILL  FILL_17_1_0
timestamp 1693479267
transform -1 0 1020 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_1_1
timestamp 1693479267
transform -1 0 1028 0 1 1705
box -2 -3 10 103
use NAND2X1  NAND2X1_191
timestamp 1693479267
transform -1 0 1052 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_298
timestamp 1693479267
transform 1 0 1052 0 1 1705
box -2 -3 18 103
use AOI21X1  AOI21X1_35
timestamp 1693479267
transform -1 0 1100 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_295
timestamp 1693479267
transform -1 0 1116 0 1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_277
timestamp 1693479267
transform -1 0 1148 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_293
timestamp 1693479267
transform -1 0 1164 0 1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_279
timestamp 1693479267
transform -1 0 1196 0 1 1705
box -2 -3 34 103
use XOR2X1  XOR2X1_6
timestamp 1693479267
transform 1 0 1196 0 1 1705
box -2 -3 58 103
use OAI21X1  OAI21X1_280
timestamp 1693479267
transform 1 0 1252 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_192
timestamp 1693479267
transform -1 0 1308 0 1 1705
box -2 -3 26 103
use OR2X2  OR2X2_14
timestamp 1693479267
transform -1 0 1340 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_171
timestamp 1693479267
transform 1 0 1340 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_278
timestamp 1693479267
transform 1 0 1364 0 1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_285
timestamp 1693479267
transform 1 0 1460 0 1 1705
box -2 -3 98 103
use FILL  FILL_17_2_0
timestamp 1693479267
transform -1 0 1564 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_2_1
timestamp 1693479267
transform -1 0 1572 0 1 1705
box -2 -3 10 103
use INVX1  INVX1_231
timestamp 1693479267
transform -1 0 1588 0 1 1705
box -2 -3 18 103
use NAND3X1  NAND3X1_75
timestamp 1693479267
transform -1 0 1620 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_149
timestamp 1693479267
transform 1 0 1620 0 1 1705
box -2 -3 34 103
use AOI22X1  AOI22X1_59
timestamp 1693479267
transform 1 0 1652 0 1 1705
box -2 -3 42 103
use BUFX4  BUFX4_233
timestamp 1693479267
transform -1 0 1724 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_232
timestamp 1693479267
transform 1 0 1724 0 1 1705
box -2 -3 18 103
use NAND3X1  NAND3X1_76
timestamp 1693479267
transform 1 0 1740 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_25
timestamp 1693479267
transform 1 0 1772 0 1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_24
timestamp 1693479267
transform -1 0 1820 0 1 1705
box -2 -3 26 103
use AND2X2  AND2X2_10
timestamp 1693479267
transform 1 0 1820 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_346
timestamp 1693479267
transform 1 0 1852 0 1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_177
timestamp 1693479267
transform -1 0 1892 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_310
timestamp 1693479267
transform 1 0 1892 0 1 1705
box -2 -3 26 103
use NAND3X1  NAND3X1_101
timestamp 1693479267
transform 1 0 1916 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_129
timestamp 1693479267
transform 1 0 1948 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_311
timestamp 1693479267
transform 1 0 1972 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_301
timestamp 1693479267
transform -1 0 2012 0 1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_70
timestamp 1693479267
transform -1 0 2036 0 1 1705
box -2 -3 26 103
use FILL  FILL_17_3_0
timestamp 1693479267
transform -1 0 2044 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_3_1
timestamp 1693479267
transform -1 0 2052 0 1 1705
box -2 -3 10 103
use NAND2X1  NAND2X1_195
timestamp 1693479267
transform -1 0 2076 0 1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_131
timestamp 1693479267
transform 1 0 2076 0 1 1705
box -2 -3 26 103
use OR2X2  OR2X2_16
timestamp 1693479267
transform -1 0 2132 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_128
timestamp 1693479267
transform -1 0 2156 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_312
timestamp 1693479267
transform 1 0 2156 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_313
timestamp 1693479267
transform 1 0 2180 0 1 1705
box -2 -3 26 103
use AND2X2  AND2X2_24
timestamp 1693479267
transform 1 0 2204 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_130
timestamp 1693479267
transform -1 0 2260 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_358
timestamp 1693479267
transform 1 0 2260 0 1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_154
timestamp 1693479267
transform -1 0 2300 0 1 1705
box -2 -3 26 103
use INVX2  INVX2_51
timestamp 1693479267
transform -1 0 2316 0 1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_155
timestamp 1693479267
transform -1 0 2340 0 1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_132
timestamp 1693479267
transform -1 0 2364 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_347
timestamp 1693479267
transform 1 0 2364 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_349
timestamp 1693479267
transform -1 0 2412 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_372
timestamp 1693479267
transform 1 0 2412 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_351
timestamp 1693479267
transform -1 0 2468 0 1 1705
box -2 -3 26 103
use AND2X2  AND2X2_26
timestamp 1693479267
transform -1 0 2500 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_347
timestamp 1693479267
transform 1 0 2500 0 1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_314
timestamp 1693479267
transform 1 0 2516 0 1 1705
box -2 -3 26 103
use FILL  FILL_17_4_0
timestamp 1693479267
transform -1 0 2548 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_4_1
timestamp 1693479267
transform -1 0 2556 0 1 1705
box -2 -3 10 103
use NOR2X1  NOR2X1_262
timestamp 1693479267
transform -1 0 2580 0 1 1705
box -2 -3 26 103
use AOI22X1  AOI22X1_93
timestamp 1693479267
transform -1 0 2620 0 1 1705
box -2 -3 42 103
use AOI21X1  AOI21X1_44
timestamp 1693479267
transform -1 0 2652 0 1 1705
box -2 -3 34 103
use AOI22X1  AOI22X1_94
timestamp 1693479267
transform -1 0 2692 0 1 1705
box -2 -3 42 103
use AOI21X1  AOI21X1_49
timestamp 1693479267
transform 1 0 2692 0 1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_55
timestamp 1693479267
transform 1 0 2724 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_377
timestamp 1693479267
transform 1 0 2756 0 1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_185
timestamp 1693479267
transform -1 0 2796 0 1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_183
timestamp 1693479267
transform 1 0 2796 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_340
timestamp 1693479267
transform 1 0 2820 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_264
timestamp 1693479267
transform -1 0 2876 0 1 1705
box -2 -3 26 103
use OR2X2  OR2X2_31
timestamp 1693479267
transform 1 0 2876 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_348
timestamp 1693479267
transform 1 0 2908 0 1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_493
timestamp 1693479267
transform 1 0 2924 0 1 1705
box -2 -3 26 103
use AND2X2  AND2X2_43
timestamp 1693479267
transform 1 0 2948 0 1 1705
box -2 -3 34 103
use OAI22X1  OAI22X1_25
timestamp 1693479267
transform 1 0 2980 0 1 1705
box -2 -3 42 103
use AOI21X1  AOI21X1_106
timestamp 1693479267
transform -1 0 3052 0 1 1705
box -2 -3 34 103
use FILL  FILL_17_5_0
timestamp 1693479267
transform -1 0 3060 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_5_1
timestamp 1693479267
transform -1 0 3068 0 1 1705
box -2 -3 10 103
use AOI21X1  AOI21X1_105
timestamp 1693479267
transform -1 0 3100 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_391
timestamp 1693479267
transform -1 0 3116 0 1 1705
box -2 -3 18 103
use NAND3X1  NAND3X1_128
timestamp 1693479267
transform -1 0 3148 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_338
timestamp 1693479267
transform 1 0 3148 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_360
timestamp 1693479267
transform -1 0 3204 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_410
timestamp 1693479267
transform 1 0 3204 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_706
timestamp 1693479267
transform 1 0 3236 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_699
timestamp 1693479267
transform 1 0 3268 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_573
timestamp 1693479267
transform -1 0 3324 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_387
timestamp 1693479267
transform -1 0 3356 0 1 1705
box -2 -3 34 103
use INVX2  INVX2_50
timestamp 1693479267
transform -1 0 3372 0 1 1705
box -2 -3 18 103
use INVX1  INVX1_363
timestamp 1693479267
transform 1 0 3372 0 1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_574
timestamp 1693479267
transform -1 0 3412 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_725
timestamp 1693479267
transform 1 0 3412 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_584
timestamp 1693479267
transform -1 0 3468 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_594
timestamp 1693479267
transform -1 0 3492 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_746
timestamp 1693479267
transform -1 0 3524 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_452
timestamp 1693479267
transform -1 0 3548 0 1 1705
box -2 -3 26 103
use AND2X2  AND2X2_28
timestamp 1693479267
transform -1 0 3580 0 1 1705
box -2 -3 34 103
use FILL  FILL_17_6_0
timestamp 1693479267
transform 1 0 3580 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_6_1
timestamp 1693479267
transform 1 0 3588 0 1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_766
timestamp 1693479267
transform 1 0 3596 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_372
timestamp 1693479267
transform -1 0 3652 0 1 1705
box -2 -3 26 103
use OAI22X1  OAI22X1_44
timestamp 1693479267
transform 1 0 3652 0 1 1705
box -2 -3 42 103
use OAI21X1  OAI21X1_436
timestamp 1693479267
transform 1 0 3692 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_418
timestamp 1693479267
transform 1 0 3724 0 1 1705
box -2 -3 26 103
use AND2X2  AND2X2_73
timestamp 1693479267
transform 1 0 3748 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_440
timestamp 1693479267
transform -1 0 3812 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_589
timestamp 1693479267
transform -1 0 3836 0 1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_235
timestamp 1693479267
transform -1 0 3860 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_366
timestamp 1693479267
transform -1 0 3884 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_380
timestamp 1693479267
transform 1 0 3884 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_707
timestamp 1693479267
transform -1 0 3948 0 1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_183
timestamp 1693479267
transform -1 0 3980 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_93
timestamp 1693479267
transform 1 0 3980 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_276
timestamp 1693479267
transform 1 0 4012 0 1 1705
box -2 -3 34 103
use AND2X2  AND2X2_70
timestamp 1693479267
transform 1 0 4044 0 1 1705
box -2 -3 34 103
use FILL  FILL_17_7_0
timestamp 1693479267
transform -1 0 4084 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_7_1
timestamp 1693479267
transform -1 0 4092 0 1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_720
timestamp 1693479267
transform -1 0 4124 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_77
timestamp 1693479267
transform 1 0 4124 0 1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_79
timestamp 1693479267
transform 1 0 4148 0 1 1705
box -2 -3 26 103
use AOI22X1  AOI22X1_104
timestamp 1693479267
transform 1 0 4172 0 1 1705
box -2 -3 42 103
use AOI22X1  AOI22X1_105
timestamp 1693479267
transform -1 0 4252 0 1 1705
box -2 -3 42 103
use OAI22X1  OAI22X1_41
timestamp 1693479267
transform 1 0 4252 0 1 1705
box -2 -3 42 103
use NOR2X1  NOR2X1_361
timestamp 1693479267
transform 1 0 4292 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_599
timestamp 1693479267
transform 1 0 4316 0 1 1705
box -2 -3 26 103
use OAI22X1  OAI22X1_43
timestamp 1693479267
transform 1 0 4340 0 1 1705
box -2 -3 42 103
use OAI21X1  OAI21X1_749
timestamp 1693479267
transform 1 0 4380 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_596
timestamp 1693479267
transform -1 0 4436 0 1 1705
box -2 -3 26 103
use NAND3X1  NAND3X1_167
timestamp 1693479267
transform -1 0 4468 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_735
timestamp 1693479267
transform -1 0 4500 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_587
timestamp 1693479267
transform -1 0 4524 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_729
timestamp 1693479267
transform -1 0 4556 0 1 1705
box -2 -3 34 103
use INVX2  INVX2_18
timestamp 1693479267
transform -1 0 4572 0 1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_74
timestamp 1693479267
transform 1 0 4572 0 1 1705
box -2 -3 26 103
use FILL  FILL_18_1
timestamp 1693479267
transform 1 0 4596 0 1 1705
box -2 -3 10 103
use BUFX2  BUFX2_68
timestamp 1693479267
transform -1 0 28 0 -1 1905
box -2 -3 26 103
use BUFX2  BUFX2_3
timestamp 1693479267
transform -1 0 52 0 -1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_160
timestamp 1693479267
transform -1 0 148 0 -1 1905
box -2 -3 98 103
use CLKBUF1  CLKBUF1_5
timestamp 1693479267
transform -1 0 220 0 -1 1905
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_441
timestamp 1693479267
transform 1 0 220 0 -1 1905
box -2 -3 98 103
use INVX1  INVX1_489
timestamp 1693479267
transform -1 0 332 0 -1 1905
box -2 -3 18 103
use INVX1  INVX1_488
timestamp 1693479267
transform -1 0 348 0 -1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_865
timestamp 1693479267
transform 1 0 348 0 -1 1905
box -2 -3 34 103
use INVX8  INVX8_1
timestamp 1693479267
transform 1 0 380 0 -1 1905
box -2 -3 42 103
use OAI21X1  OAI21X1_188
timestamp 1693479267
transform -1 0 452 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_61
timestamp 1693479267
transform -1 0 484 0 -1 1905
box -2 -3 34 103
use FILL  FILL_18_0_0
timestamp 1693479267
transform 1 0 484 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_0_1
timestamp 1693479267
transform 1 0 492 0 -1 1905
box -2 -3 10 103
use XOR2X1  XOR2X1_9
timestamp 1693479267
transform 1 0 500 0 -1 1905
box -2 -3 58 103
use OAI21X1  OAI21X1_859
timestamp 1693479267
transform 1 0 556 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_187
timestamp 1693479267
transform -1 0 620 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_190
timestamp 1693479267
transform -1 0 652 0 -1 1905
box -2 -3 34 103
use BUFX4  BUFX4_13
timestamp 1693479267
transform -1 0 684 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_497
timestamp 1693479267
transform 1 0 684 0 -1 1905
box -2 -3 98 103
use NAND3X1  NAND3X1_65
timestamp 1693479267
transform 1 0 780 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_501
timestamp 1693479267
transform 1 0 812 0 -1 1905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_469
timestamp 1693479267
transform 1 0 908 0 -1 1905
box -2 -3 98 103
use FILL  FILL_18_1_0
timestamp 1693479267
transform 1 0 1004 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_1_1
timestamp 1693479267
transform 1 0 1012 0 -1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_283
timestamp 1693479267
transform 1 0 1020 0 -1 1905
box -2 -3 98 103
use INVX1  INVX1_294
timestamp 1693479267
transform 1 0 1116 0 -1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_64
timestamp 1693479267
transform -1 0 1156 0 -1 1905
box -2 -3 26 103
use INVX1  INVX1_290
timestamp 1693479267
transform 1 0 1156 0 -1 1905
box -2 -3 18 103
use AOI21X1  AOI21X1_32
timestamp 1693479267
transform -1 0 1204 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_59
timestamp 1693479267
transform 1 0 1204 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_275
timestamp 1693479267
transform -1 0 1260 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_278
timestamp 1693479267
transform 1 0 1260 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_292
timestamp 1693479267
transform 1 0 1292 0 -1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_63
timestamp 1693479267
transform -1 0 1332 0 -1 1905
box -2 -3 26 103
use NAND3X1  NAND3X1_87
timestamp 1693479267
transform 1 0 1332 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_300
timestamp 1693479267
transform -1 0 1380 0 -1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_62
timestamp 1693479267
transform 1 0 1380 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_189
timestamp 1693479267
transform -1 0 1428 0 -1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_284
timestamp 1693479267
transform 1 0 1428 0 -1 1905
box -2 -3 98 103
use FILL  FILL_18_2_0
timestamp 1693479267
transform 1 0 1524 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_2_1
timestamp 1693479267
transform 1 0 1532 0 -1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_302
timestamp 1693479267
transform 1 0 1540 0 -1 1905
box -2 -3 98 103
use XNOR2X1  XNOR2X1_48
timestamp 1693479267
transform -1 0 1692 0 -1 1905
box -2 -3 58 103
use AND2X2  AND2X2_12
timestamp 1693479267
transform -1 0 1724 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_291
timestamp 1693479267
transform -1 0 1740 0 -1 1905
box -2 -3 18 103
use AOI22X1  AOI22X1_66
timestamp 1693479267
transform 1 0 1740 0 -1 1905
box -2 -3 42 103
use AOI22X1  AOI22X1_68
timestamp 1693479267
transform 1 0 1780 0 -1 1905
box -2 -3 42 103
use NOR3X1  NOR3X1_48
timestamp 1693479267
transform -1 0 1884 0 -1 1905
box -2 -3 66 103
use INVX1  INVX1_238
timestamp 1693479267
transform 1 0 1884 0 -1 1905
box -2 -3 18 103
use NAND2X1  NAND2X1_126
timestamp 1693479267
transform -1 0 1924 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_204
timestamp 1693479267
transform -1 0 1948 0 -1 1905
box -2 -3 26 103
use INVX1  INVX1_236
timestamp 1693479267
transform 1 0 1948 0 -1 1905
box -2 -3 18 103
use NOR3X1  NOR3X1_47
timestamp 1693479267
transform 1 0 1964 0 -1 1905
box -2 -3 66 103
use FILL  FILL_18_3_0
timestamp 1693479267
transform -1 0 2036 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_3_1
timestamp 1693479267
transform -1 0 2044 0 -1 1905
box -2 -3 10 103
use INVX1  INVX1_237
timestamp 1693479267
transform -1 0 2060 0 -1 1905
box -2 -3 18 103
use NAND2X1  NAND2X1_194
timestamp 1693479267
transform -1 0 2084 0 -1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_379
timestamp 1693479267
transform -1 0 2108 0 -1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_71
timestamp 1693479267
transform 1 0 2108 0 -1 1905
box -2 -3 26 103
use OR2X2  OR2X2_44
timestamp 1693479267
transform 1 0 2132 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_199
timestamp 1693479267
transform -1 0 2188 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_203
timestamp 1693479267
transform -1 0 2212 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_371
timestamp 1693479267
transform -1 0 2244 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_102
timestamp 1693479267
transform 1 0 2244 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_350
timestamp 1693479267
transform -1 0 2300 0 -1 1905
box -2 -3 26 103
use AND2X2  AND2X2_25
timestamp 1693479267
transform -1 0 2332 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_174
timestamp 1693479267
transform 1 0 2332 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_348
timestamp 1693479267
transform -1 0 2380 0 -1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_175
timestamp 1693479267
transform -1 0 2404 0 -1 1905
box -2 -3 26 103
use INVX1  INVX1_359
timestamp 1693479267
transform 1 0 2404 0 -1 1905
box -2 -3 18 103
use NAND2X1  NAND2X1_354
timestamp 1693479267
transform 1 0 2420 0 -1 1905
box -2 -3 26 103
use MUX2X1  MUX2X1_13
timestamp 1693479267
transform -1 0 2492 0 -1 1905
box -2 -3 50 103
use AOI21X1  AOI21X1_236
timestamp 1693479267
transform -1 0 2524 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_984
timestamp 1693479267
transform 1 0 2524 0 -1 1905
box -2 -3 26 103
use FILL  FILL_18_4_0
timestamp 1693479267
transform 1 0 2548 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_4_1
timestamp 1693479267
transform 1 0 2556 0 -1 1905
box -2 -3 10 103
use INVX1  INVX1_688
timestamp 1693479267
transform 1 0 2564 0 -1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_435
timestamp 1693479267
transform -1 0 2604 0 -1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_135
timestamp 1693479267
transform -1 0 2628 0 -1 1905
box -2 -3 26 103
use INVX1  INVX1_390
timestamp 1693479267
transform 1 0 2628 0 -1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_257
timestamp 1693479267
transform -1 0 2668 0 -1 1905
box -2 -3 26 103
use NAND3X1  NAND3X1_125
timestamp 1693479267
transform -1 0 2700 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_126
timestamp 1693479267
transform 1 0 2700 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_356
timestamp 1693479267
transform -1 0 2748 0 -1 1905
box -2 -3 18 103
use NAND2X1  NAND2X1_344
timestamp 1693479267
transform -1 0 2772 0 -1 1905
box -2 -3 26 103
use INVX1  INVX1_376
timestamp 1693479267
transform 1 0 2772 0 -1 1905
box -2 -3 18 103
use INVX2  INVX2_56
timestamp 1693479267
transform -1 0 2804 0 -1 1905
box -2 -3 18 103
use NAND2X1  NAND2X1_435
timestamp 1693479267
transform 1 0 2804 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_462
timestamp 1693479267
transform 1 0 2828 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_355
timestamp 1693479267
transform -1 0 2884 0 -1 1905
box -2 -3 26 103
use INVX2  INVX2_49
timestamp 1693479267
transform 1 0 2884 0 -1 1905
box -2 -3 18 103
use INVX1  INVX1_352
timestamp 1693479267
transform 1 0 2900 0 -1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_136
timestamp 1693479267
transform -1 0 2940 0 -1 1905
box -2 -3 26 103
use NAND3X1  NAND3X1_92
timestamp 1693479267
transform -1 0 2972 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_978
timestamp 1693479267
transform 1 0 2972 0 -1 1905
box -2 -3 26 103
use INVX1  INVX1_672
timestamp 1693479267
transform 1 0 2996 0 -1 1905
box -2 -3 18 103
use NAND2X1  NAND2X1_941
timestamp 1693479267
transform 1 0 3012 0 -1 1905
box -2 -3 26 103
use INVX1  INVX1_673
timestamp 1693479267
transform -1 0 3052 0 -1 1905
box -2 -3 18 103
use FILL  FILL_18_5_0
timestamp 1693479267
transform 1 0 3052 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_5_1
timestamp 1693479267
transform 1 0 3060 0 -1 1905
box -2 -3 10 103
use BUFX4  BUFX4_188
timestamp 1693479267
transform 1 0 3068 0 -1 1905
box -2 -3 34 103
use BUFX4  BUFX4_88
timestamp 1693479267
transform 1 0 3100 0 -1 1905
box -2 -3 34 103
use INVX8  INVX8_12
timestamp 1693479267
transform -1 0 3172 0 -1 1905
box -2 -3 42 103
use OAI21X1  OAI21X1_285
timestamp 1693479267
transform -1 0 3204 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_409
timestamp 1693479267
transform -1 0 3236 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_158
timestamp 1693479267
transform 1 0 3236 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_357
timestamp 1693479267
transform 1 0 3260 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_159
timestamp 1693479267
transform 1 0 3292 0 -1 1905
box -2 -3 26 103
use INVX1  INVX1_421
timestamp 1693479267
transform 1 0 3316 0 -1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_358
timestamp 1693479267
transform -1 0 3364 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_408
timestamp 1693479267
transform 1 0 3364 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_395
timestamp 1693479267
transform 1 0 3396 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_745
timestamp 1693479267
transform 1 0 3420 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_355
timestamp 1693479267
transform -1 0 3484 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_765
timestamp 1693479267
transform 1 0 3484 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_356
timestamp 1693479267
transform -1 0 3548 0 -1 1905
box -2 -3 34 103
use FILL  FILL_18_6_0
timestamp 1693479267
transform 1 0 3548 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_6_1
timestamp 1693479267
transform 1 0 3556 0 -1 1905
box -2 -3 10 103
use MUX2X1  MUX2X1_48
timestamp 1693479267
transform 1 0 3564 0 -1 1905
box -2 -3 50 103
use INVX1  INVX1_361
timestamp 1693479267
transform 1 0 3612 0 -1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_381
timestamp 1693479267
transform 1 0 3628 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_382
timestamp 1693479267
transform -1 0 3692 0 -1 1905
box -2 -3 34 103
use OR2X2  OR2X2_25
timestamp 1693479267
transform -1 0 3724 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_439
timestamp 1693479267
transform 1 0 3724 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_379
timestamp 1693479267
transform 1 0 3756 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_736
timestamp 1693479267
transform -1 0 3820 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_80
timestamp 1693479267
transform -1 0 3844 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_200
timestamp 1693479267
transform -1 0 3868 0 -1 1905
box -2 -3 26 103
use INVX1  INVX1_416
timestamp 1693479267
transform 1 0 3868 0 -1 1905
box -2 -3 18 103
use NAND2X1  NAND2X1_319
timestamp 1693479267
transform 1 0 3884 0 -1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_343
timestamp 1693479267
transform -1 0 3932 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_335
timestamp 1693479267
transform 1 0 3932 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_194
timestamp 1693479267
transform 1 0 3964 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_349
timestamp 1693479267
transform -1 0 4020 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_318
timestamp 1693479267
transform -1 0 4044 0 -1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_78
timestamp 1693479267
transform -1 0 4068 0 -1 1905
box -2 -3 26 103
use INVX1  INVX1_307
timestamp 1693479267
transform -1 0 4084 0 -1 1905
box -2 -3 18 103
use FILL  FILL_18_7_0
timestamp 1693479267
transform -1 0 4092 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_7_1
timestamp 1693479267
transform -1 0 4100 0 -1 1905
box -2 -3 10 103
use NOR2X1  NOR2X1_163
timestamp 1693479267
transform -1 0 4124 0 -1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_190
timestamp 1693479267
transform 1 0 4124 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_96
timestamp 1693479267
transform -1 0 4188 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_303
timestamp 1693479267
transform -1 0 4204 0 -1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_75
timestamp 1693479267
transform 1 0 4204 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_317
timestamp 1693479267
transform 1 0 4228 0 -1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_195
timestamp 1693479267
transform 1 0 4252 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_283
timestamp 1693479267
transform 1 0 4284 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_422
timestamp 1693479267
transform 1 0 4316 0 -1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_741
timestamp 1693479267
transform -1 0 4364 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_166
timestamp 1693479267
transform 1 0 4364 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_593
timestamp 1693479267
transform 1 0 4396 0 -1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_199
timestamp 1693479267
transform 1 0 4420 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_196
timestamp 1693479267
transform -1 0 4484 0 -1 1905
box -2 -3 34 103
use INVX2  INVX2_17
timestamp 1693479267
transform 1 0 4484 0 -1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_354
timestamp 1693479267
transform -1 0 4524 0 -1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_73
timestamp 1693479267
transform -1 0 4548 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_734
timestamp 1693479267
transform 1 0 4548 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_72
timestamp 1693479267
transform 1 0 4580 0 -1 1905
box -2 -3 26 103
use BUFX2  BUFX2_29
timestamp 1693479267
transform -1 0 28 0 1 1905
box -2 -3 26 103
use BUFX2  BUFX2_64
timestamp 1693479267
transform -1 0 52 0 1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_186
timestamp 1693479267
transform -1 0 148 0 1 1905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_187
timestamp 1693479267
transform -1 0 244 0 1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_862
timestamp 1693479267
transform 1 0 244 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_691
timestamp 1693479267
transform -1 0 300 0 1 1905
box -2 -3 26 103
use NAND3X1  NAND3X1_9
timestamp 1693479267
transform 1 0 300 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_688
timestamp 1693479267
transform -1 0 356 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_692
timestamp 1693479267
transform 1 0 356 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_189
timestamp 1693479267
transform -1 0 412 0 1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_500
timestamp 1693479267
transform -1 0 508 0 1 1905
box -2 -3 98 103
use FILL  FILL_19_0_0
timestamp 1693479267
transform -1 0 516 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_0_1
timestamp 1693479267
transform -1 0 524 0 1 1905
box -2 -3 10 103
use NAND3X1  NAND3X1_63
timestamp 1693479267
transform -1 0 556 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_858
timestamp 1693479267
transform 1 0 556 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_687
timestamp 1693479267
transform 1 0 588 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_186
timestamp 1693479267
transform -1 0 644 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_57
timestamp 1693479267
transform -1 0 676 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_56
timestamp 1693479267
transform -1 0 708 0 1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_465
timestamp 1693479267
transform 1 0 708 0 1 1905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_255
timestamp 1693479267
transform 1 0 804 0 1 1905
box -2 -3 98 103
use CLKBUF1  CLKBUF1_36
timestamp 1693479267
transform 1 0 900 0 1 1905
box -2 -3 74 103
use XNOR2X1  XNOR2X1_47
timestamp 1693479267
transform 1 0 972 0 1 1905
box -2 -3 58 103
use FILL  FILL_19_1_0
timestamp 1693479267
transform 1 0 1028 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_1_1
timestamp 1693479267
transform 1 0 1036 0 1 1905
box -2 -3 10 103
use NOR2X1  NOR2X1_61
timestamp 1693479267
transform 1 0 1044 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_60
timestamp 1693479267
transform 1 0 1068 0 1 1905
box -2 -3 26 103
use AND2X2  AND2X2_17
timestamp 1693479267
transform -1 0 1124 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_289
timestamp 1693479267
transform 1 0 1124 0 1 1905
box -2 -3 18 103
use AOI21X1  AOI21X1_31
timestamp 1693479267
transform -1 0 1172 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_187
timestamp 1693479267
transform -1 0 1196 0 1 1905
box -2 -3 26 103
use AND2X2  AND2X2_19
timestamp 1693479267
transform -1 0 1228 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_190
timestamp 1693479267
transform -1 0 1252 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_65
timestamp 1693479267
transform -1 0 1276 0 1 1905
box -2 -3 26 103
use INVX1  INVX1_297
timestamp 1693479267
transform 1 0 1276 0 1 1905
box -2 -3 18 103
use INVX1  INVX1_274
timestamp 1693479267
transform 1 0 1292 0 1 1905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_279
timestamp 1693479267
transform 1 0 1308 0 1 1905
box -2 -3 98 103
use XNOR2X1  XNOR2X1_5
timestamp 1693479267
transform 1 0 1404 0 1 1905
box -2 -3 58 103
use AOI21X1  AOI21X1_6
timestamp 1693479267
transform 1 0 1460 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_121
timestamp 1693479267
transform 1 0 1492 0 1 1905
box -2 -3 26 103
use FILL  FILL_19_2_0
timestamp 1693479267
transform 1 0 1516 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_2_1
timestamp 1693479267
transform 1 0 1524 0 1 1905
box -2 -3 10 103
use NOR2X1  NOR2X1_26
timestamp 1693479267
transform 1 0 1532 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_120
timestamp 1693479267
transform -1 0 1580 0 1 1905
box -2 -3 26 103
use OR2X2  OR2X2_9
timestamp 1693479267
transform 1 0 1580 0 1 1905
box -2 -3 34 103
use AND2X2  AND2X2_13
timestamp 1693479267
transform 1 0 1612 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_230
timestamp 1693479267
transform -1 0 1676 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_229
timestamp 1693479267
transform -1 0 1708 0 1 1905
box -2 -3 34 103
use AND2X2  AND2X2_11
timestamp 1693479267
transform -1 0 1740 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_148
timestamp 1693479267
transform 1 0 1740 0 1 1905
box -2 -3 34 103
use AOI22X1  AOI22X1_42
timestamp 1693479267
transform 1 0 1772 0 1 1905
box -2 -3 42 103
use AOI22X1  AOI22X1_63
timestamp 1693479267
transform -1 0 1852 0 1 1905
box -2 -3 42 103
use AOI22X1  AOI22X1_67
timestamp 1693479267
transform -1 0 1892 0 1 1905
box -2 -3 42 103
use NAND2X1  NAND2X1_125
timestamp 1693479267
transform -1 0 1916 0 1 1905
box -2 -3 26 103
use AND2X2  AND2X2_9
timestamp 1693479267
transform -1 0 1948 0 1 1905
box -2 -3 34 103
use AND2X2  AND2X2_20
timestamp 1693479267
transform 1 0 1948 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_205
timestamp 1693479267
transform -1 0 2004 0 1 1905
box -2 -3 26 103
use INVX1  INVX1_314
timestamp 1693479267
transform 1 0 2004 0 1 1905
box -2 -3 18 103
use FILL  FILL_19_3_0
timestamp 1693479267
transform 1 0 2020 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_3_1
timestamp 1693479267
transform 1 0 2028 0 1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_290
timestamp 1693479267
transform 1 0 2036 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_289
timestamp 1693479267
transform -1 0 2100 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_313
timestamp 1693479267
transform -1 0 2116 0 1 1905
box -2 -3 18 103
use NAND2X1  NAND2X1_196
timestamp 1693479267
transform -1 0 2140 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_281
timestamp 1693479267
transform -1 0 2172 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_302
timestamp 1693479267
transform -1 0 2188 0 1 1905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_349
timestamp 1693479267
transform 1 0 2188 0 1 1905
box -2 -3 98 103
use NAND2X1  NAND2X1_198
timestamp 1693479267
transform -1 0 2308 0 1 1905
box -2 -3 26 103
use OR2X2  OR2X2_61
timestamp 1693479267
transform 1 0 2308 0 1 1905
box -2 -3 34 103
use AOI22X1  AOI22X1_131
timestamp 1693479267
transform -1 0 2380 0 1 1905
box -2 -3 42 103
use NAND2X1  NAND2X1_954
timestamp 1693479267
transform -1 0 2404 0 1 1905
box -2 -3 26 103
use OR2X2  OR2X2_60
timestamp 1693479267
transform -1 0 2436 0 1 1905
box -2 -3 34 103
use INVX2  INVX2_85
timestamp 1693479267
transform 1 0 2436 0 1 1905
box -2 -3 18 103
use INVX2  INVX2_48
timestamp 1693479267
transform 1 0 2452 0 1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_436
timestamp 1693479267
transform -1 0 2492 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_962
timestamp 1693479267
transform 1 0 2492 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_928
timestamp 1693479267
transform 1 0 2516 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_4_0
timestamp 1693479267
transform 1 0 2548 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_4_1
timestamp 1693479267
transform 1 0 2556 0 1 1905
box -2 -3 10 103
use INVX1  INVX1_355
timestamp 1693479267
transform 1 0 2564 0 1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_172
timestamp 1693479267
transform -1 0 2604 0 1 1905
box -2 -3 26 103
use AND2X2  AND2X2_23
timestamp 1693479267
transform 1 0 2604 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_315
timestamp 1693479267
transform -1 0 2660 0 1 1905
box -2 -3 26 103
use INVX1  INVX1_686
timestamp 1693479267
transform 1 0 2660 0 1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_284
timestamp 1693479267
transform -1 0 2708 0 1 1905
box -2 -3 34 103
use AND2X2  AND2X2_94
timestamp 1693479267
transform 1 0 2708 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_687
timestamp 1693479267
transform 1 0 2740 0 1 1905
box -2 -3 18 103
use OR2X2  OR2X2_65
timestamp 1693479267
transform 1 0 2756 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_927
timestamp 1693479267
transform 1 0 2788 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_708
timestamp 1693479267
transform -1 0 2836 0 1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_433
timestamp 1693479267
transform -1 0 2860 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_434
timestamp 1693479267
transform -1 0 2884 0 1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_234
timestamp 1693479267
transform -1 0 2916 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_960
timestamp 1693479267
transform -1 0 2940 0 1 1905
box -2 -3 26 103
use INVX1  INVX1_701
timestamp 1693479267
transform 1 0 2940 0 1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_448
timestamp 1693479267
transform -1 0 2980 0 1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_241
timestamp 1693479267
transform 1 0 2980 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_449
timestamp 1693479267
transform -1 0 3036 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_940
timestamp 1693479267
transform 1 0 3036 0 1 1905
box -2 -3 26 103
use FILL  FILL_19_5_0
timestamp 1693479267
transform -1 0 3068 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_5_1
timestamp 1693479267
transform -1 0 3076 0 1 1905
box -2 -3 10 103
use AOI22X1  AOI22X1_128
timestamp 1693479267
transform -1 0 3116 0 1 1905
box -2 -3 42 103
use OR2X2  OR2X2_56
timestamp 1693479267
transform -1 0 3148 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_942
timestamp 1693479267
transform 1 0 3148 0 1 1905
box -2 -3 26 103
use INVX1  INVX1_711
timestamp 1693479267
transform 1 0 3172 0 1 1905
box -2 -3 18 103
use AND2X2  AND2X2_21
timestamp 1693479267
transform 1 0 3188 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_338
timestamp 1693479267
transform -1 0 3252 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_38
timestamp 1693479267
transform 1 0 3252 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_583
timestamp 1693479267
transform 1 0 3284 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_724
timestamp 1693479267
transform -1 0 3340 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_53
timestamp 1693479267
transform 1 0 3340 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_40
timestamp 1693479267
transform 1 0 3372 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_157
timestamp 1693479267
transform 1 0 3404 0 1 1905
box -2 -3 26 103
use INVX4  INVX4_3
timestamp 1693479267
transform 1 0 3428 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_334
timestamp 1693479267
transform -1 0 3476 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_335
timestamp 1693479267
transform 1 0 3476 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_421
timestamp 1693479267
transform 1 0 3500 0 1 1905
box -2 -3 26 103
use INVX2  INVX2_25
timestamp 1693479267
transform 1 0 3524 0 1 1905
box -2 -3 18 103
use INVX4  INVX4_2
timestamp 1693479267
transform -1 0 3564 0 1 1905
box -2 -3 26 103
use FILL  FILL_19_6_0
timestamp 1693479267
transform 1 0 3564 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_6_1
timestamp 1693479267
transform 1 0 3572 0 1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_378
timestamp 1693479267
transform 1 0 3580 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_364
timestamp 1693479267
transform -1 0 3636 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_189
timestamp 1693479267
transform 1 0 3636 0 1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_205
timestamp 1693479267
transform 1 0 3660 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_165
timestamp 1693479267
transform -1 0 3724 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_190
timestamp 1693479267
transform 1 0 3724 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_365
timestamp 1693479267
transform 1 0 3748 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_81
timestamp 1693479267
transform 1 0 3772 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_713
timestamp 1693479267
transform 1 0 3796 0 1 1905
box -2 -3 34 103
use INVX2  INVX2_19
timestamp 1693479267
transform -1 0 3844 0 1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_709
timestamp 1693479267
transform 1 0 3844 0 1 1905
box -2 -3 34 103
use AND2X2  AND2X2_65
timestamp 1693479267
transform -1 0 3908 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_419
timestamp 1693479267
transform -1 0 3924 0 1 1905
box -2 -3 18 103
use AOI21X1  AOI21X1_187
timestamp 1693479267
transform 1 0 3924 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_714
timestamp 1693479267
transform 1 0 3956 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_732
timestamp 1693479267
transform 1 0 3988 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_733
timestamp 1693479267
transform 1 0 4020 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_191
timestamp 1693479267
transform 1 0 4052 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_7_0
timestamp 1693479267
transform 1 0 4084 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_7_1
timestamp 1693479267
transform 1 0 4092 0 1 1905
box -2 -3 10 103
use NOR2X1  NOR2X1_350
timestamp 1693479267
transform 1 0 4100 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_82
timestamp 1693479267
transform 1 0 4124 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_578
timestamp 1693479267
transform 1 0 4148 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_201
timestamp 1693479267
transform 1 0 4172 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_76
timestamp 1693479267
transform -1 0 4220 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_139
timestamp 1693479267
transform 1 0 4220 0 1 1905
box -2 -3 26 103
use AOI22X1  AOI22X1_75
timestamp 1693479267
transform -1 0 4284 0 1 1905
box -2 -3 42 103
use INVX1  INVX1_349
timestamp 1693479267
transform -1 0 4300 0 1 1905
box -2 -3 18 103
use INVX1  INVX1_305
timestamp 1693479267
transform -1 0 4316 0 1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_750
timestamp 1693479267
transform 1 0 4316 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_202
timestamp 1693479267
transform -1 0 4380 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_334
timestamp 1693479267
transform -1 0 4412 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_355
timestamp 1693479267
transform -1 0 4436 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_592
timestamp 1693479267
transform -1 0 4460 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_351
timestamp 1693479267
transform -1 0 4484 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_723
timestamp 1693479267
transform 1 0 4484 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_192
timestamp 1693479267
transform -1 0 4548 0 1 1905
box -2 -3 34 103
use INVX2  INVX2_16
timestamp 1693479267
transform 1 0 4548 0 1 1905
box -2 -3 18 103
use NAND2X1  NAND2X1_588
timestamp 1693479267
transform -1 0 4588 0 1 1905
box -2 -3 26 103
use FILL  FILL_20_1
timestamp 1693479267
transform 1 0 4588 0 1 1905
box -2 -3 10 103
use FILL  FILL_20_2
timestamp 1693479267
transform 1 0 4596 0 1 1905
box -2 -3 10 103
use BUFX2  BUFX2_40
timestamp 1693479267
transform -1 0 28 0 -1 2105
box -2 -3 26 103
use BUFX2  BUFX2_27
timestamp 1693479267
transform -1 0 52 0 -1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_184
timestamp 1693479267
transform -1 0 148 0 -1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_473
timestamp 1693479267
transform -1 0 244 0 -1 2105
box -2 -3 98 103
use INVX1  INVX1_469
timestamp 1693479267
transform 1 0 244 0 -1 2105
box -2 -3 18 103
use AOI21X1  AOI21X1_2
timestamp 1693479267
transform -1 0 292 0 -1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_1
timestamp 1693479267
transform -1 0 324 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_8
timestamp 1693479267
transform 1 0 324 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_816
timestamp 1693479267
transform 1 0 356 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_162
timestamp 1693479267
transform -1 0 420 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_161
timestamp 1693479267
transform 1 0 420 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_60
timestamp 1693479267
transform -1 0 484 0 -1 2105
box -2 -3 34 103
use FILL  FILL_20_0_0
timestamp 1693479267
transform -1 0 492 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_0_1
timestamp 1693479267
transform -1 0 500 0 -1 2105
box -2 -3 10 103
use NAND3X1  NAND3X1_62
timestamp 1693479267
transform -1 0 532 0 -1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_468
timestamp 1693479267
transform 1 0 532 0 -1 2105
box -2 -3 98 103
use BUFX4  BUFX4_112
timestamp 1693479267
transform -1 0 660 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_640
timestamp 1693479267
transform 1 0 660 0 -1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_281
timestamp 1693479267
transform 1 0 684 0 -1 2105
box -2 -3 98 103
use INVX1  INVX1_663
timestamp 1693479267
transform 1 0 780 0 -1 2105
box -2 -3 18 103
use NAND3X1  NAND3X1_328
timestamp 1693479267
transform -1 0 828 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_902
timestamp 1693479267
transform 1 0 828 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_662
timestamp 1693479267
transform -1 0 876 0 -1 2105
box -2 -3 18 103
use NAND3X1  NAND3X1_329
timestamp 1693479267
transform 1 0 876 0 -1 2105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_46
timestamp 1693479267
transform 1 0 908 0 -1 2105
box -2 -3 58 103
use NAND2X1  NAND2X1_184
timestamp 1693479267
transform -1 0 988 0 -1 2105
box -2 -3 26 103
use INVX1  INVX1_284
timestamp 1693479267
transform -1 0 1004 0 -1 2105
box -2 -3 18 103
use FILL  FILL_20_1_0
timestamp 1693479267
transform 1 0 1004 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_1_1
timestamp 1693479267
transform 1 0 1012 0 -1 2105
box -2 -3 10 103
use AOI21X1  AOI21X1_30
timestamp 1693479267
transform 1 0 1020 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_183
timestamp 1693479267
transform -1 0 1076 0 -1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_55
timestamp 1693479267
transform 1 0 1076 0 -1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_57
timestamp 1693479267
transform 1 0 1100 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_274
timestamp 1693479267
transform 1 0 1124 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_281
timestamp 1693479267
transform 1 0 1156 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_272
timestamp 1693479267
transform -1 0 1204 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_282
timestamp 1693479267
transform -1 0 1220 0 -1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_54
timestamp 1693479267
transform -1 0 1244 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_270
timestamp 1693479267
transform 1 0 1244 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_296
timestamp 1693479267
transform 1 0 1276 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_271
timestamp 1693479267
transform 1 0 1292 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_180
timestamp 1693479267
transform -1 0 1348 0 -1 2105
box -2 -3 26 103
use INVX2  INVX2_15
timestamp 1693479267
transform -1 0 1364 0 -1 2105
box -2 -3 18 103
use NAND2X1  NAND2X1_179
timestamp 1693479267
transform -1 0 1388 0 -1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_52
timestamp 1693479267
transform -1 0 1412 0 -1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_254
timestamp 1693479267
transform 1 0 1412 0 -1 2105
box -2 -3 98 103
use NOR2X1  NOR2X1_69
timestamp 1693479267
transform 1 0 1508 0 -1 2105
box -2 -3 26 103
use FILL  FILL_20_2_0
timestamp 1693479267
transform -1 0 1540 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_2_1
timestamp 1693479267
transform -1 0 1548 0 -1 2105
box -2 -3 10 103
use NOR2X1  NOR2X1_68
timestamp 1693479267
transform -1 0 1572 0 -1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_193
timestamp 1693479267
transform -1 0 1596 0 -1 2105
box -2 -3 26 103
use INVX1  INVX1_230
timestamp 1693479267
transform 1 0 1596 0 -1 2105
box -2 -3 18 103
use AOI21X1  AOI21X1_5
timestamp 1693479267
transform -1 0 1644 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_119
timestamp 1693479267
transform 1 0 1644 0 -1 2105
box -2 -3 26 103
use AOI22X1  AOI22X1_61
timestamp 1693479267
transform 1 0 1668 0 -1 2105
box -2 -3 42 103
use NAND2X1  NAND2X1_116
timestamp 1693479267
transform -1 0 1732 0 -1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_197
timestamp 1693479267
transform -1 0 1756 0 -1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_301
timestamp 1693479267
transform 1 0 1756 0 -1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_366
timestamp 1693479267
transform -1 0 1948 0 -1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_350
timestamp 1693479267
transform -1 0 2044 0 -1 2105
box -2 -3 98 103
use FILL  FILL_20_3_0
timestamp 1693479267
transform -1 0 2052 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_3_1
timestamp 1693479267
transform -1 0 2060 0 -1 2105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_364
timestamp 1693479267
transform -1 0 2156 0 -1 2105
box -2 -3 98 103
use INVX1  INVX1_690
timestamp 1693479267
transform 1 0 2156 0 -1 2105
box -2 -3 18 103
use XNOR2X1  XNOR2X1_55
timestamp 1693479267
transform 1 0 2172 0 -1 2105
box -2 -3 58 103
use NOR2X1  NOR2X1_438
timestamp 1693479267
transform -1 0 2252 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_929
timestamp 1693479267
transform -1 0 2284 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_709
timestamp 1693479267
transform -1 0 2300 0 -1 2105
box -2 -3 18 103
use NAND2X1  NAND2X1_955
timestamp 1693479267
transform 1 0 2300 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_930
timestamp 1693479267
transform -1 0 2356 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_689
timestamp 1693479267
transform -1 0 2372 0 -1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_437
timestamp 1693479267
transform -1 0 2396 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_237
timestamp 1693479267
transform -1 0 2428 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_335
timestamp 1693479267
transform -1 0 2460 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_961
timestamp 1693479267
transform 1 0 2460 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_908
timestamp 1693479267
transform -1 0 2516 0 -1 2105
box -2 -3 34 103
use AND2X2  AND2X2_95
timestamp 1693479267
transform 1 0 2516 0 -1 2105
box -2 -3 34 103
use FILL  FILL_20_4_0
timestamp 1693479267
transform 1 0 2548 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_4_1
timestamp 1693479267
transform 1 0 2556 0 -1 2105
box -2 -3 10 103
use AOI21X1  AOI21X1_247
timestamp 1693479267
transform 1 0 2564 0 -1 2105
box -2 -3 34 103
use OR2X2  OR2X2_62
timestamp 1693479267
transform 1 0 2596 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_956
timestamp 1693479267
transform 1 0 2628 0 -1 2105
box -2 -3 26 103
use AOI22X1  AOI22X1_132
timestamp 1693479267
transform 1 0 2652 0 -1 2105
box -2 -3 42 103
use INVX1  INVX1_306
timestamp 1693479267
transform 1 0 2692 0 -1 2105
box -2 -3 18 103
use NAND2X1  NAND2X1_957
timestamp 1693479267
transform -1 0 2732 0 -1 2105
box -2 -3 26 103
use OR2X2  OR2X2_63
timestamp 1693479267
transform -1 0 2764 0 -1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_246
timestamp 1693479267
transform 1 0 2764 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_958
timestamp 1693479267
transform 1 0 2796 0 -1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_457
timestamp 1693479267
transform -1 0 2844 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_926
timestamp 1693479267
transform 1 0 2844 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_458
timestamp 1693479267
transform 1 0 2876 0 -1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_991
timestamp 1693479267
transform 1 0 2900 0 -1 2105
box -2 -3 26 103
use INVX1  INVX1_707
timestamp 1693479267
transform -1 0 2940 0 -1 2105
box -2 -3 18 103
use NAND3X1  NAND3X1_339
timestamp 1693479267
transform 1 0 2940 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_684
timestamp 1693479267
transform 1 0 2972 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_907
timestamp 1693479267
transform 1 0 2988 0 -1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_235
timestamp 1693479267
transform 1 0 3020 0 -1 2105
box -2 -3 34 103
use FILL  FILL_20_5_0
timestamp 1693479267
transform -1 0 3060 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_5_1
timestamp 1693479267
transform -1 0 3068 0 -1 2105
box -2 -3 10 103
use INVX1  INVX1_700
timestamp 1693479267
transform -1 0 3084 0 -1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_450
timestamp 1693479267
transform -1 0 3108 0 -1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_938
timestamp 1693479267
transform 1 0 3108 0 -1 2105
box -2 -3 26 103
use INVX1  INVX1_671
timestamp 1693479267
transform 1 0 3132 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_904
timestamp 1693479267
transform 1 0 3148 0 -1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_242
timestamp 1693479267
transform 1 0 3180 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_425
timestamp 1693479267
transform 1 0 3212 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_252
timestamp 1693479267
transform -1 0 3268 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_308
timestamp 1693479267
transform -1 0 3284 0 -1 2105
box -2 -3 18 103
use NAND2X1  NAND2X1_989
timestamp 1693479267
transform -1 0 3308 0 -1 2105
box -2 -3 26 103
use AND2X2  AND2X2_83
timestamp 1693479267
transform -1 0 3340 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_340
timestamp 1693479267
transform 1 0 3340 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_202
timestamp 1693479267
transform -1 0 3396 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_287
timestamp 1693479267
transform -1 0 3428 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_310
timestamp 1693479267
transform -1 0 3444 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_286
timestamp 1693479267
transform -1 0 3476 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_309
timestamp 1693479267
transform -1 0 3492 0 -1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_460
timestamp 1693479267
transform 1 0 3492 0 -1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_462
timestamp 1693479267
transform -1 0 3540 0 -1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_990
timestamp 1693479267
transform -1 0 3564 0 -1 2105
box -2 -3 26 103
use FILL  FILL_20_6_0
timestamp 1693479267
transform -1 0 3572 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_6_1
timestamp 1693479267
transform -1 0 3580 0 -1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_282
timestamp 1693479267
transform -1 0 3612 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_309
timestamp 1693479267
transform -1 0 3636 0 -1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_88
timestamp 1693479267
transform -1 0 3660 0 -1 2105
box -2 -3 26 103
use INVX1  INVX1_312
timestamp 1693479267
transform -1 0 3676 0 -1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_89
timestamp 1693479267
transform -1 0 3700 0 -1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_90
timestamp 1693479267
transform -1 0 3724 0 -1 2105
box -2 -3 26 103
use INVX1  INVX1_433
timestamp 1693479267
transform 1 0 3724 0 -1 2105
box -2 -3 18 103
use AOI22X1  AOI22X1_109
timestamp 1693479267
transform 1 0 3740 0 -1 2105
box -2 -3 42 103
use OAI21X1  OAI21X1_781
timestamp 1693479267
transform 1 0 3780 0 -1 2105
box -2 -3 34 103
use INVX2  INVX2_24
timestamp 1693479267
transform 1 0 3812 0 -1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_162
timestamp 1693479267
transform 1 0 3828 0 -1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_91
timestamp 1693479267
transform -1 0 3876 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_721
timestamp 1693479267
transform -1 0 3908 0 -1 2105
box -2 -3 34 103
use AND2X2  AND2X2_64
timestamp 1693479267
transform -1 0 3940 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_710
timestamp 1693479267
transform 1 0 3940 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_431
timestamp 1693479267
transform 1 0 3972 0 -1 2105
box -2 -3 18 103
use AOI22X1  AOI22X1_108
timestamp 1693479267
transform 1 0 3988 0 -1 2105
box -2 -3 42 103
use OAI21X1  OAI21X1_771
timestamp 1693479267
transform -1 0 4060 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_430
timestamp 1693479267
transform -1 0 4076 0 -1 2105
box -2 -3 18 103
use FILL  FILL_20_7_0
timestamp 1693479267
transform -1 0 4084 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_7_1
timestamp 1693479267
transform -1 0 4092 0 -1 2105
box -2 -3 10 103
use OR2X2  OR2X2_15
timestamp 1693479267
transform -1 0 4124 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_582
timestamp 1693479267
transform 1 0 4124 0 -1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_87
timestamp 1693479267
transform -1 0 4172 0 -1 2105
box -2 -3 26 103
use NAND3X1  NAND3X1_95
timestamp 1693479267
transform -1 0 4204 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_137
timestamp 1693479267
transform -1 0 4228 0 -1 2105
box -2 -3 26 103
use INVX2  INVX2_23
timestamp 1693479267
transform -1 0 4244 0 -1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_86
timestamp 1693479267
transform 1 0 4244 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_751
timestamp 1693479267
transform 1 0 4268 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_426
timestamp 1693479267
transform 1 0 4300 0 -1 2105
box -2 -3 18 103
use AOI21X1  AOI21X1_203
timestamp 1693479267
transform 1 0 4316 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_427
timestamp 1693479267
transform -1 0 4364 0 -1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_364
timestamp 1693479267
transform 1 0 4364 0 -1 2105
box -2 -3 26 103
use INVX2  INVX2_71
timestamp 1693479267
transform 1 0 4388 0 -1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_83
timestamp 1693479267
transform -1 0 4428 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_207
timestamp 1693479267
transform -1 0 4460 0 -1 2105
box -2 -3 34 103
use INVX2  INVX2_21
timestamp 1693479267
transform 1 0 4460 0 -1 2105
box -2 -3 18 103
use INVX2  INVX2_20
timestamp 1693479267
transform 1 0 4476 0 -1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_84
timestamp 1693479267
transform 1 0 4492 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_742
timestamp 1693479267
transform -1 0 4548 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_722
timestamp 1693479267
transform -1 0 4580 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_356
timestamp 1693479267
transform -1 0 4604 0 -1 2105
box -2 -3 26 103
use BUFX2  BUFX2_26
timestamp 1693479267
transform -1 0 28 0 1 2105
box -2 -3 26 103
use BUFX2  BUFX2_30
timestamp 1693479267
transform -1 0 52 0 1 2105
box -2 -3 26 103
use BUFX2  BUFX2_39
timestamp 1693479267
transform -1 0 76 0 1 2105
box -2 -3 26 103
use BUFX2  BUFX2_67
timestamp 1693479267
transform -1 0 100 0 1 2105
box -2 -3 26 103
use INVX1  INVX1_168
timestamp 1693479267
transform -1 0 116 0 1 2105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_472
timestamp 1693479267
transform -1 0 212 0 1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_440
timestamp 1693479267
transform 1 0 212 0 1 2105
box -2 -3 98 103
use INVX1  INVX1_468
timestamp 1693479267
transform 1 0 308 0 1 2105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_183
timestamp 1693479267
transform -1 0 420 0 1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_815
timestamp 1693479267
transform 1 0 420 0 1 2105
box -2 -3 34 103
use BUFX2  BUFX2_98
timestamp 1693479267
transform -1 0 476 0 1 2105
box -2 -3 26 103
use FILL  FILL_21_0_0
timestamp 1693479267
transform -1 0 484 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_0_1
timestamp 1693479267
transform -1 0 492 0 1 2105
box -2 -3 10 103
use NOR3X1  NOR3X1_27
timestamp 1693479267
transform -1 0 556 0 1 2105
box -2 -3 66 103
use NAND2X1  NAND2X1_685
timestamp 1693479267
transform 1 0 556 0 1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_300
timestamp 1693479267
transform 1 0 580 0 1 2105
box -2 -3 98 103
use NOR2X1  NOR2X1_133
timestamp 1693479267
transform -1 0 700 0 1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_420
timestamp 1693479267
transform 1 0 700 0 1 2105
box -2 -3 98 103
use BUFX4  BUFX4_248
timestamp 1693479267
transform 1 0 796 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_639
timestamp 1693479267
transform -1 0 852 0 1 2105
box -2 -3 26 103
use BUFX2  BUFX2_84
timestamp 1693479267
transform -1 0 876 0 1 2105
box -2 -3 26 103
use NOR3X1  NOR3X1_7
timestamp 1693479267
transform -1 0 940 0 1 2105
box -2 -3 66 103
use INVX1  INVX1_144
timestamp 1693479267
transform -1 0 956 0 1 2105
box -2 -3 18 103
use NOR3X1  NOR3X1_6
timestamp 1693479267
transform -1 0 1020 0 1 2105
box -2 -3 66 103
use FILL  FILL_21_1_0
timestamp 1693479267
transform 1 0 1020 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_1_1
timestamp 1693479267
transform 1 0 1028 0 1 2105
box -2 -3 10 103
use XOR2X1  XOR2X1_7
timestamp 1693479267
transform 1 0 1036 0 1 2105
box -2 -3 58 103
use NAND2X1  NAND2X1_188
timestamp 1693479267
transform 1 0 1092 0 1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_58
timestamp 1693479267
transform 1 0 1116 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_186
timestamp 1693479267
transform -1 0 1164 0 1 2105
box -2 -3 26 103
use INVX1  INVX1_286
timestamp 1693479267
transform -1 0 1180 0 1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_56
timestamp 1693479267
transform -1 0 1204 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_185
timestamp 1693479267
transform -1 0 1228 0 1 2105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_45
timestamp 1693479267
transform -1 0 1284 0 1 2105
box -2 -3 58 103
use BUFX2  BUFX2_99
timestamp 1693479267
transform 1 0 1284 0 1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_282
timestamp 1693479267
transform 1 0 1308 0 1 2105
box -2 -3 98 103
use INVX1  INVX1_278
timestamp 1693479267
transform -1 0 1420 0 1 2105
box -2 -3 18 103
use NAND2X1  NAND2X1_182
timestamp 1693479267
transform -1 0 1444 0 1 2105
box -2 -3 26 103
use INVX1  INVX1_280
timestamp 1693479267
transform -1 0 1460 0 1 2105
box -2 -3 18 103
use NAND2X1  NAND2X1_181
timestamp 1693479267
transform -1 0 1484 0 1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_53
timestamp 1693479267
transform 1 0 1484 0 1 2105
box -2 -3 26 103
use FILL  FILL_21_2_0
timestamp 1693479267
transform -1 0 1516 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_2_1
timestamp 1693479267
transform -1 0 1524 0 1 2105
box -2 -3 10 103
use CLKBUF1  CLKBUF1_17
timestamp 1693479267
transform -1 0 1596 0 1 2105
box -2 -3 74 103
use CLKBUF1  CLKBUF1_58
timestamp 1693479267
transform 1 0 1596 0 1 2105
box -2 -3 74 103
use AOI22X1  AOI22X1_64
timestamp 1693479267
transform 1 0 1668 0 1 2105
box -2 -3 42 103
use AOI22X1  AOI22X1_62
timestamp 1693479267
transform 1 0 1708 0 1 2105
box -2 -3 42 103
use AOI22X1  AOI22X1_65
timestamp 1693479267
transform 1 0 1748 0 1 2105
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_347
timestamp 1693479267
transform -1 0 1884 0 1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_365
timestamp 1693479267
transform -1 0 1980 0 1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_346
timestamp 1693479267
transform -1 0 2076 0 1 2105
box -2 -3 98 103
use FILL  FILL_21_3_0
timestamp 1693479267
transform -1 0 2084 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_3_1
timestamp 1693479267
transform -1 0 2092 0 1 2105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_348
timestamp 1693479267
transform -1 0 2188 0 1 2105
box -2 -3 98 103
use INVX2  INVX2_82
timestamp 1693479267
transform 1 0 2188 0 1 2105
box -2 -3 18 103
use NAND2X1  NAND2X1_609
timestamp 1693479267
transform 1 0 2204 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_611
timestamp 1693479267
transform 1 0 2228 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_788
timestamp 1693479267
transform -1 0 2284 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_786
timestamp 1693479267
transform -1 0 2316 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_441
timestamp 1693479267
transform -1 0 2332 0 1 2105
box -2 -3 18 103
use INVX1  INVX1_439
timestamp 1693479267
transform -1 0 2348 0 1 2105
box -2 -3 18 103
use NAND2X1  NAND2X1_627
timestamp 1693479267
transform 1 0 2348 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_804
timestamp 1693479267
transform -1 0 2404 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_180
timestamp 1693479267
transform -1 0 2436 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_629
timestamp 1693479267
transform -1 0 2460 0 1 2105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_54
timestamp 1693479267
transform -1 0 2516 0 1 2105
box -2 -3 58 103
use FILL  FILL_21_4_0
timestamp 1693479267
transform -1 0 2524 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_4_1
timestamp 1693479267
transform -1 0 2532 0 1 2105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_344
timestamp 1693479267
transform -1 0 2628 0 1 2105
box -2 -3 98 103
use BUFX4  BUFX4_177
timestamp 1693479267
transform 1 0 2628 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_806
timestamp 1693479267
transform -1 0 2692 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_785
timestamp 1693479267
transform -1 0 2724 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_438
timestamp 1693479267
transform -1 0 2740 0 1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_931
timestamp 1693479267
transform -1 0 2772 0 1 2105
box -2 -3 34 103
use OR2X2  OR2X2_64
timestamp 1693479267
transform 1 0 2772 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_683
timestamp 1693479267
transform 1 0 2804 0 1 2105
box -2 -3 18 103
use NAND2X1  NAND2X1_959
timestamp 1693479267
transform 1 0 2820 0 1 2105
box -2 -3 26 103
use AOI22X1  AOI22X1_133
timestamp 1693479267
transform -1 0 2884 0 1 2105
box -2 -3 42 103
use INVX1  INVX1_685
timestamp 1693479267
transform -1 0 2900 0 1 2105
box -2 -3 18 103
use INVX1  INVX1_459
timestamp 1693479267
transform -1 0 2916 0 1 2105
box -2 -3 18 103
use INVX1  INVX1_457
timestamp 1693479267
transform -1 0 2932 0 1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_461
timestamp 1693479267
transform 1 0 2932 0 1 2105
box -2 -3 26 103
use OR2X2  OR2X2_68
timestamp 1693479267
transform 1 0 2956 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_939
timestamp 1693479267
transform 1 0 2988 0 1 2105
box -2 -3 26 103
use AOI22X1  AOI22X1_135
timestamp 1693479267
transform 1 0 3012 0 1 2105
box -2 -3 42 103
use FILL  FILL_21_5_0
timestamp 1693479267
transform 1 0 3052 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_5_1
timestamp 1693479267
transform 1 0 3060 0 1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_903
timestamp 1693479267
transform 1 0 3068 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_337
timestamp 1693479267
transform 1 0 3100 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_699
timestamp 1693479267
transform -1 0 3148 0 1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_447
timestamp 1693479267
transform -1 0 3172 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_918
timestamp 1693479267
transform 1 0 3172 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_712
timestamp 1693479267
transform 1 0 3204 0 1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_909
timestamp 1693479267
transform 1 0 3220 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_992
timestamp 1693479267
transform 1 0 3252 0 1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_255
timestamp 1693479267
transform -1 0 3308 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_713
timestamp 1693479267
transform -1 0 3324 0 1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_938
timestamp 1693479267
transform 1 0 3324 0 1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_455
timestamp 1693479267
transform -1 0 3380 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_993
timestamp 1693479267
transform -1 0 3404 0 1 2105
box -2 -3 26 103
use AOI22X1  AOI22X1_136
timestamp 1693479267
transform -1 0 3444 0 1 2105
box -2 -3 42 103
use NAND3X1  NAND3X1_343
timestamp 1693479267
transform -1 0 3476 0 1 2105
box -2 -3 34 103
use OR2X2  OR2X2_67
timestamp 1693479267
transform -1 0 3508 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_342
timestamp 1693479267
transform 1 0 3508 0 1 2105
box -2 -3 34 103
use OR2X2  OR2X2_66
timestamp 1693479267
transform -1 0 3572 0 1 2105
box -2 -3 34 103
use FILL  FILL_21_6_0
timestamp 1693479267
transform 1 0 3572 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_6_1
timestamp 1693479267
transform 1 0 3580 0 1 2105
box -2 -3 10 103
use NOR2X1  NOR2X1_456
timestamp 1693479267
transform 1 0 3588 0 1 2105
box -2 -3 26 103
use INVX1  INVX1_706
timestamp 1693479267
transform -1 0 3628 0 1 2105
box -2 -3 18 103
use INVX1  INVX1_304
timestamp 1693479267
transform -1 0 3644 0 1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_465
timestamp 1693479267
transform 1 0 3644 0 1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_181
timestamp 1693479267
transform 1 0 3668 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_432
timestamp 1693479267
transform 1 0 3700 0 1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_698
timestamp 1693479267
transform -1 0 3748 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_159
timestamp 1693479267
transform -1 0 3780 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_695
timestamp 1693479267
transform 1 0 3780 0 1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_177
timestamp 1693479267
transform 1 0 3812 0 1 2105
box -2 -3 34 103
use INVX2  INVX2_27
timestamp 1693479267
transform 1 0 3844 0 1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_374
timestamp 1693479267
transform -1 0 3884 0 1 2105
box -2 -3 26 103
use INVX1  INVX1_315
timestamp 1693479267
transform 1 0 3884 0 1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_92
timestamp 1693479267
transform -1 0 3924 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_337
timestamp 1693479267
transform 1 0 3924 0 1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_45
timestamp 1693479267
transform -1 0 3988 0 1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_93
timestamp 1693479267
transform 1 0 3988 0 1 2105
box -2 -3 26 103
use NAND3X1  NAND3X1_178
timestamp 1693479267
transform -1 0 4044 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_175
timestamp 1693479267
transform 1 0 4044 0 1 2105
box -2 -3 34 103
use FILL  FILL_21_7_0
timestamp 1693479267
transform -1 0 4084 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_7_1
timestamp 1693479267
transform -1 0 4092 0 1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_774
timestamp 1693479267
transform -1 0 4124 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_174
timestamp 1693479267
transform 1 0 4124 0 1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_138
timestamp 1693479267
transform -1 0 4180 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_316
timestamp 1693479267
transform -1 0 4204 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_333
timestamp 1693479267
transform 1 0 4204 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_336
timestamp 1693479267
transform -1 0 4268 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_428
timestamp 1693479267
transform 1 0 4268 0 1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_288
timestamp 1693479267
transform -1 0 4316 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_762
timestamp 1693479267
transform 1 0 4316 0 1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_211
timestamp 1693479267
transform -1 0 4380 0 1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_204
timestamp 1693479267
transform 1 0 4380 0 1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_85
timestamp 1693479267
transform 1 0 4412 0 1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_367
timestamp 1693479267
transform 1 0 4436 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_755
timestamp 1693479267
transform -1 0 4492 0 1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_200
timestamp 1693479267
transform 1 0 4492 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_424
timestamp 1693479267
transform 1 0 4524 0 1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_743
timestamp 1693479267
transform -1 0 4572 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_423
timestamp 1693479267
transform -1 0 4588 0 1 2105
box -2 -3 18 103
use FILL  FILL_22_1
timestamp 1693479267
transform 1 0 4588 0 1 2105
box -2 -3 10 103
use FILL  FILL_22_2
timestamp 1693479267
transform 1 0 4596 0 1 2105
box -2 -3 10 103
use BUFX2  BUFX2_28
timestamp 1693479267
transform -1 0 28 0 -1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_185
timestamp 1693479267
transform -1 0 124 0 -1 2305
box -2 -3 98 103
use INVX1  INVX1_187
timestamp 1693479267
transform 1 0 124 0 -1 2305
box -2 -3 18 103
use NOR3X1  NOR3X1_46
timestamp 1693479267
transform -1 0 204 0 -1 2305
box -2 -3 66 103
use DFFPOSX1  DFFPOSX1_439
timestamp 1693479267
transform 1 0 204 0 -1 2305
box -2 -3 98 103
use NAND2X1  NAND2X1_103
timestamp 1693479267
transform -1 0 324 0 -1 2305
box -2 -3 26 103
use AND2X2  AND2X2_2
timestamp 1693479267
transform -1 0 356 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_47
timestamp 1693479267
transform 1 0 356 0 -1 2305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_47
timestamp 1693479267
transform -1 0 460 0 -1 2305
box -2 -3 74 103
use BUFX4  BUFX4_140
timestamp 1693479267
transform -1 0 492 0 -1 2305
box -2 -3 34 103
use FILL  FILL_22_0_0
timestamp 1693479267
transform -1 0 500 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_0_1
timestamp 1693479267
transform -1 0 508 0 -1 2305
box -2 -3 10 103
use NOR3X1  NOR3X1_5
timestamp 1693479267
transform -1 0 572 0 -1 2305
box -2 -3 66 103
use INVX1  INVX1_142
timestamp 1693479267
transform -1 0 588 0 -1 2305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_296
timestamp 1693479267
transform 1 0 588 0 -1 2305
box -2 -3 98 103
use INVX1  INVX1_139
timestamp 1693479267
transform 1 0 684 0 -1 2305
box -2 -3 18 103
use NOR3X1  NOR3X1_2
timestamp 1693479267
transform -1 0 764 0 -1 2305
box -2 -3 66 103
use DFFPOSX1  DFFPOSX1_297
timestamp 1693479267
transform 1 0 764 0 -1 2305
box -2 -3 98 103
use NOR2X1  NOR2X1_134
timestamp 1693479267
transform 1 0 860 0 -1 2305
box -2 -3 26 103
use INVX1  INVX1_147
timestamp 1693479267
transform 1 0 884 0 -1 2305
box -2 -3 18 103
use INVX1  INVX1_146
timestamp 1693479267
transform 1 0 900 0 -1 2305
box -2 -3 18 103
use NOR3X1  NOR3X1_10
timestamp 1693479267
transform -1 0 980 0 -1 2305
box -2 -3 66 103
use INVX1  INVX1_143
timestamp 1693479267
transform 1 0 980 0 -1 2305
box -2 -3 18 103
use FILL  FILL_22_1_0
timestamp 1693479267
transform 1 0 996 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_1_1
timestamp 1693479267
transform 1 0 1004 0 -1 2305
box -2 -3 10 103
use NOR3X1  NOR3X1_9
timestamp 1693479267
transform 1 0 1012 0 -1 2305
box -2 -3 66 103
use INVX1  INVX1_283
timestamp 1693479267
transform -1 0 1092 0 -1 2305
box -2 -3 18 103
use INVX1  INVX1_288
timestamp 1693479267
transform -1 0 1108 0 -1 2305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_293
timestamp 1693479267
transform 1 0 1108 0 -1 2305
box -2 -3 98 103
use CLKBUF1  CLKBUF1_25
timestamp 1693479267
transform 1 0 1204 0 -1 2305
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_334
timestamp 1693479267
transform 1 0 1276 0 -1 2305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_294
timestamp 1693479267
transform 1 0 1372 0 -1 2305
box -2 -3 98 103
use INVX1  INVX1_279
timestamp 1693479267
transform 1 0 1468 0 -1 2305
box -2 -3 18 103
use CLKBUF1  CLKBUF1_4
timestamp 1693479267
transform 1 0 1484 0 -1 2305
box -2 -3 74 103
use FILL  FILL_22_2_0
timestamp 1693479267
transform -1 0 1564 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_2_1
timestamp 1693479267
transform -1 0 1572 0 -1 2305
box -2 -3 10 103
use INVX2  INVX2_5
timestamp 1693479267
transform -1 0 1588 0 -1 2305
box -2 -3 18 103
use CLKBUF1  CLKBUF1_2
timestamp 1693479267
transform 1 0 1588 0 -1 2305
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_159
timestamp 1693479267
transform 1 0 1660 0 -1 2305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_129
timestamp 1693479267
transform 1 0 1756 0 -1 2305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_367
timestamp 1693479267
transform -1 0 1948 0 -1 2305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_231
timestamp 1693479267
transform -1 0 2044 0 -1 2305
box -2 -3 98 103
use FILL  FILL_22_3_0
timestamp 1693479267
transform 1 0 2044 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_3_1
timestamp 1693479267
transform 1 0 2052 0 -1 2305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_360
timestamp 1693479267
transform 1 0 2060 0 -1 2305
box -2 -3 98 103
use NAND2X1  NAND2X1_625
timestamp 1693479267
transform 1 0 2156 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_802
timestamp 1693479267
transform -1 0 2212 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_610
timestamp 1693479267
transform 1 0 2212 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_628
timestamp 1693479267
transform 1 0 2236 0 -1 2305
box -2 -3 26 103
use INVX1  INVX1_442
timestamp 1693479267
transform 1 0 2260 0 -1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_789
timestamp 1693479267
transform 1 0 2276 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_805
timestamp 1693479267
transform -1 0 2340 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_801
timestamp 1693479267
transform -1 0 2372 0 -1 2305
box -2 -3 34 103
use INVX1  INVX1_454
timestamp 1693479267
transform -1 0 2388 0 -1 2305
box -2 -3 18 103
use INVX1  INVX1_458
timestamp 1693479267
transform -1 0 2404 0 -1 2305
box -2 -3 18 103
use BUFX4  BUFX4_264
timestamp 1693479267
transform 1 0 2404 0 -1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_345
timestamp 1693479267
transform -1 0 2532 0 -1 2305
box -2 -3 98 103
use NOR2X1  NOR2X1_377
timestamp 1693479267
transform 1 0 2532 0 -1 2305
box -2 -3 26 103
use FILL  FILL_22_4_0
timestamp 1693479267
transform 1 0 2556 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_4_1
timestamp 1693479267
transform 1 0 2564 0 -1 2305
box -2 -3 10 103
use NOR2X1  NOR2X1_378
timestamp 1693479267
transform 1 0 2572 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_607
timestamp 1693479267
transform -1 0 2620 0 -1 2305
box -2 -3 26 103
use INVX1  INVX1_437
timestamp 1693479267
transform -1 0 2636 0 -1 2305
box -2 -3 18 103
use NOR2X1  NOR2X1_376
timestamp 1693479267
transform -1 0 2660 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_608
timestamp 1693479267
transform 1 0 2660 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_605
timestamp 1693479267
transform 1 0 2684 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_784
timestamp 1693479267
transform -1 0 2740 0 -1 2305
box -2 -3 34 103
use INVX1  INVX1_435
timestamp 1693479267
transform -1 0 2756 0 -1 2305
box -2 -3 18 103
use NAND2X1  NAND2X1_616
timestamp 1693479267
transform 1 0 2756 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_944
timestamp 1693479267
transform 1 0 2780 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_445
timestamp 1693479267
transform -1 0 2828 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_905
timestamp 1693479267
transform 1 0 2828 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_916
timestamp 1693479267
transform 1 0 2860 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_943
timestamp 1693479267
transform 1 0 2892 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_906
timestamp 1693479267
transform 1 0 2916 0 -1 2305
box -2 -3 34 103
use NOR3X1  NOR3X1_70
timestamp 1693479267
transform -1 0 3012 0 -1 2305
box -2 -3 66 103
use AND2X2  AND2X2_85
timestamp 1693479267
transform 1 0 3012 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_427
timestamp 1693479267
transform -1 0 3068 0 -1 2305
box -2 -3 26 103
use FILL  FILL_22_5_0
timestamp 1693479267
transform 1 0 3068 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_5_1
timestamp 1693479267
transform 1 0 3076 0 -1 2305
box -2 -3 10 103
use INVX1  INVX1_697
timestamp 1693479267
transform 1 0 3084 0 -1 2305
box -2 -3 18 103
use NAND2X1  NAND2X1_974
timestamp 1693479267
transform 1 0 3100 0 -1 2305
box -2 -3 26 103
use AOI22X1  AOI22X1_134
timestamp 1693479267
transform -1 0 3164 0 -1 2305
box -2 -3 42 103
use NAND2X1  NAND2X1_975
timestamp 1693479267
transform 1 0 3164 0 -1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_251
timestamp 1693479267
transform 1 0 3188 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_934
timestamp 1693479267
transform 1 0 3220 0 -1 2305
box -2 -3 34 103
use INVX1  INVX1_714
timestamp 1693479267
transform 1 0 3252 0 -1 2305
box -2 -3 18 103
use NAND2X1  NAND2X1_977
timestamp 1693479267
transform -1 0 3292 0 -1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_243
timestamp 1693479267
transform -1 0 3324 0 -1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_332
timestamp 1693479267
transform 1 0 3324 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_983
timestamp 1693479267
transform 1 0 3356 0 -1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_250
timestamp 1693479267
transform 1 0 3380 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_937
timestamp 1693479267
transform 1 0 3412 0 -1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_240
timestamp 1693479267
transform -1 0 3476 0 -1 2305
box -2 -3 34 103
use AND2X2  AND2X2_93
timestamp 1693479267
transform -1 0 3508 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_968
timestamp 1693479267
transform 1 0 3508 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_429
timestamp 1693479267
transform -1 0 3556 0 -1 2305
box -2 -3 26 103
use INVX1  INVX1_676
timestamp 1693479267
transform -1 0 3572 0 -1 2305
box -2 -3 18 103
use FILL  FILL_22_6_0
timestamp 1693479267
transform 1 0 3572 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_6_1
timestamp 1693479267
transform 1 0 3580 0 -1 2305
box -2 -3 10 103
use INVX1  INVX1_675
timestamp 1693479267
transform 1 0 3588 0 -1 2305
box -2 -3 18 103
use NAND2X1  NAND2X1_987
timestamp 1693479267
transform 1 0 3604 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_986
timestamp 1693479267
transform -1 0 3652 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_428
timestamp 1693479267
transform -1 0 3676 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_430
timestamp 1693479267
transform 1 0 3676 0 -1 2305
box -2 -3 26 103
use INVX1  INVX1_695
timestamp 1693479267
transform 1 0 3700 0 -1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_913
timestamp 1693479267
transform -1 0 3748 0 -1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_239
timestamp 1693479267
transform -1 0 3780 0 -1 2305
box -2 -3 34 103
use INVX1  INVX1_691
timestamp 1693479267
transform -1 0 3796 0 -1 2305
box -2 -3 18 103
use INVX1  INVX1_710
timestamp 1693479267
transform 1 0 3796 0 -1 2305
box -2 -3 18 103
use NOR2X1  NOR2X1_432
timestamp 1693479267
transform -1 0 3836 0 -1 2305
box -2 -3 26 103
use INVX1  INVX1_680
timestamp 1693479267
transform 1 0 3836 0 -1 2305
box -2 -3 18 103
use NAND2X1  NAND2X1_948
timestamp 1693479267
transform -1 0 3876 0 -1 2305
box -2 -3 26 103
use INVX1  INVX1_679
timestamp 1693479267
transform 1 0 3876 0 -1 2305
box -2 -3 18 103
use NOR2X1  NOR2X1_441
timestamp 1693479267
transform -1 0 3916 0 -1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_238
timestamp 1693479267
transform -1 0 3948 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_967
timestamp 1693479267
transform -1 0 3972 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_440
timestamp 1693479267
transform 1 0 3972 0 -1 2305
box -2 -3 26 103
use INVX1  INVX1_694
timestamp 1693479267
transform -1 0 4012 0 -1 2305
box -2 -3 18 103
use INVX2  INVX2_26
timestamp 1693479267
transform -1 0 4028 0 -1 2305
box -2 -3 18 103
use NAND3X1  NAND3X1_177
timestamp 1693479267
transform 1 0 4028 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_783
timestamp 1693479267
transform -1 0 4092 0 -1 2305
box -2 -3 34 103
use FILL  FILL_22_7_0
timestamp 1693479267
transform 1 0 4092 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_7_1
timestamp 1693479267
transform 1 0 4100 0 -1 2305
box -2 -3 10 103
use INVX1  INVX1_434
timestamp 1693479267
transform 1 0 4108 0 -1 2305
box -2 -3 18 103
use NAND3X1  NAND3X1_176
timestamp 1693479267
transform 1 0 4124 0 -1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_88
timestamp 1693479267
transform 1 0 4156 0 -1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_172
timestamp 1693479267
transform 1 0 4188 0 -1 2305
box -2 -3 34 103
use OR2X2  OR2X2_43
timestamp 1693479267
transform -1 0 4252 0 -1 2305
box -2 -3 34 103
use INVX1  INVX1_311
timestamp 1693479267
transform -1 0 4268 0 -1 2305
box -2 -3 18 103
use AOI21X1  AOI21X1_214
timestamp 1693479267
transform -1 0 4300 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_773
timestamp 1693479267
transform -1 0 4332 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_597
timestamp 1693479267
transform 1 0 4332 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_362
timestamp 1693479267
transform -1 0 4380 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_363
timestamp 1693479267
transform -1 0 4404 0 -1 2305
box -2 -3 26 103
use AND2X2  AND2X2_69
timestamp 1693479267
transform 1 0 4404 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_756
timestamp 1693479267
transform -1 0 4468 0 -1 2305
box -2 -3 34 103
use INVX2  INVX2_22
timestamp 1693479267
transform -1 0 4484 0 -1 2305
box -2 -3 18 103
use NAND3X1  NAND3X1_171
timestamp 1693479267
transform -1 0 4516 0 -1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_170
timestamp 1693479267
transform 1 0 4516 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_754
timestamp 1693479267
transform -1 0 4580 0 -1 2305
box -2 -3 34 103
use FILL  FILL_23_1
timestamp 1693479267
transform -1 0 4588 0 -1 2305
box -2 -3 10 103
use FILL  FILL_23_2
timestamp 1693479267
transform -1 0 4596 0 -1 2305
box -2 -3 10 103
use FILL  FILL_23_3
timestamp 1693479267
transform -1 0 4604 0 -1 2305
box -2 -3 10 103
use INVX1  INVX1_181
timestamp 1693479267
transform 1 0 4 0 1 2305
box -2 -3 18 103
use INVX1  INVX1_169
timestamp 1693479267
transform 1 0 20 0 1 2305
box -2 -3 18 103
use CLKBUF1  CLKBUF1_44
timestamp 1693479267
transform -1 0 108 0 1 2305
box -2 -3 74 103
use NOR3X1  NOR3X1_40
timestamp 1693479267
transform -1 0 172 0 1 2305
box -2 -3 66 103
use NOR3X1  NOR3X1_28
timestamp 1693479267
transform -1 0 236 0 1 2305
box -2 -3 66 103
use DFFPOSX1  DFFPOSX1_433
timestamp 1693479267
transform 1 0 236 0 1 2305
box -2 -3 98 103
use BUFX4  BUFX4_50
timestamp 1693479267
transform -1 0 364 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_421
timestamp 1693479267
transform 1 0 364 0 1 2305
box -2 -3 98 103
use BUFX4  BUFX4_246
timestamp 1693479267
transform 1 0 460 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_0_0
timestamp 1693479267
transform 1 0 492 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_0_1
timestamp 1693479267
transform 1 0 500 0 1 2305
box -2 -3 10 103
use BUFX2  BUFX2_85
timestamp 1693479267
transform 1 0 508 0 1 2305
box -2 -3 26 103
use INVX8  INVX8_14
timestamp 1693479267
transform 1 0 532 0 1 2305
box -2 -3 42 103
use INVX1  INVX1_131
timestamp 1693479267
transform 1 0 572 0 1 2305
box -2 -3 18 103
use NOR3X1  NOR3X1_1
timestamp 1693479267
transform 1 0 588 0 1 2305
box -2 -3 66 103
use BUFX2  BUFX2_92
timestamp 1693479267
transform 1 0 652 0 1 2305
box -2 -3 26 103
use BUFX2  BUFX2_96
timestamp 1693479267
transform 1 0 676 0 1 2305
box -2 -3 26 103
use BUFX2  BUFX2_93
timestamp 1693479267
transform -1 0 724 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_883
timestamp 1693479267
transform -1 0 756 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_654
timestamp 1693479267
transform -1 0 772 0 1 2305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_315
timestamp 1693479267
transform 1 0 772 0 1 2305
box -2 -3 98 103
use INVX1  INVX1_652
timestamp 1693479267
transform 1 0 868 0 1 2305
box -2 -3 18 103
use INVX1  INVX1_655
timestamp 1693479267
transform 1 0 884 0 1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_884
timestamp 1693479267
transform 1 0 900 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_649
timestamp 1693479267
transform 1 0 932 0 1 2305
box -2 -3 18 103
use NOR2X1  NOR2X1_417
timestamp 1693479267
transform 1 0 948 0 1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_414
timestamp 1693479267
transform 1 0 972 0 1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_415
timestamp 1693479267
transform 1 0 996 0 1 2305
box -2 -3 26 103
use FILL  FILL_23_1_0
timestamp 1693479267
transform 1 0 1020 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_1_1
timestamp 1693479267
transform 1 0 1028 0 1 2305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_310
timestamp 1693479267
transform 1 0 1036 0 1 2305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_309
timestamp 1693479267
transform 1 0 1132 0 1 2305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_312
timestamp 1693479267
transform 1 0 1228 0 1 2305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_316
timestamp 1693479267
transform 1 0 1324 0 1 2305
box -2 -3 98 103
use BUFX4  BUFX4_6
timestamp 1693479267
transform 1 0 1420 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_150
timestamp 1693479267
transform 1 0 1452 0 1 2305
box -2 -3 98 103
use FILL  FILL_23_2_0
timestamp 1693479267
transform 1 0 1548 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_2_1
timestamp 1693479267
transform 1 0 1556 0 1 2305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_130
timestamp 1693479267
transform 1 0 1564 0 1 2305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_18
timestamp 1693479267
transform -1 0 1756 0 1 2305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_17
timestamp 1693479267
transform -1 0 1852 0 1 2305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_361
timestamp 1693479267
transform -1 0 1948 0 1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_23
timestamp 1693479267
transform -1 0 1980 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_23
timestamp 1693479267
transform -1 0 1996 0 1 2305
box -2 -3 18 103
use FILL  FILL_23_3_0
timestamp 1693479267
transform -1 0 2004 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_3_1
timestamp 1693479267
transform -1 0 2012 0 1 2305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_368
timestamp 1693479267
transform -1 0 2108 0 1 2305
box -2 -3 98 103
use OAI21X1  OAI21X1_25
timestamp 1693479267
transform -1 0 2140 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_25
timestamp 1693479267
transform -1 0 2156 0 1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_3
timestamp 1693479267
transform -1 0 2188 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_3
timestamp 1693479267
transform -1 0 2204 0 1 2305
box -2 -3 18 103
use INVX1  INVX1_5
timestamp 1693479267
transform 1 0 2204 0 1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_5
timestamp 1693479267
transform 1 0 2220 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_787
timestamp 1693479267
transform -1 0 2284 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_440
timestamp 1693479267
transform -1 0 2300 0 1 2305
box -2 -3 18 103
use NAND2X1  NAND2X1_612
timestamp 1693479267
transform -1 0 2324 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_624
timestamp 1693479267
transform -1 0 2348 0 1 2305
box -2 -3 26 103
use INVX1  INVX1_455
timestamp 1693479267
transform -1 0 2364 0 1 2305
box -2 -3 18 103
use BUFX4  BUFX4_265
timestamp 1693479267
transform -1 0 2396 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_613
timestamp 1693479267
transform 1 0 2396 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_790
timestamp 1693479267
transform -1 0 2452 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_443
timestamp 1693479267
transform -1 0 2468 0 1 2305
box -2 -3 18 103
use BUFX4  BUFX4_181
timestamp 1693479267
transform 1 0 2468 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_4_0
timestamp 1693479267
transform -1 0 2508 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_4_1
timestamp 1693479267
transform -1 0 2516 0 1 2305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_356
timestamp 1693479267
transform -1 0 2612 0 1 2305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_357
timestamp 1693479267
transform -1 0 2708 0 1 2305
box -2 -3 98 103
use NAND2X1  NAND2X1_606
timestamp 1693479267
transform -1 0 2732 0 1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_375
timestamp 1693479267
transform 1 0 2732 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_638
timestamp 1693479267
transform 1 0 2756 0 1 2305
box -2 -3 26 103
use INVX1  INVX1_436
timestamp 1693479267
transform 1 0 2780 0 1 2305
box -2 -3 18 103
use INVX2  INVX2_83
timestamp 1693479267
transform 1 0 2796 0 1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_793
timestamp 1693479267
transform -1 0 2844 0 1 2305
box -2 -3 34 103
use BUFX4  BUFX4_268
timestamp 1693479267
transform -1 0 2876 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_614
timestamp 1693479267
transform 1 0 2876 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_619
timestamp 1693479267
transform -1 0 2924 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_791
timestamp 1693479267
transform -1 0 2956 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_796
timestamp 1693479267
transform -1 0 2988 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_426
timestamp 1693479267
transform -1 0 3012 0 1 2305
box -2 -3 26 103
use OAI22X1  OAI22X1_50
timestamp 1693479267
transform 1 0 3012 0 1 2305
box -2 -3 42 103
use FILL  FILL_23_5_0
timestamp 1693479267
transform -1 0 3060 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_5_1
timestamp 1693479267
transform -1 0 3068 0 1 2305
box -2 -3 10 103
use AND2X2  AND2X2_84
timestamp 1693479267
transform -1 0 3100 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_698
timestamp 1693479267
transform 1 0 3100 0 1 2305
box -2 -3 18 103
use NAND2X1  NAND2X1_972
timestamp 1693479267
transform 1 0 3116 0 1 2305
box -2 -3 26 103
use INVX1  INVX1_75
timestamp 1693479267
transform -1 0 3156 0 1 2305
box -2 -3 18 103
use NOR2X1  NOR2X1_446
timestamp 1693479267
transform -1 0 3180 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_917
timestamp 1693479267
transform -1 0 3212 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_973
timestamp 1693479267
transform -1 0 3236 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_933
timestamp 1693479267
transform -1 0 3268 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_696
timestamp 1693479267
transform -1 0 3284 0 1 2305
box -2 -3 18 103
use NAND2X1  NAND2X1_976
timestamp 1693479267
transform 1 0 3284 0 1 2305
box -2 -3 26 103
use AND2X2  AND2X2_91
timestamp 1693479267
transform 1 0 3308 0 1 2305
box -2 -3 34 103
use INVX2  INVX2_86
timestamp 1693479267
transform -1 0 3356 0 1 2305
box -2 -3 18 103
use INVX1  INVX1_449
timestamp 1693479267
transform -1 0 3372 0 1 2305
box -2 -3 18 103
use AOI21X1  AOI21X1_254
timestamp 1693479267
transform 1 0 3372 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_941
timestamp 1693479267
transform -1 0 3436 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_245
timestamp 1693479267
transform -1 0 3468 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_338
timestamp 1693479267
transform 1 0 3468 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_925
timestamp 1693479267
transform 1 0 3500 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_924
timestamp 1693479267
transform 1 0 3532 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_6_0
timestamp 1693479267
transform 1 0 3564 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_6_1
timestamp 1693479267
transform 1 0 3572 0 1 2305
box -2 -3 10 103
use INVX1  INVX1_677
timestamp 1693479267
transform 1 0 3580 0 1 2305
box -2 -3 18 103
use NAND2X1  NAND2X1_945
timestamp 1693479267
transform -1 0 3620 0 1 2305
box -2 -3 26 103
use INVX1  INVX1_678
timestamp 1693479267
transform 1 0 3620 0 1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_912
timestamp 1693479267
transform -1 0 3668 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_946
timestamp 1693479267
transform -1 0 3692 0 1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_459
timestamp 1693479267
transform 1 0 3692 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_988
timestamp 1693479267
transform -1 0 3740 0 1 2305
box -2 -3 26 103
use AND2X2  AND2X2_86
timestamp 1693479267
transform 1 0 3740 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_966
timestamp 1693479267
transform -1 0 3796 0 1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_249
timestamp 1693479267
transform -1 0 3828 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_932
timestamp 1693479267
transform -1 0 3860 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_333
timestamp 1693479267
transform 1 0 3860 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_947
timestamp 1693479267
transform 1 0 3892 0 1 2305
box -2 -3 26 103
use AOI22X1  AOI22X1_129
timestamp 1693479267
transform -1 0 3956 0 1 2305
box -2 -3 42 103
use NAND2X1  NAND2X1_949
timestamp 1693479267
transform -1 0 3980 0 1 2305
box -2 -3 26 103
use OR2X2  OR2X2_57
timestamp 1693479267
transform -1 0 4012 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_248
timestamp 1693479267
transform -1 0 4044 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_963
timestamp 1693479267
transform 1 0 4044 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_965
timestamp 1693479267
transform 1 0 4068 0 1 2305
box -2 -3 26 103
use FILL  FILL_23_7_0
timestamp 1693479267
transform -1 0 4100 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_7_1
timestamp 1693479267
transform -1 0 4108 0 1 2305
box -2 -3 10 103
use AND2X2  AND2X2_88
timestamp 1693479267
transform -1 0 4140 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_985
timestamp 1693479267
transform -1 0 4164 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_603
timestamp 1693479267
transform 1 0 4164 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_602
timestamp 1693479267
transform 1 0 4188 0 1 2305
box -2 -3 26 103
use NAND3X1  NAND3X1_173
timestamp 1693479267
transform -1 0 4244 0 1 2305
box -2 -3 34 103
use INVX2  INVX2_28
timestamp 1693479267
transform 1 0 4244 0 1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_764
timestamp 1693479267
transform 1 0 4260 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_370
timestamp 1693479267
transform -1 0 4316 0 1 2305
box -2 -3 26 103
use NAND3X1  NAND3X1_169
timestamp 1693479267
transform -1 0 4348 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_752
timestamp 1693479267
transform 1 0 4348 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_208
timestamp 1693479267
transform -1 0 4412 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_964
timestamp 1693479267
transform 1 0 4412 0 1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_366
timestamp 1693479267
transform -1 0 4460 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_600
timestamp 1693479267
transform -1 0 4484 0 1 2305
box -2 -3 26 103
use INVX1  INVX1_429
timestamp 1693479267
transform -1 0 4500 0 1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_763
timestamp 1693479267
transform -1 0 4532 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_744
timestamp 1693479267
transform 1 0 4532 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_358
timestamp 1693479267
transform 1 0 4564 0 1 2305
box -2 -3 26 103
use FILL  FILL_24_1
timestamp 1693479267
transform 1 0 4588 0 1 2305
box -2 -3 10 103
use FILL  FILL_24_2
timestamp 1693479267
transform 1 0 4596 0 1 2305
box -2 -3 10 103
use INVX1  INVX1_185
timestamp 1693479267
transform 1 0 4 0 -1 2505
box -2 -3 18 103
use NOR3X1  NOR3X1_44
timestamp 1693479267
transform -1 0 84 0 -1 2505
box -2 -3 66 103
use DFFPOSX1  DFFPOSX1_437
timestamp 1693479267
transform 1 0 84 0 -1 2505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_438
timestamp 1693479267
transform 1 0 180 0 -1 2505
box -2 -3 98 103
use BUFX2  BUFX2_97
timestamp 1693479267
transform 1 0 276 0 -1 2505
box -2 -3 26 103
use NOR3X1  NOR3X1_3
timestamp 1693479267
transform -1 0 364 0 -1 2505
box -2 -3 66 103
use INVX1  INVX1_140
timestamp 1693479267
transform -1 0 380 0 -1 2505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_298
timestamp 1693479267
transform 1 0 380 0 -1 2505
box -2 -3 98 103
use INVX1  INVX1_148
timestamp 1693479267
transform 1 0 476 0 -1 2505
box -2 -3 18 103
use FILL  FILL_24_0_0
timestamp 1693479267
transform 1 0 492 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_0_1
timestamp 1693479267
transform 1 0 500 0 -1 2505
box -2 -3 10 103
use NOR3X1  NOR3X1_11
timestamp 1693479267
transform 1 0 508 0 -1 2505
box -2 -3 66 103
use OR2X2  OR2X2_17
timestamp 1693479267
transform 1 0 572 0 -1 2505
box -2 -3 34 103
use NOR3X1  NOR3X1_4
timestamp 1693479267
transform 1 0 604 0 -1 2505
box -2 -3 66 103
use DFFPOSX1  DFFPOSX1_324
timestamp 1693479267
transform 1 0 668 0 -1 2505
box -2 -3 98 103
use CLKBUF1  CLKBUF1_56
timestamp 1693479267
transform -1 0 836 0 -1 2505
box -2 -3 74 103
use AOI22X1  AOI22X1_125
timestamp 1693479267
transform 1 0 836 0 -1 2505
box -2 -3 42 103
use AOI22X1  AOI22X1_120
timestamp 1693479267
transform 1 0 876 0 -1 2505
box -2 -3 42 103
use OAI21X1  OAI21X1_896
timestamp 1693479267
transform -1 0 948 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_901
timestamp 1693479267
transform 1 0 948 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_650
timestamp 1693479267
transform 1 0 980 0 -1 2505
box -2 -3 18 103
use INVX2  INVX2_14
timestamp 1693479267
transform -1 0 1012 0 -1 2505
box -2 -3 18 103
use FILL  FILL_24_1_0
timestamp 1693479267
transform -1 0 1020 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_1_1
timestamp 1693479267
transform -1 0 1028 0 -1 2505
box -2 -3 10 103
use INVX1  INVX1_271
timestamp 1693479267
transform -1 0 1044 0 -1 2505
box -2 -3 18 103
use BUFX4  BUFX4_260
timestamp 1693479267
transform 1 0 1044 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_653
timestamp 1693479267
transform 1 0 1076 0 -1 2505
box -2 -3 18 103
use INVX1  INVX1_648
timestamp 1693479267
transform 1 0 1092 0 -1 2505
box -2 -3 18 103
use NOR2X1  NOR2X1_418
timestamp 1693479267
transform 1 0 1108 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_413
timestamp 1693479267
transform -1 0 1156 0 -1 2505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_313
timestamp 1693479267
transform 1 0 1156 0 -1 2505
box -2 -3 98 103
use INVX1  INVX1_285
timestamp 1693479267
transform -1 0 1268 0 -1 2505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_328
timestamp 1693479267
transform 1 0 1268 0 -1 2505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_333
timestamp 1693479267
transform 1 0 1364 0 -1 2505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_308
timestamp 1693479267
transform 1 0 1460 0 -1 2505
box -2 -3 98 103
use FILL  FILL_24_2_0
timestamp 1693479267
transform 1 0 1556 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_2_1
timestamp 1693479267
transform 1 0 1564 0 -1 2505
box -2 -3 10 103
use CLKBUF1  CLKBUF1_12
timestamp 1693479267
transform 1 0 1572 0 -1 2505
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_38
timestamp 1693479267
transform -1 0 1740 0 -1 2505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_132
timestamp 1693479267
transform -1 0 1836 0 -1 2505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_133
timestamp 1693479267
transform -1 0 1932 0 -1 2505
box -2 -3 98 103
use OAI21X1  OAI21X1_4
timestamp 1693479267
transform -1 0 1964 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_4
timestamp 1693479267
transform -1 0 1980 0 -1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_18
timestamp 1693479267
transform -1 0 2012 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_18
timestamp 1693479267
transform -1 0 2028 0 -1 2505
box -2 -3 18 103
use FILL  FILL_24_3_0
timestamp 1693479267
transform -1 0 2036 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_3_1
timestamp 1693479267
transform -1 0 2044 0 -1 2505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_225
timestamp 1693479267
transform -1 0 2140 0 -1 2505
box -2 -3 98 103
use OAI21X1  OAI21X1_21
timestamp 1693479267
transform 1 0 2140 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_21
timestamp 1693479267
transform -1 0 2188 0 -1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_24
timestamp 1693479267
transform -1 0 2220 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_24
timestamp 1693479267
transform -1 0 2236 0 -1 2505
box -2 -3 18 103
use BUFX4  BUFX4_21
timestamp 1693479267
transform -1 0 2268 0 -1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_244
timestamp 1693479267
transform 1 0 2268 0 -1 2505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_363
timestamp 1693479267
transform 1 0 2364 0 -1 2505
box -2 -3 98 103
use NAND2X1  NAND2X1_626
timestamp 1693479267
transform 1 0 2460 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_803
timestamp 1693479267
transform -1 0 2516 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_623
timestamp 1693479267
transform 1 0 2516 0 -1 2505
box -2 -3 26 103
use FILL  FILL_24_4_0
timestamp 1693479267
transform -1 0 2548 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_4_1
timestamp 1693479267
transform -1 0 2556 0 -1 2505
box -2 -3 10 103
use OAI21X1  OAI21X1_800
timestamp 1693479267
transform -1 0 2588 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_622
timestamp 1693479267
transform 1 0 2588 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_799
timestamp 1693479267
transform -1 0 2644 0 -1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_359
timestamp 1693479267
transform 1 0 2644 0 -1 2505
box -2 -3 98 103
use NAND2X1  NAND2X1_620
timestamp 1693479267
transform -1 0 2764 0 -1 2505
box -2 -3 26 103
use INVX1  INVX1_453
timestamp 1693479267
transform -1 0 2780 0 -1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_8
timestamp 1693479267
transform -1 0 2812 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_8
timestamp 1693479267
transform -1 0 2828 0 -1 2505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_351
timestamp 1693479267
transform 1 0 2828 0 -1 2505
box -2 -3 98 103
use INVX1  INVX1_10
timestamp 1693479267
transform -1 0 2940 0 -1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_2
timestamp 1693479267
transform -1 0 2972 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_456
timestamp 1693479267
transform -1 0 2988 0 -1 2505
box -2 -3 18 103
use INVX1  INVX1_2
timestamp 1693479267
transform -1 0 3004 0 -1 2505
box -2 -3 18 103
use NAND2X1  NAND2X1_80
timestamp 1693479267
transform 1 0 3004 0 -1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_79
timestamp 1693479267
transform -1 0 3052 0 -1 2505
box -2 -3 26 103
use FILL  FILL_24_5_0
timestamp 1693479267
transform -1 0 3060 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_5_1
timestamp 1693479267
transform -1 0 3068 0 -1 2505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_375
timestamp 1693479267
transform -1 0 3164 0 -1 2505
box -2 -3 98 103
use NAND2X1  NAND2X1_76
timestamp 1693479267
transform -1 0 3188 0 -1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_77
timestamp 1693479267
transform 1 0 3188 0 -1 2505
box -2 -3 26 103
use INVX1  INVX1_452
timestamp 1693479267
transform -1 0 3228 0 -1 2505
box -2 -3 18 103
use INVX1  INVX1_674
timestamp 1693479267
transform -1 0 3244 0 -1 2505
box -2 -3 18 103
use INVX1  INVX1_444
timestamp 1693479267
transform -1 0 3260 0 -1 2505
box -2 -3 18 103
use BUFX4  BUFX4_267
timestamp 1693479267
transform 1 0 3260 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_637
timestamp 1693479267
transform 1 0 3292 0 -1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_618
timestamp 1693479267
transform 1 0 3316 0 -1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_615
timestamp 1693479267
transform 1 0 3340 0 -1 2505
box -2 -3 26 103
use BUFX4  BUFX4_266
timestamp 1693479267
transform 1 0 3364 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_446
timestamp 1693479267
transform -1 0 3412 0 -1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_795
timestamp 1693479267
transform -1 0 3444 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_792
timestamp 1693479267
transform -1 0 3476 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_448
timestamp 1693479267
transform -1 0 3492 0 -1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_814
timestamp 1693479267
transform -1 0 3524 0 -1 2505
box -2 -3 34 103
use BUFX4  BUFX4_179
timestamp 1693479267
transform 1 0 3524 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_467
timestamp 1693479267
transform -1 0 3572 0 -1 2505
box -2 -3 18 103
use FILL  FILL_24_6_0
timestamp 1693479267
transform 1 0 3572 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_6_1
timestamp 1693479267
transform 1 0 3580 0 -1 2505
box -2 -3 10 103
use NAND2X1  NAND2X1_929
timestamp 1693479267
transform 1 0 3588 0 -1 2505
box -2 -3 26 103
use INVX1  INVX1_666
timestamp 1693479267
transform -1 0 3628 0 -1 2505
box -2 -3 18 103
use INVX1  INVX1_665
timestamp 1693479267
transform 1 0 3628 0 -1 2505
box -2 -3 18 103
use NAND2X1  NAND2X1_969
timestamp 1693479267
transform 1 0 3644 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_421
timestamp 1693479267
transform -1 0 3692 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_922
timestamp 1693479267
transform 1 0 3692 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_970
timestamp 1693479267
transform 1 0 3724 0 -1 2505
box -2 -3 26 103
use INVX1  INVX1_664
timestamp 1693479267
transform 1 0 3748 0 -1 2505
box -2 -3 18 103
use NAND2X1  NAND2X1_928
timestamp 1693479267
transform -1 0 3788 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_422
timestamp 1693479267
transform -1 0 3812 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_420
timestamp 1693479267
transform -1 0 3836 0 -1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_981
timestamp 1693479267
transform 1 0 3836 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_923
timestamp 1693479267
transform 1 0 3860 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_705
timestamp 1693479267
transform -1 0 3908 0 -1 2505
box -2 -3 18 103
use NAND3X1  NAND3X1_341
timestamp 1693479267
transform 1 0 3908 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_454
timestamp 1693479267
transform 1 0 3940 0 -1 2505
box -2 -3 26 103
use NAND3X1  NAND3X1_330
timestamp 1693479267
transform 1 0 3964 0 -1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_336
timestamp 1693479267
transform 1 0 3996 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_936
timestamp 1693479267
transform -1 0 4060 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_452
timestamp 1693479267
transform -1 0 4084 0 -1 2505
box -2 -3 26 103
use FILL  FILL_24_7_0
timestamp 1693479267
transform -1 0 4092 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_7_1
timestamp 1693479267
transform -1 0 4100 0 -1 2505
box -2 -3 10 103
use INVX1  INVX1_445
timestamp 1693479267
transform -1 0 4116 0 -1 2505
box -2 -3 18 103
use NOR2X1  NOR2X1_424
timestamp 1693479267
transform -1 0 4140 0 -1 2505
box -2 -3 26 103
use AND2X2  AND2X2_96
timestamp 1693479267
transform 1 0 4140 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_463
timestamp 1693479267
transform 1 0 4172 0 -1 2505
box -2 -3 26 103
use OAI22X1  OAI22X1_52
timestamp 1693479267
transform 1 0 4196 0 -1 2505
box -2 -3 42 103
use NOR2X1  NOR2X1_464
timestamp 1693479267
transform -1 0 4260 0 -1 2505
box -2 -3 26 103
use NOR3X1  NOR3X1_72
timestamp 1693479267
transform 1 0 4260 0 -1 2505
box -2 -3 66 103
use OAI21X1  OAI21X1_939
timestamp 1693479267
transform 1 0 4324 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_940
timestamp 1693479267
transform 1 0 4356 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_953
timestamp 1693479267
transform 1 0 4388 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_910
timestamp 1693479267
transform -1 0 4444 0 -1 2505
box -2 -3 34 103
use AND2X2  AND2X2_87
timestamp 1693479267
transform 1 0 4444 0 -1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_334
timestamp 1693479267
transform 1 0 4476 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_693
timestamp 1693479267
transform -1 0 4524 0 -1 2505
box -2 -3 18 103
use NOR2X1  NOR2X1_439
timestamp 1693479267
transform -1 0 4548 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_911
timestamp 1693479267
transform -1 0 4580 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_692
timestamp 1693479267
transform 1 0 4580 0 -1 2505
box -2 -3 18 103
use FILL  FILL_25_1
timestamp 1693479267
transform -1 0 4604 0 -1 2505
box -2 -3 10 103
use INVX1  INVX1_170
timestamp 1693479267
transform 1 0 4 0 1 2505
box -2 -3 18 103
use INVX1  INVX1_186
timestamp 1693479267
transform 1 0 20 0 1 2505
box -2 -3 18 103
use NOR3X1  NOR3X1_29
timestamp 1693479267
transform -1 0 100 0 1 2505
box -2 -3 66 103
use NOR3X1  NOR3X1_45
timestamp 1693479267
transform -1 0 164 0 1 2505
box -2 -3 66 103
use DFFPOSX1  DFFPOSX1_422
timestamp 1693479267
transform 1 0 164 0 1 2505
box -2 -3 98 103
use BUFX4  BUFX4_249
timestamp 1693479267
transform -1 0 292 0 1 2505
box -2 -3 34 103
use BUFX2  BUFX2_86
timestamp 1693479267
transform 1 0 292 0 1 2505
box -2 -3 26 103
use CLKBUF1  CLKBUF1_13
timestamp 1693479267
transform 1 0 316 0 1 2505
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_295
timestamp 1693479267
transform 1 0 388 0 1 2505
box -2 -3 98 103
use INVX1  INVX1_656
timestamp 1693479267
transform 1 0 484 0 1 2505
box -2 -3 18 103
use FILL  FILL_25_0_0
timestamp 1693479267
transform -1 0 508 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_0_1
timestamp 1693479267
transform -1 0 516 0 1 2505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_299
timestamp 1693479267
transform -1 0 612 0 1 2505
box -2 -3 98 103
use INVX1  INVX1_141
timestamp 1693479267
transform 1 0 612 0 1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_885
timestamp 1693479267
transform 1 0 628 0 1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_317
timestamp 1693479267
transform 1 0 660 0 1 2505
box -2 -3 98 103
use BUFX4  BUFX4_263
timestamp 1693479267
transform 1 0 756 0 1 2505
box -2 -3 34 103
use AOI22X1  AOI22X1_124
timestamp 1693479267
transform 1 0 788 0 1 2505
box -2 -3 42 103
use OAI21X1  OAI21X1_900
timestamp 1693479267
transform -1 0 860 0 1 2505
box -2 -3 34 103
use AOI22X1  AOI22X1_122
timestamp 1693479267
transform 1 0 860 0 1 2505
box -2 -3 42 103
use OAI21X1  OAI21X1_898
timestamp 1693479267
transform -1 0 932 0 1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_332
timestamp 1693479267
transform 1 0 932 0 1 2505
box -2 -3 98 103
use FILL  FILL_25_1_0
timestamp 1693479267
transform 1 0 1028 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_1_1
timestamp 1693479267
transform 1 0 1036 0 1 2505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_330
timestamp 1693479267
transform 1 0 1044 0 1 2505
box -2 -3 98 103
use CLKBUF1  CLKBUF1_1
timestamp 1693479267
transform -1 0 1212 0 1 2505
box -2 -3 74 103
use CLKBUF1  CLKBUF1_32
timestamp 1693479267
transform -1 0 1284 0 1 2505
box -2 -3 74 103
use CLKBUF1  CLKBUF1_18
timestamp 1693479267
transform 1 0 1284 0 1 2505
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_127
timestamp 1693479267
transform 1 0 1356 0 1 2505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_20
timestamp 1693479267
transform -1 0 1548 0 1 2505
box -2 -3 98 103
use FILL  FILL_25_2_0
timestamp 1693479267
transform -1 0 1556 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_2_1
timestamp 1693479267
transform -1 0 1564 0 1 2505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_21
timestamp 1693479267
transform -1 0 1660 0 1 2505
box -2 -3 98 103
use BUFX4  BUFX4_7
timestamp 1693479267
transform 1 0 1660 0 1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_87
timestamp 1693479267
transform 1 0 1692 0 1 2505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_229
timestamp 1693479267
transform -1 0 1884 0 1 2505
box -2 -3 98 103
use NAND2X1  NAND2X1_23
timestamp 1693479267
transform 1 0 1884 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_4
timestamp 1693479267
transform 1 0 1908 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_22
timestamp 1693479267
transform 1 0 1932 0 1 2505
box -2 -3 34 103
use INVX1  INVX1_22
timestamp 1693479267
transform -1 0 1980 0 1 2505
box -2 -3 18 103
use NAND2X1  NAND2X1_18
timestamp 1693479267
transform 1 0 1980 0 1 2505
box -2 -3 26 103
use FILL  FILL_25_3_0
timestamp 1693479267
transform 1 0 2004 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_3_1
timestamp 1693479267
transform 1 0 2012 0 1 2505
box -2 -3 10 103
use CLKBUF1  CLKBUF1_53
timestamp 1693479267
transform 1 0 2020 0 1 2505
box -2 -3 74 103
use NAND2X1  NAND2X1_25
timestamp 1693479267
transform 1 0 2092 0 1 2505
box -2 -3 26 103
use BUFX4  BUFX4_18
timestamp 1693479267
transform -1 0 2148 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_21
timestamp 1693479267
transform 1 0 2148 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_24
timestamp 1693479267
transform 1 0 2172 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_70
timestamp 1693479267
transform 1 0 2196 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_68
timestamp 1693479267
transform -1 0 2252 0 1 2505
box -2 -3 34 103
use INVX1  INVX1_69
timestamp 1693479267
transform -1 0 2268 0 1 2505
box -2 -3 18 103
use NAND2X1  NAND2X1_5
timestamp 1693479267
transform 1 0 2268 0 1 2505
box -2 -3 26 103
use INVX1  INVX1_88
timestamp 1693479267
transform 1 0 2292 0 1 2505
box -2 -3 18 103
use INVX1  INVX1_73
timestamp 1693479267
transform 1 0 2308 0 1 2505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_358
timestamp 1693479267
transform -1 0 2420 0 1 2505
box -2 -3 98 103
use NAND2X1  NAND2X1_74
timestamp 1693479267
transform 1 0 2420 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_72
timestamp 1693479267
transform 1 0 2444 0 1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_352
timestamp 1693479267
transform -1 0 2572 0 1 2505
box -2 -3 98 103
use FILL  FILL_25_4_0
timestamp 1693479267
transform -1 0 2580 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_4_1
timestamp 1693479267
transform -1 0 2588 0 1 2505
box -2 -3 10 103
use OAI21X1  OAI21X1_13
timestamp 1693479267
transform -1 0 2620 0 1 2505
box -2 -3 34 103
use INVX1  INVX1_13
timestamp 1693479267
transform -1 0 2636 0 1 2505
box -2 -3 18 103
use INVX1  INVX1_16
timestamp 1693479267
transform 1 0 2636 0 1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_16
timestamp 1693479267
transform 1 0 2652 0 1 2505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_48
timestamp 1693479267
transform 1 0 2684 0 1 2505
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_353
timestamp 1693479267
transform -1 0 2852 0 1 2505
box -2 -3 98 103
use OAI21X1  OAI21X1_10
timestamp 1693479267
transform -1 0 2884 0 1 2505
box -2 -3 34 103
use INVX1  INVX1_1
timestamp 1693479267
transform 1 0 2884 0 1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_1
timestamp 1693479267
transform 1 0 2900 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_2
timestamp 1693479267
transform 1 0 2932 0 1 2505
box -2 -3 26 103
use INVX1  INVX1_79
timestamp 1693479267
transform 1 0 2956 0 1 2505
box -2 -3 18 103
use NAND2X1  NAND2X1_97
timestamp 1693479267
transform 1 0 2972 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_78
timestamp 1693479267
transform 1 0 2996 0 1 2505
box -2 -3 34 103
use FILL  FILL_25_5_0
timestamp 1693479267
transform -1 0 3036 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_5_1
timestamp 1693479267
transform -1 0 3044 0 1 2505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_374
timestamp 1693479267
transform -1 0 3140 0 1 2505
box -2 -3 98 103
use OAI21X1  OAI21X1_74
timestamp 1693479267
transform 1 0 3140 0 1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_354
timestamp 1693479267
transform 1 0 3172 0 1 2505
box -2 -3 98 103
use NAND2X1  NAND2X1_621
timestamp 1693479267
transform 1 0 3268 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_617
timestamp 1693479267
transform 1 0 3292 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_636
timestamp 1693479267
transform 1 0 3316 0 1 2505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_355
timestamp 1693479267
transform 1 0 3340 0 1 2505
box -2 -3 98 103
use NAND2X1  NAND2X1_635
timestamp 1693479267
transform 1 0 3436 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_813
timestamp 1693479267
transform -1 0 3492 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_797
timestamp 1693479267
transform -1 0 3524 0 1 2505
box -2 -3 34 103
use INVX1  INVX1_450
timestamp 1693479267
transform -1 0 3540 0 1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_812
timestamp 1693479267
transform -1 0 3572 0 1 2505
box -2 -3 34 103
use FILL  FILL_25_6_0
timestamp 1693479267
transform -1 0 3580 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_6_1
timestamp 1693479267
transform -1 0 3588 0 1 2505
box -2 -3 10 103
use INVX1  INVX1_466
timestamp 1693479267
transform -1 0 3604 0 1 2505
box -2 -3 18 103
use BUFX4  BUFX4_178
timestamp 1693479267
transform 1 0 3604 0 1 2505
box -2 -3 34 103
use INVX1  INVX1_465
timestamp 1693479267
transform -1 0 3652 0 1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_794
timestamp 1693479267
transform -1 0 3684 0 1 2505
box -2 -3 34 103
use INVX1  INVX1_447
timestamp 1693479267
transform -1 0 3700 0 1 2505
box -2 -3 18 103
use INVX1  INVX1_667
timestamp 1693479267
transform 1 0 3700 0 1 2505
box -2 -3 18 103
use NAND2X1  NAND2X1_930
timestamp 1693479267
transform -1 0 3740 0 1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_442
timestamp 1693479267
transform 1 0 3740 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_971
timestamp 1693479267
transform -1 0 3788 0 1 2505
box -2 -3 26 103
use AND2X2  AND2X2_81
timestamp 1693479267
transform 1 0 3788 0 1 2505
box -2 -3 34 103
use INVX2  INVX2_80
timestamp 1693479267
transform 1 0 3820 0 1 2505
box -2 -3 18 103
use NAND2X1  NAND2X1_982
timestamp 1693479267
transform -1 0 3860 0 1 2505
box -2 -3 26 103
use AND2X2  AND2X2_92
timestamp 1693479267
transform -1 0 3892 0 1 2505
box -2 -3 34 103
use INVX1  INVX1_668
timestamp 1693479267
transform 1 0 3892 0 1 2505
box -2 -3 18 103
use NAND2X1  NAND2X1_933
timestamp 1693479267
transform 1 0 3908 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_935
timestamp 1693479267
transform 1 0 3932 0 1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_253
timestamp 1693479267
transform -1 0 3996 0 1 2505
box -2 -3 34 103
use NOR3X1  NOR3X1_71
timestamp 1693479267
transform -1 0 4060 0 1 2505
box -2 -3 66 103
use OAI21X1  OAI21X1_915
timestamp 1693479267
transform -1 0 4092 0 1 2505
box -2 -3 34 103
use FILL  FILL_25_7_0
timestamp 1693479267
transform 1 0 4092 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_7_1
timestamp 1693479267
transform 1 0 4100 0 1 2505
box -2 -3 10 103
use NOR2X1  NOR2X1_423
timestamp 1693479267
transform 1 0 4108 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_919
timestamp 1693479267
transform 1 0 4132 0 1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_244
timestamp 1693479267
transform 1 0 4164 0 1 2505
box -2 -3 34 103
use AND2X2  AND2X2_97
timestamp 1693479267
transform 1 0 4196 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_979
timestamp 1693479267
transform 1 0 4228 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_920
timestamp 1693479267
transform -1 0 4284 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_451
timestamp 1693479267
transform -1 0 4308 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_980
timestamp 1693479267
transform 1 0 4308 0 1 2505
box -2 -3 26 103
use INVX2  INVX2_84
timestamp 1693479267
transform 1 0 4332 0 1 2505
box -2 -3 18 103
use INVX1  INVX1_682
timestamp 1693479267
transform 1 0 4348 0 1 2505
box -2 -3 18 103
use NAND2X1  NAND2X1_952
timestamp 1693479267
transform -1 0 4388 0 1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_431
timestamp 1693479267
transform 1 0 4388 0 1 2505
box -2 -3 26 103
use INVX1  INVX1_681
timestamp 1693479267
transform 1 0 4412 0 1 2505
box -2 -3 18 103
use AOI21X1  AOI21X1_233
timestamp 1693479267
transform 1 0 4428 0 1 2505
box -2 -3 34 103
use OR2X2  OR2X2_59
timestamp 1693479267
transform 1 0 4460 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_951
timestamp 1693479267
transform 1 0 4492 0 1 2505
box -2 -3 26 103
use AOI22X1  AOI22X1_130
timestamp 1693479267
transform -1 0 4556 0 1 2505
box -2 -3 42 103
use NAND2X1  NAND2X1_950
timestamp 1693479267
transform -1 0 4580 0 1 2505
box -2 -3 26 103
use FILL  FILL_26_1
timestamp 1693479267
transform 1 0 4580 0 1 2505
box -2 -3 10 103
use FILL  FILL_26_2
timestamp 1693479267
transform 1 0 4588 0 1 2505
box -2 -3 10 103
use FILL  FILL_26_3
timestamp 1693479267
transform 1 0 4596 0 1 2505
box -2 -3 10 103
use INVX1  INVX1_183
timestamp 1693479267
transform 1 0 4 0 -1 2705
box -2 -3 18 103
use INVX1  INVX1_180
timestamp 1693479267
transform 1 0 20 0 -1 2705
box -2 -3 18 103
use NOR3X1  NOR3X1_39
timestamp 1693479267
transform -1 0 100 0 -1 2705
box -2 -3 66 103
use NOR3X1  NOR3X1_42
timestamp 1693479267
transform -1 0 164 0 -1 2705
box -2 -3 66 103
use BUFX4  BUFX4_49
timestamp 1693479267
transform -1 0 196 0 -1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_435
timestamp 1693479267
transform 1 0 196 0 -1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_434
timestamp 1693479267
transform 1 0 292 0 -1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_436
timestamp 1693479267
transform 1 0 388 0 -1 2705
box -2 -3 98 103
use NOR2X1  NOR2X1_419
timestamp 1693479267
transform -1 0 508 0 -1 2705
box -2 -3 26 103
use FILL  FILL_26_0_0
timestamp 1693479267
transform -1 0 516 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_0_1
timestamp 1693479267
transform -1 0 524 0 -1 2705
box -2 -3 10 103
use BUFX2  BUFX2_94
timestamp 1693479267
transform -1 0 548 0 -1 2705
box -2 -3 26 103
use BUFX2  BUFX2_95
timestamp 1693479267
transform -1 0 572 0 -1 2705
box -2 -3 26 103
use INVX1  INVX1_651
timestamp 1693479267
transform 1 0 572 0 -1 2705
box -2 -3 18 103
use AOI22X1  AOI22X1_123
timestamp 1693479267
transform 1 0 588 0 -1 2705
box -2 -3 42 103
use NOR2X1  NOR2X1_416
timestamp 1693479267
transform 1 0 628 0 -1 2705
box -2 -3 26 103
use INVX4  INVX4_11
timestamp 1693479267
transform 1 0 652 0 -1 2705
box -2 -3 26 103
use AOI22X1  AOI22X1_121
timestamp 1693479267
transform -1 0 716 0 -1 2705
box -2 -3 42 103
use OAI21X1  OAI21X1_899
timestamp 1693479267
transform -1 0 748 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_897
timestamp 1693479267
transform -1 0 780 0 -1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_331
timestamp 1693479267
transform 1 0 780 0 -1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_311
timestamp 1693479267
transform 1 0 876 0 -1 2705
box -2 -3 98 103
use FILL  FILL_26_1_0
timestamp 1693479267
transform 1 0 972 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_1_1
timestamp 1693479267
transform 1 0 980 0 -1 2705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_329
timestamp 1693479267
transform 1 0 988 0 -1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_142
timestamp 1693479267
transform 1 0 1084 0 -1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_145
timestamp 1693479267
transform 1 0 1180 0 -1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_128
timestamp 1693479267
transform 1 0 1276 0 -1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_16
timestamp 1693479267
transform 1 0 1372 0 -1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_15
timestamp 1693479267
transform 1 0 1468 0 -1 2705
box -2 -3 98 103
use FILL  FILL_26_2_0
timestamp 1693479267
transform 1 0 1564 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_2_1
timestamp 1693479267
transform 1 0 1572 0 -1 2705
box -2 -3 10 103
use OAI21X1  OAI21X1_193
timestamp 1693479267
transform 1 0 1580 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_203
timestamp 1693479267
transform 1 0 1612 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_201
timestamp 1693479267
transform -1 0 1660 0 -1 2705
box -2 -3 18 103
use AOI22X1  AOI22X1_18
timestamp 1693479267
transform -1 0 1700 0 -1 2705
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_88
timestamp 1693479267
transform -1 0 1796 0 -1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_56
timestamp 1693479267
transform -1 0 1892 0 -1 2705
box -2 -3 98 103
use INVX1  INVX1_188
timestamp 1693479267
transform -1 0 1908 0 -1 2705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_78
timestamp 1693479267
transform -1 0 2004 0 -1 2705
box -2 -3 98 103
use FILL  FILL_26_3_0
timestamp 1693479267
transform -1 0 2012 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_3_1
timestamp 1693479267
transform -1 0 2020 0 -1 2705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_222
timestamp 1693479267
transform -1 0 2116 0 -1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_252
timestamp 1693479267
transform -1 0 2212 0 -1 2705
box -2 -3 98 103
use INVX1  INVX1_7
timestamp 1693479267
transform 1 0 2212 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_7
timestamp 1693479267
transform 1 0 2228 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_20
timestamp 1693479267
transform 1 0 2260 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_20
timestamp 1693479267
transform 1 0 2276 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_17
timestamp 1693479267
transform 1 0 2308 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_17
timestamp 1693479267
transform 1 0 2324 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_24
timestamp 1693479267
transform -1 0 2388 0 -1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_232
timestamp 1693479267
transform -1 0 2484 0 -1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_235
timestamp 1693479267
transform -1 0 2580 0 -1 2705
box -2 -3 98 103
use FILL  FILL_26_4_0
timestamp 1693479267
transform 1 0 2580 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_4_1
timestamp 1693479267
transform 1 0 2588 0 -1 2705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_362
timestamp 1693479267
transform 1 0 2596 0 -1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_370
timestamp 1693479267
transform 1 0 2692 0 -1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_369
timestamp 1693479267
transform -1 0 2884 0 -1 2705
box -2 -3 98 103
use OAI21X1  OAI21X1_14
timestamp 1693479267
transform -1 0 2916 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_14
timestamp 1693479267
transform -1 0 2932 0 -1 2705
box -2 -3 18 103
use NAND2X1  NAND2X1_92
timestamp 1693479267
transform 1 0 2932 0 -1 2705
box -2 -3 26 103
use BUFX4  BUFX4_23
timestamp 1693479267
transform -1 0 2988 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_95
timestamp 1693479267
transform -1 0 3020 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_96
timestamp 1693479267
transform -1 0 3036 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_77
timestamp 1693479267
transform -1 0 3068 0 -1 2705
box -2 -3 34 103
use FILL  FILL_26_5_0
timestamp 1693479267
transform -1 0 3076 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_5_1
timestamp 1693479267
transform -1 0 3084 0 -1 2705
box -2 -3 10 103
use INVX1  INVX1_78
timestamp 1693479267
transform -1 0 3100 0 -1 2705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_234
timestamp 1693479267
transform -1 0 3196 0 -1 2705
box -2 -3 98 103
use OAI21X1  OAI21X1_75
timestamp 1693479267
transform -1 0 3228 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_76
timestamp 1693479267
transform 1 0 3228 0 -1 2705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_373
timestamp 1693479267
transform 1 0 3244 0 -1 2705
box -2 -3 98 103
use NAND2X1  NAND2X1_630
timestamp 1693479267
transform 1 0 3340 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_633
timestamp 1693479267
transform 1 0 3364 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_631
timestamp 1693479267
transform 1 0 3388 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_632
timestamp 1693479267
transform 1 0 3412 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_634
timestamp 1693479267
transform 1 0 3436 0 -1 2705
box -2 -3 26 103
use CLKBUF1  CLKBUF1_57
timestamp 1693479267
transform 1 0 3460 0 -1 2705
box -2 -3 74 103
use CLKBUF1  CLKBUF1_46
timestamp 1693479267
transform 1 0 3532 0 -1 2705
box -2 -3 74 103
use FILL  FILL_26_6_0
timestamp 1693479267
transform -1 0 3612 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_6_1
timestamp 1693479267
transform -1 0 3620 0 -1 2705
box -2 -3 10 103
use OAI21X1  OAI21X1_808
timestamp 1693479267
transform -1 0 3652 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_461
timestamp 1693479267
transform -1 0 3668 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_798
timestamp 1693479267
transform -1 0 3700 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_451
timestamp 1693479267
transform -1 0 3716 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_811
timestamp 1693479267
transform -1 0 3748 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_810
timestamp 1693479267
transform -1 0 3780 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_464
timestamp 1693479267
transform -1 0 3796 0 -1 2705
box -2 -3 18 103
use INVX1  INVX1_463
timestamp 1693479267
transform -1 0 3812 0 -1 2705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_387
timestamp 1693479267
transform 1 0 3812 0 -1 2705
box -2 -3 98 103
use OAI21X1  OAI21X1_921
timestamp 1693479267
transform 1 0 3908 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_932
timestamp 1693479267
transform 1 0 3940 0 -1 2705
box -2 -3 26 103
use AOI22X1  AOI22X1_126
timestamp 1693479267
transform -1 0 4004 0 -1 2705
box -2 -3 42 103
use OR2X2  OR2X2_53
timestamp 1693479267
transform -1 0 4036 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_670
timestamp 1693479267
transform 1 0 4036 0 -1 2705
box -2 -3 18 103
use NAND2X1  NAND2X1_937
timestamp 1693479267
transform 1 0 4052 0 -1 2705
box -2 -3 26 103
use FILL  FILL_26_7_0
timestamp 1693479267
transform 1 0 4076 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_7_1
timestamp 1693479267
transform 1 0 4084 0 -1 2705
box -2 -3 10 103
use OAI21X1  OAI21X1_914
timestamp 1693479267
transform 1 0 4092 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_936
timestamp 1693479267
transform 1 0 4124 0 -1 2705
box -2 -3 26 103
use AND2X2  AND2X2_82
timestamp 1693479267
transform 1 0 4148 0 -1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_331
timestamp 1693479267
transform -1 0 4212 0 -1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_232
timestamp 1693479267
transform -1 0 4244 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_669
timestamp 1693479267
transform 1 0 4244 0 -1 2705
box -2 -3 18 103
use INVX1  INVX1_702
timestamp 1693479267
transform 1 0 4260 0 -1 2705
box -2 -3 18 103
use OAI22X1  OAI22X1_51
timestamp 1693479267
transform 1 0 4276 0 -1 2705
box -2 -3 42 103
use NOR2X1  NOR2X1_444
timestamp 1693479267
transform -1 0 4340 0 -1 2705
box -2 -3 26 103
use INVX1  INVX1_703
timestamp 1693479267
transform -1 0 4356 0 -1 2705
box -2 -3 18 103
use AND2X2  AND2X2_90
timestamp 1693479267
transform -1 0 4388 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_935
timestamp 1693479267
transform -1 0 4412 0 -1 2705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_216
timestamp 1693479267
transform -1 0 4508 0 -1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_201
timestamp 1693479267
transform 1 0 4508 0 -1 2705
box -2 -3 98 103
use INVX1  INVX1_182
timestamp 1693479267
transform 1 0 4 0 1 2705
box -2 -3 18 103
use INVX1  INVX1_184
timestamp 1693479267
transform 1 0 20 0 1 2705
box -2 -3 18 103
use NOR3X1  NOR3X1_41
timestamp 1693479267
transform -1 0 100 0 1 2705
box -2 -3 66 103
use NOR3X1  NOR3X1_43
timestamp 1693479267
transform -1 0 164 0 1 2705
box -2 -3 66 103
use DFFPOSX1  DFFPOSX1_432
timestamp 1693479267
transform 1 0 164 0 1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_335
timestamp 1693479267
transform 1 0 260 0 1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_336
timestamp 1693479267
transform 1 0 356 0 1 2705
box -2 -3 98 103
use NAND2X1  NAND2X1_927
timestamp 1693479267
transform 1 0 452 0 1 2705
box -2 -3 26 103
use FILL  FILL_27_0_0
timestamp 1693479267
transform -1 0 484 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_0_1
timestamp 1693479267
transform -1 0 492 0 1 2705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_337
timestamp 1693479267
transform -1 0 588 0 1 2705
box -2 -3 98 103
use AOI22X1  AOI22X1_119
timestamp 1693479267
transform 1 0 588 0 1 2705
box -2 -3 42 103
use OAI21X1  OAI21X1_895
timestamp 1693479267
transform -1 0 660 0 1 2705
box -2 -3 34 103
use BUFX4  BUFX4_261
timestamp 1693479267
transform -1 0 692 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_892
timestamp 1693479267
transform -1 0 724 0 1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_303
timestamp 1693479267
transform 1 0 724 0 1 2705
box -2 -3 98 103
use OAI21X1  OAI21X1_893
timestamp 1693479267
transform -1 0 852 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_891
timestamp 1693479267
transform -1 0 884 0 1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_323
timestamp 1693479267
transform 1 0 884 0 1 2705
box -2 -3 98 103
use FILL  FILL_27_1_0
timestamp 1693479267
transform 1 0 980 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_1_1
timestamp 1693479267
transform 1 0 988 0 1 2705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_325
timestamp 1693479267
transform 1 0 996 0 1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_327
timestamp 1693479267
transform 1 0 1092 0 1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_120
timestamp 1693479267
transform 1 0 1188 0 1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_8
timestamp 1693479267
transform 1 0 1284 0 1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_135
timestamp 1693479267
transform 1 0 1380 0 1 2705
box -2 -3 98 103
use FILL  FILL_27_2_0
timestamp 1693479267
transform 1 0 1476 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_2_1
timestamp 1693479267
transform 1 0 1484 0 1 2705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_23
timestamp 1693479267
transform 1 0 1492 0 1 2705
box -2 -3 98 103
use AOI22X1  AOI22X1_8
timestamp 1693479267
transform -1 0 1628 0 1 2705
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_46
timestamp 1693479267
transform -1 0 1724 0 1 2705
box -2 -3 98 103
use AOI22X1  AOI22X1_23
timestamp 1693479267
transform -1 0 1764 0 1 2705
box -2 -3 42 103
use AOI22X1  AOI22X1_16
timestamp 1693479267
transform -1 0 1804 0 1 2705
box -2 -3 42 103
use AOI22X1  AOI22X1_17
timestamp 1693479267
transform -1 0 1844 0 1 2705
box -2 -3 42 103
use INVX1  INVX1_200
timestamp 1693479267
transform 1 0 1844 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_202
timestamp 1693479267
transform 1 0 1860 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_109
timestamp 1693479267
transform 1 0 1892 0 1 2705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_54
timestamp 1693479267
transform -1 0 2004 0 1 2705
box -2 -3 98 103
use FILL  FILL_27_3_0
timestamp 1693479267
transform -1 0 2012 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_3_1
timestamp 1693479267
transform -1 0 2020 0 1 2705
box -2 -3 10 103
use CLKBUF1  CLKBUF1_15
timestamp 1693479267
transform -1 0 2092 0 1 2705
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_61
timestamp 1693479267
transform -1 0 2188 0 1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_247
timestamp 1693479267
transform -1 0 2284 0 1 2705
box -2 -3 98 103
use NAND2X1  NAND2X1_89
timestamp 1693479267
transform 1 0 2284 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_87
timestamp 1693479267
transform 1 0 2308 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_20
timestamp 1693479267
transform 1 0 2340 0 1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_22
timestamp 1693479267
transform 1 0 2364 0 1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_3
timestamp 1693479267
transform 1 0 2388 0 1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_17
timestamp 1693479267
transform 1 0 2412 0 1 2705
box -2 -3 26 103
use INVX1  INVX1_6
timestamp 1693479267
transform 1 0 2436 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_6
timestamp 1693479267
transform 1 0 2452 0 1 2705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_21
timestamp 1693479267
transform 1 0 2484 0 1 2705
box -2 -3 74 103
use FILL  FILL_27_4_0
timestamp 1693479267
transform 1 0 2556 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_4_1
timestamp 1693479267
transform 1 0 2564 0 1 2705
box -2 -3 10 103
use INVX1  INVX1_15
timestamp 1693479267
transform 1 0 2572 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_15
timestamp 1693479267
transform 1 0 2588 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_19
timestamp 1693479267
transform 1 0 2620 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_19
timestamp 1693479267
transform 1 0 2636 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_27
timestamp 1693479267
transform 1 0 2668 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_27
timestamp 1693479267
transform 1 0 2684 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_16
timestamp 1693479267
transform 1 0 2716 0 1 2705
box -2 -3 26 103
use BUFX4  BUFX4_19
timestamp 1693479267
transform -1 0 2772 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_8
timestamp 1693479267
transform -1 0 2796 0 1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_13
timestamp 1693479267
transform 1 0 2796 0 1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_7
timestamp 1693479267
transform 1 0 2820 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_9
timestamp 1693479267
transform -1 0 2876 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_9
timestamp 1693479267
transform -1 0 2892 0 1 2705
box -2 -3 18 103
use NAND2X1  NAND2X1_14
timestamp 1693479267
transform 1 0 2892 0 1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_75
timestamp 1693479267
transform 1 0 2916 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_90
timestamp 1693479267
transform -1 0 2972 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_91
timestamp 1693479267
transform -1 0 2988 0 1 2705
box -2 -3 18 103
use NAND2X1  NAND2X1_67
timestamp 1693479267
transform 1 0 2988 0 1 2705
box -2 -3 26 103
use BUFX4  BUFX4_163
timestamp 1693479267
transform -1 0 3044 0 1 2705
box -2 -3 34 103
use FILL  FILL_27_5_0
timestamp 1693479267
transform -1 0 3052 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_5_1
timestamp 1693479267
transform -1 0 3060 0 1 2705
box -2 -3 10 103
use OAI21X1  OAI21X1_65
timestamp 1693479267
transform -1 0 3092 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_65
timestamp 1693479267
transform -1 0 3108 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_31
timestamp 1693479267
transform -1 0 3140 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_31
timestamp 1693479267
transform -1 0 3156 0 1 2705
box -2 -3 18 103
use INVX1  INVX1_11
timestamp 1693479267
transform 1 0 3156 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_11
timestamp 1693479267
transform 1 0 3172 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_28
timestamp 1693479267
transform 1 0 3204 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_28
timestamp 1693479267
transform 1 0 3220 0 1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_371
timestamp 1693479267
transform 1 0 3252 0 1 2705
box -2 -3 98 103
use OAI21X1  OAI21X1_12
timestamp 1693479267
transform -1 0 3380 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_12
timestamp 1693479267
transform -1 0 3396 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_29
timestamp 1693479267
transform -1 0 3428 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_29
timestamp 1693479267
transform -1 0 3444 0 1 2705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_386
timestamp 1693479267
transform 1 0 3444 0 1 2705
box -2 -3 98 103
use FILL  FILL_27_6_0
timestamp 1693479267
transform 1 0 3540 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_6_1
timestamp 1693479267
transform 1 0 3548 0 1 2705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_372
timestamp 1693479267
transform 1 0 3556 0 1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_397
timestamp 1693479267
transform 1 0 3652 0 1 2705
box -2 -3 98 103
use OAI21X1  OAI21X1_807
timestamp 1693479267
transform -1 0 3780 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_460
timestamp 1693479267
transform -1 0 3796 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_809
timestamp 1693479267
transform -1 0 3828 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_462
timestamp 1693479267
transform -1 0 3844 0 1 2705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_402
timestamp 1693479267
transform 1 0 3844 0 1 2705
box -2 -3 98 103
use INVX1  INVX1_704
timestamp 1693479267
transform 1 0 3940 0 1 2705
box -2 -3 18 103
use NOR2X1  NOR2X1_453
timestamp 1693479267
transform -1 0 3980 0 1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_931
timestamp 1693479267
transform -1 0 4004 0 1 2705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_378
timestamp 1693479267
transform 1 0 4004 0 1 2705
box -2 -3 98 103
use FILL  FILL_27_7_0
timestamp 1693479267
transform 1 0 4100 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_7_1
timestamp 1693479267
transform 1 0 4108 0 1 2705
box -2 -3 10 103
use INVX2  INVX2_81
timestamp 1693479267
transform 1 0 4116 0 1 2705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_158
timestamp 1693479267
transform 1 0 4132 0 1 2705
box -2 -3 98 103
use AND2X2  AND2X2_89
timestamp 1693479267
transform 1 0 4228 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_443
timestamp 1693479267
transform -1 0 4284 0 1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_934
timestamp 1693479267
transform 1 0 4284 0 1 2705
box -2 -3 26 103
use OR2X2  OR2X2_54
timestamp 1693479267
transform 1 0 4308 0 1 2705
box -2 -3 34 103
use AOI22X1  AOI22X1_127
timestamp 1693479267
transform 1 0 4340 0 1 2705
box -2 -3 42 103
use OR2X2  OR2X2_55
timestamp 1693479267
transform -1 0 4412 0 1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_211
timestamp 1693479267
transform -1 0 4508 0 1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_200
timestamp 1693479267
transform 1 0 4508 0 1 2705
box -2 -3 98 103
use INVX1  INVX1_177
timestamp 1693479267
transform 1 0 4 0 -1 2905
box -2 -3 18 103
use NOR3X1  NOR3X1_36
timestamp 1693479267
transform -1 0 84 0 -1 2905
box -2 -3 66 103
use INVX1  INVX1_159
timestamp 1693479267
transform 1 0 84 0 -1 2905
box -2 -3 18 103
use NOR3X1  NOR3X1_19
timestamp 1693479267
transform -1 0 164 0 -1 2905
box -2 -3 66 103
use DFFPOSX1  DFFPOSX1_411
timestamp 1693479267
transform 1 0 164 0 -1 2905
box -2 -3 98 103
use NOR3X1  NOR3X1_13
timestamp 1693479267
transform -1 0 324 0 -1 2905
box -2 -3 66 103
use INVX1  INVX1_152
timestamp 1693479267
transform -1 0 340 0 -1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_289
timestamp 1693479267
transform 1 0 340 0 -1 2905
box -2 -3 98 103
use INVX2  INVX2_79
timestamp 1693479267
transform 1 0 436 0 -1 2905
box -2 -3 18 103
use NOR2X1  NOR2X1_411
timestamp 1693479267
transform -1 0 476 0 -1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_918
timestamp 1693479267
transform 1 0 476 0 -1 2905
box -2 -3 26 103
use FILL  FILL_28_0_0
timestamp 1693479267
transform 1 0 500 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_0_1
timestamp 1693479267
transform 1 0 508 0 -1 2905
box -2 -3 10 103
use AOI21X1  AOI21X1_230
timestamp 1693479267
transform 1 0 516 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_882
timestamp 1693479267
transform 1 0 548 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_917
timestamp 1693479267
transform 1 0 580 0 -1 2905
box -2 -3 26 103
use INVX1  INVX1_642
timestamp 1693479267
transform -1 0 620 0 -1 2905
box -2 -3 18 103
use NOR3X1  NOR3X1_69
timestamp 1693479267
transform -1 0 684 0 -1 2905
box -2 -3 66 103
use OAI21X1  OAI21X1_894
timestamp 1693479267
transform -1 0 716 0 -1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_326
timestamp 1693479267
transform 1 0 716 0 -1 2905
box -2 -3 98 103
use NOR2X1  NOR2X1_7
timestamp 1693479267
transform -1 0 836 0 -1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_102
timestamp 1693479267
transform -1 0 860 0 -1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_5
timestamp 1693479267
transform 1 0 860 0 -1 2905
box -2 -3 26 103
use AND2X2  AND2X2_1
timestamp 1693479267
transform 1 0 884 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_66
timestamp 1693479267
transform 1 0 916 0 -1 2905
box -2 -3 18 103
use NOR2X1  NOR2X1_1
timestamp 1693479267
transform -1 0 956 0 -1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_66
timestamp 1693479267
transform 1 0 956 0 -1 2905
box -2 -3 26 103
use FILL  FILL_28_1_0
timestamp 1693479267
transform 1 0 980 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_1_1
timestamp 1693479267
transform 1 0 988 0 -1 2905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_134
timestamp 1693479267
transform 1 0 996 0 -1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_126
timestamp 1693479267
transform -1 0 1188 0 -1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_30
timestamp 1693479267
transform 1 0 1188 0 -1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_33
timestamp 1693479267
transform 1 0 1284 0 -1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_147
timestamp 1693479267
transform -1 0 1476 0 -1 2905
box -2 -3 98 103
use FILL  FILL_28_2_0
timestamp 1693479267
transform -1 0 1484 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_2_1
timestamp 1693479267
transform -1 0 1492 0 -1 2905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_100
timestamp 1693479267
transform -1 0 1588 0 -1 2905
box -2 -3 98 103
use OAI21X1  OAI21X1_223
timestamp 1693479267
transform 1 0 1588 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_221
timestamp 1693479267
transform -1 0 1636 0 -1 2905
box -2 -3 18 103
use AOI22X1  AOI22X1_38
timestamp 1693479267
transform -1 0 1676 0 -1 2905
box -2 -3 42 103
use CLKBUF1  CLKBUF1_50
timestamp 1693479267
transform -1 0 1748 0 -1 2905
box -2 -3 74 103
use OAI21X1  OAI21X1_208
timestamp 1693479267
transform -1 0 1780 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_201
timestamp 1693479267
transform -1 0 1812 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_199
timestamp 1693479267
transform -1 0 1828 0 -1 2905
box -2 -3 18 103
use INVX1  INVX1_206
timestamp 1693479267
transform -1 0 1844 0 -1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_108
timestamp 1693479267
transform -1 0 1940 0 -1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_238
timestamp 1693479267
transform -1 0 2036 0 -1 2905
box -2 -3 98 103
use FILL  FILL_28_3_0
timestamp 1693479267
transform -1 0 2044 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_3_1
timestamp 1693479267
transform -1 0 2052 0 -1 2905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_93
timestamp 1693479267
transform -1 0 2148 0 -1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_86
timestamp 1693479267
transform -1 0 2244 0 -1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_233
timestamp 1693479267
transform -1 0 2340 0 -1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_237
timestamp 1693479267
transform -1 0 2436 0 -1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_230
timestamp 1693479267
transform -1 0 2532 0 -1 2905
box -2 -3 98 103
use NAND2X1  NAND2X1_91
timestamp 1693479267
transform -1 0 2556 0 -1 2905
box -2 -3 26 103
use FILL  FILL_28_4_0
timestamp 1693479267
transform -1 0 2564 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_4_1
timestamp 1693479267
transform -1 0 2572 0 -1 2905
box -2 -3 10 103
use BUFX4  BUFX4_161
timestamp 1693479267
transform -1 0 2604 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_83
timestamp 1693479267
transform 1 0 2604 0 -1 2905
box -2 -3 26 103
use INVX1  INVX1_82
timestamp 1693479267
transform 1 0 2628 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_81
timestamp 1693479267
transform 1 0 2644 0 -1 2905
box -2 -3 34 103
use BUFX4  BUFX4_157
timestamp 1693479267
transform -1 0 2708 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_71
timestamp 1693479267
transform 1 0 2708 0 -1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_69
timestamp 1693479267
transform 1 0 2732 0 -1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_81
timestamp 1693479267
transform 1 0 2756 0 -1 2905
box -2 -3 26 103
use BUFX4  BUFX4_160
timestamp 1693479267
transform -1 0 2812 0 -1 2905
box -2 -3 34 103
use BUFX4  BUFX4_17
timestamp 1693479267
transform 1 0 2812 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_26
timestamp 1693479267
transform -1 0 2876 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_26
timestamp 1693479267
transform -1 0 2892 0 -1 2905
box -2 -3 18 103
use NAND2X1  NAND2X1_73
timestamp 1693479267
transform 1 0 2892 0 -1 2905
box -2 -3 26 103
use BUFX4  BUFX4_159
timestamp 1693479267
transform -1 0 2948 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_73
timestamp 1693479267
transform -1 0 2980 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_74
timestamp 1693479267
transform 1 0 2980 0 -1 2905
box -2 -3 18 103
use NAND2X1  NAND2X1_1
timestamp 1693479267
transform -1 0 3020 0 -1 2905
box -2 -3 26 103
use BUFX4  BUFX4_162
timestamp 1693479267
transform -1 0 3052 0 -1 2905
box -2 -3 34 103
use FILL  FILL_28_5_0
timestamp 1693479267
transform 1 0 3052 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_5_1
timestamp 1693479267
transform 1 0 3060 0 -1 2905
box -2 -3 10 103
use INVX1  INVX1_32
timestamp 1693479267
transform 1 0 3068 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_32
timestamp 1693479267
transform 1 0 3084 0 -1 2905
box -2 -3 34 103
use BUFX4  BUFX4_20
timestamp 1693479267
transform -1 0 3148 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_30
timestamp 1693479267
transform 1 0 3148 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_30
timestamp 1693479267
transform 1 0 3164 0 -1 2905
box -2 -3 34 103
use BUFX4  BUFX4_22
timestamp 1693479267
transform 1 0 3196 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_94
timestamp 1693479267
transform -1 0 3252 0 -1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_78
timestamp 1693479267
transform 1 0 3252 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_76
timestamp 1693479267
transform -1 0 3308 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_77
timestamp 1693479267
transform -1 0 3324 0 -1 2905
box -2 -3 18 103
use INVX1  INVX1_93
timestamp 1693479267
transform -1 0 3340 0 -1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_249
timestamp 1693479267
transform -1 0 3436 0 -1 2905
box -2 -3 98 103
use OAI21X1  OAI21X1_43
timestamp 1693479267
transform -1 0 3468 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_43
timestamp 1693479267
transform -1 0 3484 0 -1 2905
box -2 -3 18 103
use NAND2X1  NAND2X1_35
timestamp 1693479267
transform -1 0 3508 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_63
timestamp 1693479267
transform -1 0 3540 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_63
timestamp 1693479267
transform -1 0 3556 0 -1 2905
box -2 -3 18 103
use FILL  FILL_28_6_0
timestamp 1693479267
transform 1 0 3556 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_6_1
timestamp 1693479267
transform 1 0 3564 0 -1 2905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_406
timestamp 1693479267
transform 1 0 3572 0 -1 2905
box -2 -3 98 103
use OAI21X1  OAI21X1_59
timestamp 1693479267
transform -1 0 3700 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_59
timestamp 1693479267
transform -1 0 3716 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_44
timestamp 1693479267
transform 1 0 3716 0 -1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_403
timestamp 1693479267
transform 1 0 3748 0 -1 2905
box -2 -3 98 103
use OAI21X1  OAI21X1_45
timestamp 1693479267
transform -1 0 3876 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_45
timestamp 1693479267
transform -1 0 3892 0 -1 2905
box -2 -3 18 103
use INVX1  INVX1_35
timestamp 1693479267
transform 1 0 3892 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_35
timestamp 1693479267
transform 1 0 3908 0 -1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_388
timestamp 1693479267
transform 1 0 3940 0 -1 2905
box -2 -3 98 103
use FILL  FILL_28_7_0
timestamp 1693479267
transform 1 0 4036 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_7_1
timestamp 1693479267
transform 1 0 4044 0 -1 2905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_218
timestamp 1693479267
transform 1 0 4052 0 -1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_192
timestamp 1693479267
transform 1 0 4148 0 -1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_220
timestamp 1693479267
transform 1 0 4244 0 -1 2905
box -2 -3 98 103
use NAND2X1  NAND2X1_1028
timestamp 1693479267
transform 1 0 4340 0 -1 2905
box -2 -3 26 103
use BUFX2  BUFX2_79
timestamp 1693479267
transform -1 0 4388 0 -1 2905
box -2 -3 26 103
use AOI22X1  AOI22X1_168
timestamp 1693479267
transform 1 0 4388 0 -1 2905
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_217
timestamp 1693479267
transform 1 0 4428 0 -1 2905
box -2 -3 98 103
use NAND2X1  NAND2X1_1026
timestamp 1693479267
transform 1 0 4524 0 -1 2905
box -2 -3 26 103
use NAND3X1  NAND3X1_361
timestamp 1693479267
transform 1 0 4548 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_1027
timestamp 1693479267
transform -1 0 4604 0 -1 2905
box -2 -3 26 103
use INVX1  INVX1_163
timestamp 1693479267
transform 1 0 4 0 1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_429
timestamp 1693479267
transform 1 0 20 0 1 2905
box -2 -3 98 103
use NOR3X1  NOR3X1_22
timestamp 1693479267
transform -1 0 180 0 1 2905
box -2 -3 66 103
use CLKBUF1  CLKBUF1_20
timestamp 1693479267
transform -1 0 252 0 1 2905
box -2 -3 74 103
use BUFX4  BUFX4_45
timestamp 1693479267
transform 1 0 252 0 1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_415
timestamp 1693479267
transform 1 0 284 0 1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_286
timestamp 1693479267
transform 1 0 380 0 1 2905
box -2 -3 98 103
use NAND2X1  NAND2X1_925
timestamp 1693479267
transform 1 0 476 0 1 2905
box -2 -3 26 103
use FILL  FILL_29_0_0
timestamp 1693479267
transform -1 0 508 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_0_1
timestamp 1693479267
transform -1 0 516 0 1 2905
box -2 -3 10 103
use OAI21X1  OAI21X1_881
timestamp 1693479267
transform -1 0 548 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_926
timestamp 1693479267
transform -1 0 572 0 1 2905
box -2 -3 26 103
use NAND3X1  NAND3X1_327
timestamp 1693479267
transform 1 0 572 0 1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_231
timestamp 1693479267
transform -1 0 636 0 1 2905
box -2 -3 34 103
use AOI22X1  AOI22X1_118
timestamp 1693479267
transform 1 0 636 0 1 2905
box -2 -3 42 103
use AOI22X1  AOI22X1_116
timestamp 1693479267
transform 1 0 676 0 1 2905
box -2 -3 42 103
use BUFX4  BUFX4_262
timestamp 1693479267
transform 1 0 716 0 1 2905
box -2 -3 34 103
use AOI22X1  AOI22X1_117
timestamp 1693479267
transform -1 0 788 0 1 2905
box -2 -3 42 103
use AOI22X1  AOI22X1_115
timestamp 1693479267
transform -1 0 828 0 1 2905
box -2 -3 42 103
use CLKBUF1  CLKBUF1_49
timestamp 1693479267
transform 1 0 828 0 1 2905
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_314
timestamp 1693479267
transform 1 0 900 0 1 2905
box -2 -3 98 103
use NAND2X1  NAND2X1_65
timestamp 1693479267
transform 1 0 996 0 1 2905
box -2 -3 26 103
use FILL  FILL_29_1_0
timestamp 1693479267
transform 1 0 1020 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_1_1
timestamp 1693479267
transform 1 0 1028 0 1 2905
box -2 -3 10 103
use OR2X2  OR2X2_1
timestamp 1693479267
transform 1 0 1036 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_2
timestamp 1693479267
transform -1 0 1092 0 1 2905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_144
timestamp 1693479267
transform 1 0 1092 0 1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_131
timestamp 1693479267
transform 1 0 1188 0 1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_35
timestamp 1693479267
transform -1 0 1380 0 1 2905
box -2 -3 98 103
use AOI22X1  AOI22X1_30
timestamp 1693479267
transform -1 0 1420 0 1 2905
box -2 -3 42 103
use OAI21X1  OAI21X1_215
timestamp 1693479267
transform -1 0 1452 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_213
timestamp 1693479267
transform -1 0 1468 0 1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_68
timestamp 1693479267
transform -1 0 1564 0 1 2905
box -2 -3 98 103
use FILL  FILL_29_2_0
timestamp 1693479267
transform -1 0 1572 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_2_1
timestamp 1693479267
transform -1 0 1580 0 1 2905
box -2 -3 10 103
use INVX1  INVX1_203
timestamp 1693479267
transform -1 0 1596 0 1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_90
timestamp 1693479267
transform -1 0 1692 0 1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_76
timestamp 1693479267
transform -1 0 1788 0 1 2905
box -2 -3 98 103
use BUFX4  BUFX4_258
timestamp 1693479267
transform -1 0 1820 0 1 2905
box -2 -3 34 103
use BUFX4  BUFX4_236
timestamp 1693479267
transform -1 0 1852 0 1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_245
timestamp 1693479267
transform -1 0 1948 0 1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_55
timestamp 1693479267
transform -1 0 2044 0 1 2905
box -2 -3 98 103
use FILL  FILL_29_3_0
timestamp 1693479267
transform -1 0 2052 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_3_1
timestamp 1693479267
transform -1 0 2060 0 1 2905
box -2 -3 10 103
use CLKBUF1  CLKBUF1_63
timestamp 1693479267
transform -1 0 2132 0 1 2905
box -2 -3 74 103
use INVX1  INVX1_121
timestamp 1693479267
transform 1 0 2132 0 1 2905
box -2 -3 18 103
use INVX1  INVX1_108
timestamp 1693479267
transform 1 0 2148 0 1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_224
timestamp 1693479267
transform -1 0 2260 0 1 2905
box -2 -3 98 103
use NAND2X1  NAND2X1_780
timestamp 1693479267
transform -1 0 2284 0 1 2905
box -2 -3 26 103
use INVX1  INVX1_114
timestamp 1693479267
transform 1 0 2284 0 1 2905
box -2 -3 18 103
use INVX1  INVX1_107
timestamp 1693479267
transform 1 0 2300 0 1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_226
timestamp 1693479267
transform -1 0 2412 0 1 2905
box -2 -3 98 103
use NAND2X1  NAND2X1_717
timestamp 1693479267
transform -1 0 2436 0 1 2905
box -2 -3 26 103
use INVX1  INVX1_89
timestamp 1693479267
transform 1 0 2436 0 1 2905
box -2 -3 18 103
use NAND2X1  NAND2X1_90
timestamp 1693479267
transform 1 0 2452 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_88
timestamp 1693479267
transform 1 0 2476 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_778
timestamp 1693479267
transform -1 0 2532 0 1 2905
box -2 -3 26 103
use FILL  FILL_29_4_0
timestamp 1693479267
transform -1 0 2540 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_4_1
timestamp 1693479267
transform -1 0 2548 0 1 2905
box -2 -3 10 103
use OAI21X1  OAI21X1_89
timestamp 1693479267
transform -1 0 2580 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_90
timestamp 1693479267
transform -1 0 2596 0 1 2905
box -2 -3 18 103
use NAND2X1  NAND2X1_15
timestamp 1693479267
transform 1 0 2596 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_6
timestamp 1693479267
transform 1 0 2620 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_19
timestamp 1693479267
transform -1 0 2668 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_715
timestamp 1693479267
transform -1 0 2692 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_27
timestamp 1693479267
transform -1 0 2716 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_69
timestamp 1693479267
transform -1 0 2748 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_70
timestamp 1693479267
transform -1 0 2764 0 1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_67
timestamp 1693479267
transform -1 0 2796 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_68
timestamp 1693479267
transform -1 0 2812 0 1 2905
box -2 -3 18 103
use NAND2X1  NAND2X1_747
timestamp 1693479267
transform -1 0 2836 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_26
timestamp 1693479267
transform -1 0 2860 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_9
timestamp 1693479267
transform 1 0 2860 0 1 2905
box -2 -3 26 103
use INVX1  INVX1_81
timestamp 1693479267
transform 1 0 2884 0 1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_80
timestamp 1693479267
transform 1 0 2900 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_82
timestamp 1693479267
transform -1 0 2956 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_10
timestamp 1693479267
transform -1 0 2980 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_745
timestamp 1693479267
transform -1 0 3004 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_711
timestamp 1693479267
transform 1 0 3004 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_702
timestamp 1693479267
transform -1 0 3052 0 1 2905
box -2 -3 26 103
use FILL  FILL_29_5_0
timestamp 1693479267
transform -1 0 3060 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_5_1
timestamp 1693479267
transform -1 0 3068 0 1 2905
box -2 -3 10 103
use NAND2X1  NAND2X1_11
timestamp 1693479267
transform -1 0 3092 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_31
timestamp 1693479267
transform -1 0 3116 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_32
timestamp 1693479267
transform -1 0 3140 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_28
timestamp 1693479267
transform -1 0 3164 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_30
timestamp 1693479267
transform 1 0 3164 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_29
timestamp 1693479267
transform 1 0 3188 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_92
timestamp 1693479267
transform -1 0 3244 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_12
timestamp 1693479267
transform 1 0 3244 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_63
timestamp 1693479267
transform -1 0 3292 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_43
timestamp 1693479267
transform -1 0 3316 0 1 2905
box -2 -3 26 103
use INVX1  INVX1_34
timestamp 1693479267
transform 1 0 3316 0 1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_34
timestamp 1693479267
transform 1 0 3332 0 1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_377
timestamp 1693479267
transform 1 0 3364 0 1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_390
timestamp 1693479267
transform 1 0 3460 0 1 2905
box -2 -3 98 103
use FILL  FILL_29_6_0
timestamp 1693479267
transform 1 0 3556 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_6_1
timestamp 1693479267
transform 1 0 3564 0 1 2905
box -2 -3 10 103
use CLKBUF1  CLKBUF1_37
timestamp 1693479267
transform 1 0 3572 0 1 2905
box -2 -3 74 103
use OAI21X1  OAI21X1_60
timestamp 1693479267
transform -1 0 3676 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_60
timestamp 1693479267
transform -1 0 3692 0 1 2905
box -2 -3 18 103
use INVX1  INVX1_44
timestamp 1693479267
transform 1 0 3692 0 1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_50
timestamp 1693479267
transform -1 0 3740 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_50
timestamp 1693479267
transform -1 0 3756 0 1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_393
timestamp 1693479267
transform 1 0 3756 0 1 2905
box -2 -3 98 103
use NAND2X1  NAND2X1_45
timestamp 1693479267
transform -1 0 3876 0 1 2905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_117
timestamp 1693479267
transform -1 0 3972 0 1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_207
timestamp 1693479267
transform 1 0 3972 0 1 2905
box -2 -3 98 103
use INVX1  INVX1_719
timestamp 1693479267
transform 1 0 4068 0 1 2905
box -2 -3 18 103
use FILL  FILL_29_7_0
timestamp 1693479267
transform 1 0 4084 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_7_1
timestamp 1693479267
transform 1 0 4092 0 1 2905
box -2 -3 10 103
use CLKBUF1  CLKBUF1_28
timestamp 1693479267
transform 1 0 4100 0 1 2905
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_204
timestamp 1693479267
transform 1 0 4172 0 1 2905
box -2 -3 98 103
use INVX1  INVX1_732
timestamp 1693479267
transform 1 0 4268 0 1 2905
box -2 -3 18 103
use AOI22X1  AOI22X1_170
timestamp 1693479267
transform 1 0 4284 0 1 2905
box -2 -3 42 103
use OAI21X1  OAI21X1_1052
timestamp 1693479267
transform 1 0 4324 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_723
timestamp 1693479267
transform -1 0 4372 0 1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_202
timestamp 1693479267
transform 1 0 4372 0 1 2905
box -2 -3 98 103
use INVX1  INVX1_728
timestamp 1693479267
transform 1 0 4468 0 1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_970
timestamp 1693479267
transform 1 0 4484 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_730
timestamp 1693479267
transform 1 0 4516 0 1 2905
box -2 -3 18 103
use NAND2X1  NAND2X1_1029
timestamp 1693479267
transform 1 0 4532 0 1 2905
box -2 -3 26 103
use NAND3X1  NAND3X1_362
timestamp 1693479267
transform 1 0 4556 0 1 2905
box -2 -3 34 103
use FILL  FILL_30_1
timestamp 1693479267
transform 1 0 4588 0 1 2905
box -2 -3 10 103
use FILL  FILL_30_2
timestamp 1693479267
transform 1 0 4596 0 1 2905
box -2 -3 10 103
use INVX1  INVX1_157
timestamp 1693479267
transform 1 0 4 0 -1 3105
box -2 -3 18 103
use NAND3X1  NAND3X1_71
timestamp 1693479267
transform -1 0 52 0 -1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_409
timestamp 1693479267
transform 1 0 52 0 -1 3105
box -2 -3 98 103
use INVX1  INVX1_156
timestamp 1693479267
transform 1 0 4 0 1 3105
box -2 -3 18 103
use NAND3X1  NAND3X1_70
timestamp 1693479267
transform -1 0 52 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_160
timestamp 1693479267
transform 1 0 52 0 1 3105
box -2 -3 18 103
use NAND3X1  NAND3X1_72
timestamp 1693479267
transform -1 0 100 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_158
timestamp 1693479267
transform 1 0 100 0 1 3105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_410
timestamp 1693479267
transform 1 0 148 0 -1 3105
box -2 -3 98 103
use NOR3X1  NOR3X1_18
timestamp 1693479267
transform -1 0 180 0 1 3105
box -2 -3 66 103
use INVX1  INVX1_150
timestamp 1693479267
transform 1 0 180 0 1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_108
timestamp 1693479267
transform 1 0 196 0 1 3105
box -2 -3 26 103
use INVX1  INVX1_149
timestamp 1693479267
transform 1 0 244 0 -1 3105
box -2 -3 18 103
use INVX4  INVX4_1
timestamp 1693479267
transform 1 0 260 0 -1 3105
box -2 -3 26 103
use NAND3X1  NAND3X1_5
timestamp 1693479267
transform 1 0 284 0 -1 3105
box -2 -3 34 103
use NAND3X1  NAND3X1_6
timestamp 1693479267
transform -1 0 252 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_153
timestamp 1693479267
transform 1 0 252 0 1 3105
box -2 -3 18 103
use NAND3X1  NAND3X1_7
timestamp 1693479267
transform 1 0 268 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_14
timestamp 1693479267
transform -1 0 324 0 1 3105
box -2 -3 26 103
use INVX1  INVX1_227
timestamp 1693479267
transform -1 0 332 0 -1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_113
timestamp 1693479267
transform 1 0 332 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_110
timestamp 1693479267
transform -1 0 380 0 -1 3105
box -2 -3 26 103
use INVX1  INVX1_226
timestamp 1693479267
transform -1 0 396 0 -1 3105
box -2 -3 18 103
use NOR3X1  NOR3X1_12
timestamp 1693479267
transform -1 0 460 0 -1 3105
box -2 -3 66 103
use NOR2X1  NOR2X1_21
timestamp 1693479267
transform 1 0 324 0 1 3105
box -2 -3 26 103
use NAND3X1  NAND3X1_74
timestamp 1693479267
transform -1 0 380 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_18
timestamp 1693479267
transform -1 0 404 0 1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_16
timestamp 1693479267
transform -1 0 428 0 1 3105
box -2 -3 26 103
use INVX1  INVX1_151
timestamp 1693479267
transform -1 0 476 0 -1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_114
timestamp 1693479267
transform 1 0 476 0 -1 3105
box -2 -3 26 103
use FILL  FILL_30_0_0
timestamp 1693479267
transform -1 0 508 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_0_1
timestamp 1693479267
transform -1 0 516 0 -1 3105
box -2 -3 10 103
use NAND2X1  NAND2X1_115
timestamp 1693479267
transform 1 0 428 0 1 3105
box -2 -3 26 103
use OR2X2  OR2X2_7
timestamp 1693479267
transform 1 0 452 0 1 3105
box -2 -3 34 103
use FILL  FILL_31_0_0
timestamp 1693479267
transform -1 0 492 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_0_1
timestamp 1693479267
transform -1 0 500 0 1 3105
box -2 -3 10 103
use OAI22X1  OAI22X1_6
timestamp 1693479267
transform -1 0 540 0 1 3105
box -2 -3 42 103
use CLKBUF1  CLKBUF1_34
timestamp 1693479267
transform -1 0 588 0 -1 3105
box -2 -3 74 103
use NAND3X1  NAND3X1_326
timestamp 1693479267
transform 1 0 588 0 -1 3105
box -2 -3 34 103
use OR2X2  OR2X2_5
timestamp 1693479267
transform 1 0 540 0 1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_288
timestamp 1693479267
transform 1 0 572 0 1 3105
box -2 -3 98 103
use AOI22X1  AOI22X1_114
timestamp 1693479267
transform -1 0 660 0 -1 3105
box -2 -3 42 103
use NOR2X1  NOR2X1_412
timestamp 1693479267
transform 1 0 660 0 -1 3105
box -2 -3 26 103
use INVX1  INVX1_643
timestamp 1693479267
transform 1 0 684 0 -1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_920
timestamp 1693479267
transform 1 0 700 0 -1 3105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_287
timestamp 1693479267
transform 1 0 668 0 1 3105
box -2 -3 98 103
use OAI22X1  OAI22X1_49
timestamp 1693479267
transform 1 0 724 0 -1 3105
box -2 -3 42 103
use INVX1  INVX1_641
timestamp 1693479267
transform -1 0 780 0 -1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_919
timestamp 1693479267
transform -1 0 804 0 -1 3105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_143
timestamp 1693479267
transform 1 0 804 0 -1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_305
timestamp 1693479267
transform 1 0 764 0 1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_122
timestamp 1693479267
transform 1 0 900 0 -1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_31
timestamp 1693479267
transform 1 0 860 0 1 3105
box -2 -3 98 103
use FILL  FILL_30_1_0
timestamp 1693479267
transform 1 0 996 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_1_1
timestamp 1693479267
transform 1 0 1004 0 -1 3105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_10
timestamp 1693479267
transform 1 0 1012 0 -1 3105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_24
timestamp 1693479267
transform 1 0 956 0 1 3105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_14
timestamp 1693479267
transform 1 0 1108 0 -1 3105
box -2 -3 98 103
use FILL  FILL_31_1_0
timestamp 1693479267
transform 1 0 1028 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_1_1
timestamp 1693479267
transform 1 0 1036 0 1 3105
box -2 -3 10 103
use CLKBUF1  CLKBUF1_11
timestamp 1693479267
transform 1 0 1044 0 1 3105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_32
timestamp 1693479267
transform 1 0 1204 0 -1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_146
timestamp 1693479267
transform -1 0 1212 0 1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_48
timestamp 1693479267
transform 1 0 1212 0 1 3105
box -2 -3 98 103
use AOI22X1  AOI22X1_10
timestamp 1693479267
transform 1 0 1300 0 -1 3105
box -2 -3 42 103
use AOI22X1  AOI22X1_31
timestamp 1693479267
transform 1 0 1308 0 1 3105
box -2 -3 42 103
use BUFX4  BUFX4_256
timestamp 1693479267
transform -1 0 1372 0 -1 3105
box -2 -3 34 103
use AOI22X1  AOI22X1_33
timestamp 1693479267
transform -1 0 1412 0 -1 3105
box -2 -3 42 103
use OAI21X1  OAI21X1_218
timestamp 1693479267
transform -1 0 1444 0 -1 3105
box -2 -3 34 103
use BUFX4  BUFX4_259
timestamp 1693479267
transform -1 0 1380 0 1 3105
box -2 -3 34 103
use BUFX4  BUFX4_238
timestamp 1693479267
transform -1 0 1412 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_216
timestamp 1693479267
transform -1 0 1444 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_216
timestamp 1693479267
transform -1 0 1460 0 -1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_195
timestamp 1693479267
transform -1 0 1492 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_193
timestamp 1693479267
transform -1 0 1508 0 -1 3105
box -2 -3 18 103
use FILL  FILL_30_2_0
timestamp 1693479267
transform -1 0 1516 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_2_1
timestamp 1693479267
transform -1 0 1524 0 -1 3105
box -2 -3 10 103
use BUFX4  BUFX4_144
timestamp 1693479267
transform -1 0 1476 0 1 3105
box -2 -3 34 103
use BUFX4  BUFX4_141
timestamp 1693479267
transform 1 0 1476 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_101
timestamp 1693479267
transform 1 0 1508 0 1 3105
box -2 -3 18 103
use AOI22X1  AOI22X1_20
timestamp 1693479267
transform -1 0 1564 0 -1 3105
box -2 -3 42 103
use OAI21X1  OAI21X1_205
timestamp 1693479267
transform -1 0 1596 0 -1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_80
timestamp 1693479267
transform -1 0 1692 0 -1 3105
box -2 -3 98 103
use FILL  FILL_31_2_0
timestamp 1693479267
transform -1 0 1532 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_2_1
timestamp 1693479267
transform -1 0 1540 0 1 3105
box -2 -3 10 103
use AOI22X1  AOI22X1_21
timestamp 1693479267
transform -1 0 1580 0 1 3105
box -2 -3 42 103
use AOI22X1  AOI22X1_15
timestamp 1693479267
transform -1 0 1620 0 1 3105
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_58
timestamp 1693479267
transform -1 0 1788 0 -1 3105
box -2 -3 98 103
use AOI22X1  AOI22X1_32
timestamp 1693479267
transform -1 0 1660 0 1 3105
box -2 -3 42 103
use OAI21X1  OAI21X1_200
timestamp 1693479267
transform -1 0 1692 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_217
timestamp 1693479267
transform -1 0 1724 0 1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_243
timestamp 1693479267
transform -1 0 1884 0 -1 3105
box -2 -3 98 103
use INVX1  INVX1_198
timestamp 1693479267
transform -1 0 1740 0 1 3105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_85
timestamp 1693479267
transform -1 0 1836 0 1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_103
timestamp 1693479267
transform -1 0 1980 0 -1 3105
box -2 -3 98 103
use INVX1  INVX1_215
timestamp 1693479267
transform -1 0 1852 0 1 3105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_102
timestamp 1693479267
transform -1 0 1948 0 1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_246
timestamp 1693479267
transform -1 0 2076 0 -1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_241
timestamp 1693479267
transform -1 0 2044 0 1 3105
box -2 -3 98 103
use INVX1  INVX1_129
timestamp 1693479267
transform 1 0 2060 0 1 3105
box -2 -3 18 103
use FILL  FILL_31_3_1
timestamp 1693479267
transform 1 0 2052 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_3_0
timestamp 1693479267
transform 1 0 2044 0 1 3105
box -2 -3 10 103
use OAI21X1  OAI21X1_102
timestamp 1693479267
transform 1 0 2092 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_111
timestamp 1693479267
transform 1 0 2076 0 1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_141
timestamp 1693479267
transform 1 0 2092 0 -1 3105
box -2 -3 34 103
use FILL  FILL_30_3_1
timestamp 1693479267
transform 1 0 2084 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_3_0
timestamp 1693479267
transform 1 0 2076 0 -1 3105
box -2 -3 10 103
use OAI21X1  OAI21X1_101
timestamp 1693479267
transform -1 0 2156 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_142
timestamp 1693479267
transform -1 0 2156 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_157
timestamp 1693479267
transform -1 0 2188 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_115
timestamp 1693479267
transform -1 0 2220 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_116
timestamp 1693479267
transform -1 0 2252 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_158
timestamp 1693479267
transform 1 0 2156 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_98
timestamp 1693479267
transform 1 0 2188 0 1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_98
timestamp 1693479267
transform 1 0 2204 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_118
timestamp 1693479267
transform 1 0 2252 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_117
timestamp 1693479267
transform 1 0 2284 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_128
timestamp 1693479267
transform 1 0 2316 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_97
timestamp 1693479267
transform -1 0 2268 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_147
timestamp 1693479267
transform -1 0 2300 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_85
timestamp 1693479267
transform 1 0 2300 0 1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_113
timestamp 1693479267
transform 1 0 2316 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_127
timestamp 1693479267
transform -1 0 2380 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_121
timestamp 1693479267
transform 1 0 2380 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_87
timestamp 1693479267
transform 1 0 2412 0 -1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_114
timestamp 1693479267
transform -1 0 2380 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_122
timestamp 1693479267
transform 1 0 2380 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_774
timestamp 1693479267
transform -1 0 2436 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_88
timestamp 1693479267
transform 1 0 2428 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_86
timestamp 1693479267
transform 1 0 2452 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_772
timestamp 1693479267
transform 1 0 2484 0 -1 3105
box -2 -3 26 103
use INVX1  INVX1_83
timestamp 1693479267
transform 1 0 2508 0 -1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_84
timestamp 1693479267
transform 1 0 2524 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_783
timestamp 1693479267
transform -1 0 2460 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_759
timestamp 1693479267
transform -1 0 2484 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_762
timestamp 1693479267
transform -1 0 2508 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_723
timestamp 1693479267
transform -1 0 2532 0 1 3105
box -2 -3 26 103
use FILL  FILL_31_4_1
timestamp 1693479267
transform -1 0 2572 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_4_0
timestamp 1693479267
transform -1 0 2564 0 1 3105
box -2 -3 10 103
use NAND2X1  NAND2X1_781
timestamp 1693479267
transform -1 0 2556 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_82
timestamp 1693479267
transform 1 0 2564 0 -1 3105
box -2 -3 34 103
use FILL  FILL_30_4_1
timestamp 1693479267
transform 1 0 2556 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_4_0
timestamp 1693479267
transform 1 0 2548 0 -1 3105
box -2 -3 10 103
use BUFX4  BUFX4_272
timestamp 1693479267
transform -1 0 2604 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_760
timestamp 1693479267
transform -1 0 2620 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_757
timestamp 1693479267
transform -1 0 2652 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_753
timestamp 1693479267
transform -1 0 2628 0 1 3105
box -2 -3 26 103
use BUFX4  BUFX4_134
timestamp 1693479267
transform -1 0 2652 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_870
timestamp 1693479267
transform 1 0 2652 0 -1 3105
box -2 -3 26 103
use INVX1  INVX1_92
timestamp 1693479267
transform 1 0 2676 0 -1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_91
timestamp 1693479267
transform 1 0 2692 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_93
timestamp 1693479267
transform -1 0 2748 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_872
timestamp 1693479267
transform -1 0 2676 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_721
timestamp 1693479267
transform -1 0 2700 0 1 3105
box -2 -3 26 103
use BUFX4  BUFX4_60
timestamp 1693479267
transform -1 0 2732 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_825
timestamp 1693479267
transform -1 0 2772 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_79
timestamp 1693479267
transform -1 0 2804 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_80
timestamp 1693479267
transform -1 0 2820 0 -1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_730
timestamp 1693479267
transform 1 0 2820 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_751
timestamp 1693479267
transform -1 0 2756 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_827
timestamp 1693479267
transform 1 0 2756 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_732
timestamp 1693479267
transform -1 0 2804 0 1 3105
box -2 -3 26 103
use BUFX4  BUFX4_135
timestamp 1693479267
transform 1 0 2804 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_72
timestamp 1693479267
transform 1 0 2844 0 -1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_784
timestamp 1693479267
transform -1 0 2884 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_894
timestamp 1693479267
transform -1 0 2908 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_71
timestamp 1693479267
transform 1 0 2908 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_786
timestamp 1693479267
transform -1 0 2860 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_896
timestamp 1693479267
transform -1 0 2884 0 1 3105
box -2 -3 26 103
use BUFX4  BUFX4_131
timestamp 1693479267
transform 1 0 2884 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_750
timestamp 1693479267
transform -1 0 2940 0 1 3105
box -2 -3 26 103
use BUFX4  BUFX4_132
timestamp 1693479267
transform 1 0 2940 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_748
timestamp 1693479267
transform -1 0 2996 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_799
timestamp 1693479267
transform 1 0 2996 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_909
timestamp 1693479267
transform 1 0 3020 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_738
timestamp 1693479267
transform -1 0 2964 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_736
timestamp 1693479267
transform -1 0 2988 0 1 3105
box -2 -3 26 103
use BUFX4  BUFX4_61
timestamp 1693479267
transform 1 0 2988 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_741
timestamp 1693479267
transform -1 0 3044 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_801
timestamp 1693479267
transform 1 0 3044 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_739
timestamp 1693479267
transform -1 0 3068 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_911
timestamp 1693479267
transform 1 0 3084 0 1 3105
box -2 -3 26 103
use FILL  FILL_31_5_1
timestamp 1693479267
transform 1 0 3076 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_5_0
timestamp 1693479267
transform 1 0 3068 0 1 3105
box -2 -3 10 103
use NAND2X1  NAND2X1_858
timestamp 1693479267
transform 1 0 3084 0 -1 3105
box -2 -3 26 103
use FILL  FILL_30_5_1
timestamp 1693479267
transform 1 0 3076 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_5_0
timestamp 1693479267
transform 1 0 3068 0 -1 3105
box -2 -3 10 103
use NAND2X1  NAND2X1_790
timestamp 1693479267
transform -1 0 3132 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_849
timestamp 1693479267
transform 1 0 3108 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_792
timestamp 1693479267
transform 1 0 3132 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_851
timestamp 1693479267
transform 1 0 3132 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_882
timestamp 1693479267
transform 1 0 3156 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_855
timestamp 1693479267
transform 1 0 3180 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_812
timestamp 1693479267
transform 1 0 3204 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_900
timestamp 1693479267
transform 1 0 3228 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_884
timestamp 1693479267
transform -1 0 3180 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_857
timestamp 1693479267
transform -1 0 3204 0 1 3105
box -2 -3 26 103
use BUFX4  BUFX4_59
timestamp 1693479267
transform -1 0 3236 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_54
timestamp 1693479267
transform -1 0 3276 0 -1 3105
box -2 -3 26 103
use INVX1  INVX1_54
timestamp 1693479267
transform -1 0 3292 0 -1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_54
timestamp 1693479267
transform 1 0 3292 0 -1 3105
box -2 -3 34 103
use BUFX4  BUFX4_30
timestamp 1693479267
transform 1 0 3324 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_50
timestamp 1693479267
transform -1 0 3260 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_34
timestamp 1693479267
transform -1 0 3284 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_47
timestamp 1693479267
transform -1 0 3308 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_902
timestamp 1693479267
transform 1 0 3308 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_60
timestamp 1693479267
transform -1 0 3356 0 1 3105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_394
timestamp 1693479267
transform 1 0 3356 0 -1 3105
box -2 -3 98 103
use OAI21X1  OAI21X1_37
timestamp 1693479267
transform -1 0 3388 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_37
timestamp 1693479267
transform -1 0 3404 0 1 3105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_380
timestamp 1693479267
transform 1 0 3404 0 1 3105
box -2 -3 98 103
use INVX1  INVX1_47
timestamp 1693479267
transform 1 0 3452 0 -1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_47
timestamp 1693479267
transform -1 0 3500 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_58
timestamp 1693479267
transform -1 0 3524 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_58
timestamp 1693479267
transform -1 0 3556 0 -1 3105
box -2 -3 34 103
use BUFX4  BUFX4_29
timestamp 1693479267
transform 1 0 3500 0 1 3105
box -2 -3 34 103
use FILL  FILL_31_6_0
timestamp 1693479267
transform 1 0 3532 0 1 3105
box -2 -3 10 103
use INVX1  INVX1_58
timestamp 1693479267
transform -1 0 3572 0 -1 3105
box -2 -3 18 103
use FILL  FILL_30_6_0
timestamp 1693479267
transform 1 0 3572 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_6_1
timestamp 1693479267
transform 1 0 3580 0 -1 3105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_401
timestamp 1693479267
transform 1 0 3588 0 -1 3105
box -2 -3 98 103
use FILL  FILL_31_6_1
timestamp 1693479267
transform 1 0 3540 0 1 3105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_392
timestamp 1693479267
transform 1 0 3548 0 1 3105
box -2 -3 98 103
use BUFX4  BUFX4_26
timestamp 1693479267
transform 1 0 3684 0 -1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_404
timestamp 1693479267
transform 1 0 3716 0 -1 3105
box -2 -3 98 103
use NAND2X1  NAND2X1_44
timestamp 1693479267
transform -1 0 3668 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_62
timestamp 1693479267
transform -1 0 3700 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_62
timestamp 1693479267
transform -1 0 3716 0 1 3105
box -2 -3 18 103
use INVX1  INVX1_38
timestamp 1693479267
transform 1 0 3716 0 1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_38
timestamp 1693479267
transform 1 0 3732 0 1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_119
timestamp 1693479267
transform -1 0 3908 0 -1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_405
timestamp 1693479267
transform -1 0 3860 0 1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_191
timestamp 1693479267
transform 1 0 3908 0 -1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_381
timestamp 1693479267
transform 1 0 3860 0 1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_208
timestamp 1693479267
transform 1 0 4004 0 -1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_194
timestamp 1693479267
transform 1 0 3956 0 1 3105
box -2 -3 98 103
use FILL  FILL_30_7_0
timestamp 1693479267
transform 1 0 4100 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_7_1
timestamp 1693479267
transform 1 0 4108 0 -1 3105
box -2 -3 10 103
use OAI21X1  OAI21X1_955
timestamp 1693479267
transform 1 0 4116 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_960
timestamp 1693479267
transform -1 0 4084 0 1 3105
box -2 -3 34 103
use FILL  FILL_31_7_0
timestamp 1693479267
transform 1 0 4084 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_7_1
timestamp 1693479267
transform 1 0 4092 0 1 3105
box -2 -3 10 103
use CLKBUF1  CLKBUF1_22
timestamp 1693479267
transform 1 0 4100 0 1 3105
box -2 -3 74 103
use OAI21X1  OAI21X1_954
timestamp 1693479267
transform -1 0 4180 0 -1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_215
timestamp 1693479267
transform 1 0 4180 0 -1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_195
timestamp 1693479267
transform 1 0 4172 0 1 3105
box -2 -3 98 103
use INVX1  INVX1_720
timestamp 1693479267
transform 1 0 4276 0 -1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_956
timestamp 1693479267
transform 1 0 4292 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_957
timestamp 1693479267
transform -1 0 4356 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_962
timestamp 1693479267
transform 1 0 4268 0 1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_199
timestamp 1693479267
transform 1 0 4300 0 1 3105
box -2 -3 98 103
use OAI21X1  OAI21X1_963
timestamp 1693479267
transform 1 0 4356 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_1024
timestamp 1693479267
transform 1 0 4388 0 -1 3105
box -2 -3 26 103
use BUFX2  BUFX2_78
timestamp 1693479267
transform -1 0 4436 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_1003
timestamp 1693479267
transform 1 0 4436 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_1025
timestamp 1693479267
transform 1 0 4396 0 1 3105
box -2 -3 26 103
use NAND3X1  NAND3X1_360
timestamp 1693479267
transform 1 0 4420 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_1004
timestamp 1693479267
transform 1 0 4460 0 -1 3105
box -2 -3 26 103
use INVX1  INVX1_727
timestamp 1693479267
transform 1 0 4484 0 -1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_969
timestamp 1693479267
transform 1 0 4500 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_972
timestamp 1693479267
transform 1 0 4532 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_974
timestamp 1693479267
transform 1 0 4452 0 1 3105
box -2 -3 34 103
use BUFX4  BUFX4_116
timestamp 1693479267
transform -1 0 4516 0 1 3105
box -2 -3 34 103
use BUFX2  BUFX2_82
timestamp 1693479267
transform -1 0 4540 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_1007
timestamp 1693479267
transform 1 0 4540 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_1005
timestamp 1693479267
transform 1 0 4564 0 -1 3105
box -2 -3 26 103
use FILL  FILL_31_1
timestamp 1693479267
transform -1 0 4596 0 -1 3105
box -2 -3 10 103
use FILL  FILL_31_2
timestamp 1693479267
transform -1 0 4604 0 -1 3105
box -2 -3 10 103
use NAND2X1  NAND2X1_1006
timestamp 1693479267
transform 1 0 4564 0 1 3105
box -2 -3 26 103
use FILL  FILL_32_1
timestamp 1693479267
transform 1 0 4588 0 1 3105
box -2 -3 10 103
use FILL  FILL_32_2
timestamp 1693479267
transform 1 0 4596 0 1 3105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_408
timestamp 1693479267
transform 1 0 4 0 -1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_412
timestamp 1693479267
transform 1 0 100 0 -1 3305
box -2 -3 98 103
use INVX1  INVX1_228
timestamp 1693479267
transform 1 0 196 0 -1 3305
box -2 -3 18 103
use NOR2X1  NOR2X1_19
timestamp 1693479267
transform -1 0 236 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_111
timestamp 1693479267
transform -1 0 260 0 -1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_15
timestamp 1693479267
transform 1 0 260 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_109
timestamp 1693479267
transform -1 0 308 0 -1 3305
box -2 -3 26 103
use AOI22X1  AOI22X1_41
timestamp 1693479267
transform 1 0 308 0 -1 3305
box -2 -3 42 103
use OAI21X1  OAI21X1_226
timestamp 1693479267
transform 1 0 348 0 -1 3305
box -2 -3 34 103
use INVX2  INVX2_4
timestamp 1693479267
transform 1 0 380 0 -1 3305
box -2 -3 18 103
use NOR2X1  NOR2X1_20
timestamp 1693479267
transform 1 0 396 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_112
timestamp 1693479267
transform -1 0 444 0 -1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_17
timestamp 1693479267
transform -1 0 468 0 -1 3305
box -2 -3 26 103
use OR2X2  OR2X2_6
timestamp 1693479267
transform 1 0 468 0 -1 3305
box -2 -3 34 103
use FILL  FILL_32_0_0
timestamp 1693479267
transform 1 0 500 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_0_1
timestamp 1693479267
transform 1 0 508 0 -1 3305
box -2 -3 10 103
use INVX1  INVX1_229
timestamp 1693479267
transform 1 0 516 0 -1 3305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_290
timestamp 1693479267
transform 1 0 532 0 -1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_306
timestamp 1693479267
transform 1 0 628 0 -1 3305
box -2 -3 98 103
use INVX1  INVX1_138
timestamp 1693479267
transform 1 0 724 0 -1 3305
box -2 -3 18 103
use NAND3X1  NAND3X1_4
timestamp 1693479267
transform 1 0 740 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_6
timestamp 1693479267
transform 1 0 772 0 -1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_886
timestamp 1693479267
transform -1 0 828 0 -1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_318
timestamp 1693479267
transform 1 0 828 0 -1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_123
timestamp 1693479267
transform 1 0 924 0 -1 3305
box -2 -3 98 103
use FILL  FILL_32_1_0
timestamp 1693479267
transform 1 0 1020 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_1_1
timestamp 1693479267
transform 1 0 1028 0 -1 3305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_22
timestamp 1693479267
transform 1 0 1036 0 -1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_34
timestamp 1693479267
transform 1 0 1132 0 -1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_69
timestamp 1693479267
transform 1 0 1228 0 -1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_71
timestamp 1693479267
transform 1 0 1324 0 -1 3305
box -2 -3 98 103
use INVX1  INVX1_124
timestamp 1693479267
transform 1 0 1420 0 -1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_206
timestamp 1693479267
transform 1 0 1436 0 -1 3305
box -2 -3 34 103
use INVX1  INVX1_204
timestamp 1693479267
transform -1 0 1484 0 -1 3305
box -2 -3 18 103
use INVX1  INVX1_122
timestamp 1693479267
transform 1 0 1484 0 -1 3305
box -2 -3 18 103
use FILL  FILL_32_2_0
timestamp 1693479267
transform -1 0 1508 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_2_1
timestamp 1693479267
transform -1 0 1516 0 -1 3305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_91
timestamp 1693479267
transform -1 0 1612 0 -1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_59
timestamp 1693479267
transform -1 0 1708 0 -1 3305
box -2 -3 98 103
use INVX1  INVX1_214
timestamp 1693479267
transform -1 0 1724 0 -1 3305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_101
timestamp 1693479267
transform -1 0 1820 0 -1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_228
timestamp 1693479267
transform -1 0 1916 0 -1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_144
timestamp 1693479267
transform 1 0 1916 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_143
timestamp 1693479267
transform -1 0 1980 0 -1 3305
box -2 -3 34 103
use BUFX4  BUFX4_273
timestamp 1693479267
transform -1 0 2012 0 -1 3305
box -2 -3 34 103
use FILL  FILL_32_3_0
timestamp 1693479267
transform -1 0 2020 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_3_1
timestamp 1693479267
transform -1 0 2028 0 -1 3305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_248
timestamp 1693479267
transform -1 0 2124 0 -1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_236
timestamp 1693479267
transform -1 0 2220 0 -1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_123
timestamp 1693479267
transform 1 0 2220 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_148
timestamp 1693479267
transform 1 0 2252 0 -1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_253
timestamp 1693479267
transform -1 0 2380 0 -1 3305
box -2 -3 98 103
use NAND2X1  NAND2X1_775
timestamp 1693479267
transform -1 0 2404 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_86
timestamp 1693479267
transform 1 0 2404 0 -1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_84
timestamp 1693479267
transform 1 0 2428 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_766
timestamp 1693479267
transform -1 0 2484 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_876
timestamp 1693479267
transform 1 0 2484 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_885
timestamp 1693479267
transform 1 0 2508 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_834
timestamp 1693479267
transform -1 0 2556 0 -1 3305
box -2 -3 26 103
use FILL  FILL_32_4_0
timestamp 1693479267
transform 1 0 2556 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_4_1
timestamp 1693479267
transform 1 0 2564 0 -1 3305
box -2 -3 10 103
use INVX1  INVX1_71
timestamp 1693479267
transform 1 0 2572 0 -1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_70
timestamp 1693479267
transform 1 0 2588 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_891
timestamp 1693479267
transform 1 0 2620 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_724
timestamp 1693479267
transform 1 0 2644 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_888
timestamp 1693479267
transform 1 0 2668 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_787
timestamp 1693479267
transform -1 0 2716 0 -1 3305
box -2 -3 26 103
use BUFX4  BUFX4_133
timestamp 1693479267
transform -1 0 2748 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_897
timestamp 1693479267
transform 1 0 2748 0 -1 3305
box -2 -3 26 103
use BUFX4  BUFX4_63
timestamp 1693479267
transform -1 0 2804 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_861
timestamp 1693479267
transform 1 0 2804 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_831
timestamp 1693479267
transform 1 0 2828 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_754
timestamp 1693479267
transform -1 0 2876 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_867
timestamp 1693479267
transform 1 0 2876 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_864
timestamp 1693479267
transform -1 0 2924 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_727
timestamp 1693479267
transform -1 0 2948 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_733
timestamp 1693479267
transform -1 0 2972 0 -1 3305
box -2 -3 26 103
use INVX1  INVX1_67
timestamp 1693479267
transform 1 0 2972 0 -1 3305
box -2 -3 18 103
use NAND2X1  NAND2X1_837
timestamp 1693479267
transform 1 0 2988 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_843
timestamp 1693479267
transform 1 0 3012 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_712
timestamp 1693479267
transform -1 0 3060 0 -1 3305
box -2 -3 26 103
use FILL  FILL_32_5_0
timestamp 1693479267
transform 1 0 3060 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_5_1
timestamp 1693479267
transform 1 0 3068 0 -1 3305
box -2 -3 10 103
use OAI21X1  OAI21X1_66
timestamp 1693479267
transform 1 0 3076 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_822
timestamp 1693479267
transform 1 0 3108 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_802
timestamp 1693479267
transform -1 0 3156 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_98
timestamp 1693479267
transform 1 0 3156 0 -1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_96
timestamp 1693479267
transform -1 0 3212 0 -1 3305
box -2 -3 34 103
use INVX1  INVX1_97
timestamp 1693479267
transform -1 0 3228 0 -1 3305
box -2 -3 18 103
use NAND2X1  NAND2X1_796
timestamp 1693479267
transform -1 0 3252 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_742
timestamp 1693479267
transform -1 0 3276 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_852
timestamp 1693479267
transform 1 0 3276 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_912
timestamp 1693479267
transform 1 0 3300 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_906
timestamp 1693479267
transform -1 0 3348 0 -1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_94
timestamp 1693479267
transform -1 0 3380 0 -1 3305
box -2 -3 34 103
use INVX1  INVX1_95
timestamp 1693479267
transform -1 0 3396 0 -1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_33
timestamp 1693479267
transform -1 0 3428 0 -1 3305
box -2 -3 34 103
use INVX1  INVX1_33
timestamp 1693479267
transform -1 0 3444 0 -1 3305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_376
timestamp 1693479267
transform -1 0 3540 0 -1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_49
timestamp 1693479267
transform -1 0 3572 0 -1 3305
box -2 -3 34 103
use FILL  FILL_32_6_0
timestamp 1693479267
transform -1 0 3580 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_6_1
timestamp 1693479267
transform -1 0 3588 0 -1 3305
box -2 -3 10 103
use INVX1  INVX1_49
timestamp 1693479267
transform -1 0 3604 0 -1 3305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_398
timestamp 1693479267
transform -1 0 3700 0 -1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_55
timestamp 1693479267
transform -1 0 3732 0 -1 3305
box -2 -3 34 103
use INVX1  INVX1_55
timestamp 1693479267
transform -1 0 3748 0 -1 3305
box -2 -3 18 103
use NAND2X1  NAND2X1_38
timestamp 1693479267
transform -1 0 3772 0 -1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_212
timestamp 1693479267
transform 1 0 3772 0 -1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_210
timestamp 1693479267
transform 1 0 3868 0 -1 3305
box -2 -3 98 103
use INVX1  INVX1_722
timestamp 1693479267
transform 1 0 3964 0 -1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_961
timestamp 1693479267
transform 1 0 3980 0 -1 3305
box -2 -3 34 103
use INVX1  INVX1_724
timestamp 1693479267
transform 1 0 4012 0 -1 3305
box -2 -3 18 103
use CLKBUF1  CLKBUF1_8
timestamp 1693479267
transform -1 0 4100 0 -1 3305
box -2 -3 74 103
use FILL  FILL_32_7_0
timestamp 1693479267
transform 1 0 4100 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_7_1
timestamp 1693479267
transform 1 0 4108 0 -1 3305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_219
timestamp 1693479267
transform 1 0 4116 0 -1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_965
timestamp 1693479267
transform 1 0 4212 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_964
timestamp 1693479267
transform 1 0 4244 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_1054
timestamp 1693479267
transform 1 0 4276 0 -1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_203
timestamp 1693479267
transform 1 0 4308 0 -1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_206
timestamp 1693479267
transform 1 0 4404 0 -1 3305
box -2 -3 98 103
use BUFX4  BUFX4_252
timestamp 1693479267
transform -1 0 4532 0 -1 3305
box -2 -3 34 103
use INVX1  INVX1_731
timestamp 1693479267
transform 1 0 4532 0 -1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_973
timestamp 1693479267
transform 1 0 4548 0 -1 3305
box -2 -3 34 103
use FILL  FILL_33_1
timestamp 1693479267
transform -1 0 4588 0 -1 3305
box -2 -3 10 103
use FILL  FILL_33_2
timestamp 1693479267
transform -1 0 4596 0 -1 3305
box -2 -3 10 103
use FILL  FILL_33_3
timestamp 1693479267
transform -1 0 4604 0 -1 3305
box -2 -3 10 103
use INVX1  INVX1_162
timestamp 1693479267
transform 1 0 4 0 1 3305
box -2 -3 18 103
use NOR3X1  NOR3X1_21
timestamp 1693479267
transform -1 0 84 0 1 3305
box -2 -3 66 103
use DFFPOSX1  DFFPOSX1_414
timestamp 1693479267
transform 1 0 84 0 1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_413
timestamp 1693479267
transform 1 0 180 0 1 3305
box -2 -3 98 103
use BUFX2  BUFX2_88
timestamp 1693479267
transform -1 0 300 0 1 3305
box -2 -3 26 103
use INVX1  INVX1_155
timestamp 1693479267
transform 1 0 300 0 1 3305
box -2 -3 18 103
use INVX1  INVX1_154
timestamp 1693479267
transform 1 0 316 0 1 3305
box -2 -3 18 103
use NOR3X1  NOR3X1_14
timestamp 1693479267
transform -1 0 396 0 1 3305
box -2 -3 66 103
use INVX1  INVX1_225
timestamp 1693479267
transform 1 0 396 0 1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_225
timestamp 1693479267
transform 1 0 412 0 1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_291
timestamp 1693479267
transform 1 0 444 0 1 3305
box -2 -3 98 103
use FILL  FILL_33_0_0
timestamp 1693479267
transform -1 0 548 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_0_1
timestamp 1693479267
transform -1 0 556 0 1 3305
box -2 -3 10 103
use OAI21X1  OAI21X1_880
timestamp 1693479267
transform -1 0 588 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_647
timestamp 1693479267
transform -1 0 604 0 1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_879
timestamp 1693479267
transform -1 0 636 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_646
timestamp 1693479267
transform -1 0 652 0 1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_878
timestamp 1693479267
transform -1 0 684 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_645
timestamp 1693479267
transform -1 0 700 0 1 3305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_307
timestamp 1693479267
transform 1 0 700 0 1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_322
timestamp 1693479267
transform 1 0 796 0 1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_139
timestamp 1693479267
transform 1 0 892 0 1 3305
box -2 -3 98 103
use FILL  FILL_33_1_0
timestamp 1693479267
transform 1 0 988 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_1_1
timestamp 1693479267
transform 1 0 996 0 1 3305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_27
timestamp 1693479267
transform 1 0 1004 0 1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_124
timestamp 1693479267
transform 1 0 1100 0 1 3305
box -2 -3 98 103
use AOI22X1  AOI22X1_14
timestamp 1693479267
transform 1 0 1196 0 1 3305
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_12
timestamp 1693479267
transform 1 0 1236 0 1 3305
box -2 -3 98 103
use OAI21X1  OAI21X1_199
timestamp 1693479267
transform -1 0 1364 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_197
timestamp 1693479267
transform -1 0 1380 0 1 3305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_84
timestamp 1693479267
transform -1 0 1476 0 1 3305
box -2 -3 98 103
use BUFX4  BUFX4_145
timestamp 1693479267
transform 1 0 1476 0 1 3305
box -2 -3 34 103
use FILL  FILL_33_2_0
timestamp 1693479267
transform -1 0 1516 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_2_1
timestamp 1693479267
transform -1 0 1524 0 1 3305
box -2 -3 10 103
use AOI22X1  AOI22X1_12
timestamp 1693479267
transform -1 0 1564 0 1 3305
box -2 -3 42 103
use AOI22X1  AOI22X1_22
timestamp 1693479267
transform -1 0 1604 0 1 3305
box -2 -3 42 103
use BUFX4  BUFX4_237
timestamp 1693479267
transform -1 0 1636 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_197
timestamp 1693479267
transform -1 0 1668 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_207
timestamp 1693479267
transform -1 0 1700 0 1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_70
timestamp 1693479267
transform -1 0 1796 0 1 3305
box -2 -3 98 103
use INVX1  INVX1_195
timestamp 1693479267
transform -1 0 1812 0 1 3305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_82
timestamp 1693479267
transform -1 0 1908 0 1 3305
box -2 -3 98 103
use INVX1  INVX1_205
timestamp 1693479267
transform -1 0 1924 0 1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_109
timestamp 1693479267
transform -1 0 1956 0 1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_92
timestamp 1693479267
transform -1 0 2052 0 1 3305
box -2 -3 98 103
use FILL  FILL_33_3_0
timestamp 1693479267
transform -1 0 2060 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_3_1
timestamp 1693479267
transform -1 0 2068 0 1 3305
box -2 -3 10 103
use OAI21X1  OAI21X1_125
timestamp 1693479267
transform -1 0 2100 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_145
timestamp 1693479267
transform -1 0 2132 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_123
timestamp 1693479267
transform 1 0 2132 0 1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_146
timestamp 1693479267
transform -1 0 2180 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_105
timestamp 1693479267
transform 1 0 2180 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_112
timestamp 1693479267
transform 1 0 2212 0 1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_124
timestamp 1693479267
transform 1 0 2228 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_777
timestamp 1693479267
transform -1 0 2284 0 1 3305
box -2 -3 26 103
use BUFX4  BUFX4_193
timestamp 1693479267
transform -1 0 2316 0 1 3305
box -2 -3 34 103
use BUFX4  BUFX4_195
timestamp 1693479267
transform -1 0 2348 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_508
timestamp 1693479267
transform 1 0 2348 0 1 3305
box -2 -3 18 103
use NAND2X1  NAND2X1_768
timestamp 1693479267
transform -1 0 2388 0 1 3305
box -2 -3 26 103
use CLKBUF1  CLKBUF1_23
timestamp 1693479267
transform -1 0 2460 0 1 3305
box -2 -3 74 103
use INVX1  INVX1_581
timestamp 1693479267
transform 1 0 2460 0 1 3305
box -2 -3 18 103
use BUFX4  BUFX4_158
timestamp 1693479267
transform -1 0 2508 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_887
timestamp 1693479267
transform -1 0 2532 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_836
timestamp 1693479267
transform 1 0 2532 0 1 3305
box -2 -3 26 103
use FILL  FILL_33_4_0
timestamp 1693479267
transform 1 0 2556 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_4_1
timestamp 1693479267
transform 1 0 2564 0 1 3305
box -2 -3 10 103
use NAND2X1  NAND2X1_72
timestamp 1693479267
transform 1 0 2572 0 1 3305
box -2 -3 26 103
use NAND3X1  NAND3X1_264
timestamp 1693479267
transform 1 0 2596 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_726
timestamp 1693479267
transform -1 0 2652 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_890
timestamp 1693479267
transform -1 0 2676 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_789
timestamp 1693479267
transform -1 0 2700 0 1 3305
box -2 -3 26 103
use INVX1  INVX1_534
timestamp 1693479267
transform -1 0 2716 0 1 3305
box -2 -3 18 103
use INVX1  INVX1_607
timestamp 1693479267
transform 1 0 2716 0 1 3305
box -2 -3 18 103
use NAND3X1  NAND3X1_290
timestamp 1693479267
transform 1 0 2732 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_899
timestamp 1693479267
transform 1 0 2764 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_756
timestamp 1693479267
transform -1 0 2812 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_863
timestamp 1693479267
transform 1 0 2812 0 1 3305
box -2 -3 26 103
use NAND3X1  NAND3X1_260
timestamp 1693479267
transform -1 0 2868 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_576
timestamp 1693479267
transform -1 0 2884 0 1 3305
box -2 -3 18 103
use NAND2X1  NAND2X1_729
timestamp 1693479267
transform -1 0 2908 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_833
timestamp 1693479267
transform 1 0 2908 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_735
timestamp 1693479267
transform -1 0 2956 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_866
timestamp 1693479267
transform 1 0 2956 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_869
timestamp 1693479267
transform 1 0 2980 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_714
timestamp 1693479267
transform -1 0 3028 0 1 3305
box -2 -3 26 103
use INVX1  INVX1_503
timestamp 1693479267
transform 1 0 3028 0 1 3305
box -2 -3 18 103
use FILL  FILL_33_5_0
timestamp 1693479267
transform 1 0 3044 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_5_1
timestamp 1693479267
transform 1 0 3052 0 1 3305
box -2 -3 10 103
use BUFX4  BUFX4_156
timestamp 1693479267
transform 1 0 3060 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_68
timestamp 1693479267
transform 1 0 3092 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_804
timestamp 1693479267
transform -1 0 3140 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_824
timestamp 1693479267
transform 1 0 3140 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_798
timestamp 1693479267
transform -1 0 3188 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_795
timestamp 1693479267
transform -1 0 3212 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_793
timestamp 1693479267
transform -1 0 3236 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_744
timestamp 1693479267
transform -1 0 3260 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_860
timestamp 1693479267
transform 1 0 3260 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_854
timestamp 1693479267
transform 1 0 3284 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_908
timestamp 1693479267
transform -1 0 3332 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_821
timestamp 1693479267
transform 1 0 3332 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_37
timestamp 1693479267
transform -1 0 3380 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_33
timestamp 1693479267
transform 1 0 3380 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_96
timestamp 1693479267
transform -1 0 3428 0 1 3305
box -2 -3 26 103
use BUFX4  BUFX4_28
timestamp 1693479267
transform -1 0 3460 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_48
timestamp 1693479267
transform -1 0 3484 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_59
timestamp 1693479267
transform -1 0 3508 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_55
timestamp 1693479267
transform -1 0 3532 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_49
timestamp 1693479267
transform -1 0 3556 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_62
timestamp 1693479267
transform -1 0 3580 0 1 3305
box -2 -3 26 103
use FILL  FILL_33_6_0
timestamp 1693479267
transform 1 0 3580 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_6_1
timestamp 1693479267
transform 1 0 3588 0 1 3305
box -2 -3 10 103
use INVX1  INVX1_61
timestamp 1693479267
transform 1 0 3596 0 1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_61
timestamp 1693479267
transform 1 0 3612 0 1 3305
box -2 -3 34 103
use BUFX4  BUFX4_25
timestamp 1693479267
transform -1 0 3676 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_48
timestamp 1693479267
transform -1 0 3708 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_48
timestamp 1693479267
transform -1 0 3724 0 1 3305
box -2 -3 18 103
use NAND2X1  NAND2X1_46
timestamp 1693479267
transform 1 0 3724 0 1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_391
timestamp 1693479267
transform 1 0 3748 0 1 3305
box -2 -3 98 103
use INVX1  INVX1_46
timestamp 1693479267
transform 1 0 3844 0 1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_46
timestamp 1693479267
transform 1 0 3860 0 1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_389
timestamp 1693479267
transform 1 0 3892 0 1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_193
timestamp 1693479267
transform 1 0 3988 0 1 3305
box -2 -3 98 103
use FILL  FILL_33_7_0
timestamp 1693479267
transform 1 0 4084 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_7_1
timestamp 1693479267
transform 1 0 4092 0 1 3305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_205
timestamp 1693479267
transform 1 0 4100 0 1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_196
timestamp 1693479267
transform 1 0 4196 0 1 3305
box -2 -3 98 103
use AOI22X1  AOI22X1_169
timestamp 1693479267
transform -1 0 4332 0 1 3305
box -2 -3 42 103
use OAI21X1  OAI21X1_1053
timestamp 1693479267
transform -1 0 4364 0 1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_190
timestamp 1693479267
transform 1 0 4364 0 1 3305
box -2 -3 98 103
use BUFX2  BUFX2_83
timestamp 1693479267
transform -1 0 4484 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_1009
timestamp 1693479267
transform 1 0 4484 0 1 3305
box -2 -3 26 103
use BUFX2  BUFX2_77
timestamp 1693479267
transform -1 0 4532 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_1008
timestamp 1693479267
transform 1 0 4532 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_1002
timestamp 1693479267
transform 1 0 4556 0 1 3305
box -2 -3 26 103
use FILL  FILL_34_1
timestamp 1693479267
transform 1 0 4580 0 1 3305
box -2 -3 10 103
use FILL  FILL_34_2
timestamp 1693479267
transform 1 0 4588 0 1 3305
box -2 -3 10 103
use FILL  FILL_34_3
timestamp 1693479267
transform 1 0 4596 0 1 3305
box -2 -3 10 103
use INVX1  INVX1_161
timestamp 1693479267
transform 1 0 4 0 -1 3505
box -2 -3 18 103
use NOR3X1  NOR3X1_20
timestamp 1693479267
transform -1 0 84 0 -1 3505
box -2 -3 66 103
use NOR3X1  NOR3X1_26
timestamp 1693479267
transform -1 0 148 0 -1 3505
box -2 -3 66 103
use BUFX4  BUFX4_48
timestamp 1693479267
transform -1 0 180 0 -1 3505
box -2 -3 34 103
use BUFX4  BUFX4_244
timestamp 1693479267
transform -1 0 212 0 -1 3505
box -2 -3 34 103
use BUFX4  BUFX4_242
timestamp 1693479267
transform 1 0 212 0 -1 3505
box -2 -3 34 103
use BUFX4  BUFX4_46
timestamp 1693479267
transform 1 0 244 0 -1 3505
box -2 -3 34 103
use NOR3X1  NOR3X1_15
timestamp 1693479267
transform -1 0 340 0 -1 3505
box -2 -3 66 103
use NOR3X1  NOR3X1_8
timestamp 1693479267
transform -1 0 404 0 -1 3505
box -2 -3 66 103
use INVX1  INVX1_145
timestamp 1693479267
transform -1 0 420 0 -1 3505
box -2 -3 18 103
use NAND2X1  NAND2X1_924
timestamp 1693479267
transform 1 0 420 0 -1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_921
timestamp 1693479267
transform 1 0 444 0 -1 3505
box -2 -3 26 103
use INVX1  INVX1_644
timestamp 1693479267
transform 1 0 468 0 -1 3505
box -2 -3 18 103
use FILL  FILL_34_0_0
timestamp 1693479267
transform -1 0 492 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_0_1
timestamp 1693479267
transform -1 0 500 0 -1 3505
box -2 -3 10 103
use OAI21X1  OAI21X1_877
timestamp 1693479267
transform -1 0 532 0 -1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_343
timestamp 1693479267
transform 1 0 532 0 -1 3505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_304
timestamp 1693479267
transform 1 0 628 0 -1 3505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_321
timestamp 1693479267
transform 1 0 724 0 -1 3505
box -2 -3 98 103
use INVX1  INVX1_657
timestamp 1693479267
transform -1 0 836 0 -1 3505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_138
timestamp 1693479267
transform 1 0 836 0 -1 3505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_26
timestamp 1693479267
transform 1 0 932 0 -1 3505
box -2 -3 98 103
use FILL  FILL_34_1_0
timestamp 1693479267
transform 1 0 1028 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_1_1
timestamp 1693479267
transform 1 0 1036 0 -1 3505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_11
timestamp 1693479267
transform 1 0 1044 0 -1 3505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_52
timestamp 1693479267
transform -1 0 1236 0 -1 3505
box -2 -3 98 103
use AOI22X1  AOI22X1_27
timestamp 1693479267
transform -1 0 1276 0 -1 3505
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_65
timestamp 1693479267
transform -1 0 1372 0 -1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_212
timestamp 1693479267
transform -1 0 1404 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_210
timestamp 1693479267
transform -1 0 1420 0 -1 3505
box -2 -3 18 103
use AOI22X1  AOI22X1_35
timestamp 1693479267
transform -1 0 1460 0 -1 3505
box -2 -3 42 103
use OAI21X1  OAI21X1_220
timestamp 1693479267
transform -1 0 1492 0 -1 3505
box -2 -3 34 103
use FILL  FILL_34_2_0
timestamp 1693479267
transform -1 0 1500 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_2_1
timestamp 1693479267
transform -1 0 1508 0 -1 3505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_97
timestamp 1693479267
transform -1 0 1604 0 -1 3505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_50
timestamp 1693479267
transform -1 0 1700 0 -1 3505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_60
timestamp 1693479267
transform -1 0 1796 0 -1 3505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_251
timestamp 1693479267
transform -1 0 1892 0 -1 3505
box -2 -3 98 103
use INVX1  INVX1_113
timestamp 1693479267
transform 1 0 1892 0 -1 3505
box -2 -3 18 103
use OAI21X1  OAI21X1_111
timestamp 1693479267
transform -1 0 1940 0 -1 3505
box -2 -3 34 103
use BUFX4  BUFX4_192
timestamp 1693479267
transform 1 0 1940 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_135
timestamp 1693479267
transform -1 0 2004 0 -1 3505
box -2 -3 34 103
use BUFX4  BUFX4_182
timestamp 1693479267
transform 1 0 2004 0 -1 3505
box -2 -3 34 103
use FILL  FILL_34_3_0
timestamp 1693479267
transform 1 0 2036 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_3_1
timestamp 1693479267
transform 1 0 2044 0 -1 3505
box -2 -3 10 103
use OAI21X1  OAI21X1_126
timestamp 1693479267
transform 1 0 2052 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_103
timestamp 1693479267
transform 1 0 2084 0 -1 3505
box -2 -3 18 103
use BUFX4  BUFX4_183
timestamp 1693479267
transform 1 0 2100 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_86
timestamp 1693479267
transform 1 0 2132 0 -1 3505
box -2 -3 18 103
use OAI21X1  OAI21X1_106
timestamp 1693479267
transform 1 0 2148 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_550
timestamp 1693479267
transform 1 0 2180 0 -1 3505
box -2 -3 18 103
use INVX1  INVX1_623
timestamp 1693479267
transform 1 0 2196 0 -1 3505
box -2 -3 18 103
use NAND3X1  NAND3X1_236
timestamp 1693479267
transform 1 0 2212 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_237
timestamp 1693479267
transform 1 0 2244 0 -1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_87
timestamp 1693479267
transform 1 0 2276 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_85
timestamp 1693479267
transform 1 0 2300 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_194
timestamp 1693479267
transform -1 0 2364 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_195
timestamp 1693479267
transform 1 0 2364 0 -1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_718
timestamp 1693479267
transform 1 0 2396 0 -1 3505
box -2 -3 26 103
use INVX1  INVX1_84
timestamp 1693479267
transform 1 0 2420 0 -1 3505
box -2 -3 18 103
use NAND2X1  NAND2X1_85
timestamp 1693479267
transform 1 0 2436 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_83
timestamp 1693479267
transform 1 0 2460 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_306
timestamp 1693479267
transform 1 0 2492 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_627
timestamp 1693479267
transform 1 0 2524 0 -1 3505
box -2 -3 18 103
use FILL  FILL_34_4_0
timestamp 1693479267
transform 1 0 2540 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_4_1
timestamp 1693479267
transform 1 0 2548 0 -1 3505
box -2 -3 10 103
use NAND3X1  NAND3X1_310
timestamp 1693479267
transform 1 0 2556 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_307
timestamp 1693479267
transform -1 0 2620 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_554
timestamp 1693479267
transform 1 0 2620 0 -1 3505
box -2 -3 18 103
use NAND3X1  NAND3X1_265
timestamp 1693479267
transform -1 0 2668 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_221
timestamp 1693479267
transform -1 0 2700 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_220
timestamp 1693479267
transform 1 0 2700 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_291
timestamp 1693479267
transform 1 0 2732 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_311
timestamp 1693479267
transform -1 0 2796 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_240
timestamp 1693479267
transform 1 0 2796 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_241
timestamp 1693479267
transform 1 0 2828 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_520
timestamp 1693479267
transform 1 0 2860 0 -1 3505
box -2 -3 18 103
use INVX1  INVX1_564
timestamp 1693479267
transform 1 0 2876 0 -1 3505
box -2 -3 18 103
use NAND3X1  NAND3X1_217
timestamp 1693479267
transform 1 0 2892 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_207
timestamp 1693479267
transform 1 0 2924 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_206
timestamp 1693479267
transform 1 0 2956 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_250
timestamp 1693479267
transform 1 0 2988 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_190
timestamp 1693479267
transform -1 0 3052 0 -1 3505
box -2 -3 34 103
use FILL  FILL_34_5_0
timestamp 1693479267
transform 1 0 3052 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_5_1
timestamp 1693479267
transform 1 0 3060 0 -1 3505
box -2 -3 10 103
use NAND2X1  NAND2X1_845
timestamp 1693479267
transform 1 0 3068 0 -1 3505
box -2 -3 26 103
use NAND3X1  NAND3X1_191
timestamp 1693479267
transform 1 0 3092 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_251
timestamp 1693479267
transform 1 0 3124 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_245
timestamp 1693479267
transform 1 0 3156 0 -1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_800
timestamp 1693479267
transform -1 0 3212 0 -1 3505
box -2 -3 26 103
use NAND3X1  NAND3X1_321
timestamp 1693479267
transform 1 0 3212 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_636
timestamp 1693479267
transform -1 0 3260 0 -1 3505
box -2 -3 18 103
use INVX1  INVX1_563
timestamp 1693479267
transform 1 0 3260 0 -1 3505
box -2 -3 18 103
use NAND3X1  NAND3X1_287
timestamp 1693479267
transform 1 0 3276 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_315
timestamp 1693479267
transform -1 0 3340 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_261
timestamp 1693479267
transform 1 0 3340 0 -1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_828
timestamp 1693479267
transform 1 0 3372 0 -1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_846
timestamp 1693479267
transform 1 0 3396 0 -1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_903
timestamp 1693479267
transform -1 0 3444 0 -1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_95
timestamp 1693479267
transform 1 0 3444 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_93
timestamp 1693479267
transform -1 0 3500 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_94
timestamp 1693479267
transform -1 0 3516 0 -1 3505
box -2 -3 18 103
use NAND2X1  NAND2X1_56
timestamp 1693479267
transform 1 0 3516 0 -1 3505
box -2 -3 26 103
use INVX1  INVX1_56
timestamp 1693479267
transform -1 0 3556 0 -1 3505
box -2 -3 18 103
use FILL  FILL_34_6_0
timestamp 1693479267
transform 1 0 3556 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_6_1
timestamp 1693479267
transform 1 0 3564 0 -1 3505
box -2 -3 10 103
use OAI21X1  OAI21X1_56
timestamp 1693479267
transform 1 0 3572 0 -1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_61
timestamp 1693479267
transform -1 0 3628 0 -1 3505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_399
timestamp 1693479267
transform 1 0 3628 0 -1 3505
box -2 -3 98 103
use NAND2X1  NAND2X1_64
timestamp 1693479267
transform -1 0 3748 0 -1 3505
box -2 -3 26 103
use INVX1  INVX1_64
timestamp 1693479267
transform 1 0 3748 0 -1 3505
box -2 -3 18 103
use OAI21X1  OAI21X1_64
timestamp 1693479267
transform 1 0 3764 0 -1 3505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_29
timestamp 1693479267
transform -1 0 3868 0 -1 3505
box -2 -3 74 103
use OAI21X1  OAI21X1_42
timestamp 1693479267
transform -1 0 3900 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_42
timestamp 1693479267
transform -1 0 3916 0 -1 3505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_407
timestamp 1693479267
transform 1 0 3916 0 -1 3505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_385
timestamp 1693479267
transform 1 0 4012 0 -1 3505
box -2 -3 98 103
use FILL  FILL_34_7_0
timestamp 1693479267
transform 1 0 4108 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_7_1
timestamp 1693479267
transform 1 0 4116 0 -1 3505
box -2 -3 10 103
use CLKBUF1  CLKBUF1_16
timestamp 1693479267
transform 1 0 4124 0 -1 3505
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_221
timestamp 1693479267
transform 1 0 4196 0 -1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_966
timestamp 1693479267
transform 1 0 4292 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_1055
timestamp 1693479267
transform 1 0 4324 0 -1 3505
box -2 -3 34 103
use AOI22X1  AOI22X1_171
timestamp 1693479267
transform -1 0 4396 0 -1 3505
box -2 -3 42 103
use INVX1  INVX1_733
timestamp 1693479267
transform 1 0 4396 0 -1 3505
box -2 -3 18 103
use NOR2X1  NOR2X1_479
timestamp 1693479267
transform 1 0 4412 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_968
timestamp 1693479267
transform -1 0 4468 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_726
timestamp 1693479267
transform -1 0 4484 0 -1 3505
box -2 -3 18 103
use NAND2X1  NAND2X1_1023
timestamp 1693479267
transform 1 0 4484 0 -1 3505
box -2 -3 26 103
use NAND3X1  NAND3X1_359
timestamp 1693479267
transform 1 0 4508 0 -1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_1021
timestamp 1693479267
transform -1 0 4564 0 -1 3505
box -2 -3 26 103
use INVX1  INVX1_718
timestamp 1693479267
transform 1 0 4564 0 -1 3505
box -2 -3 18 103
use FILL  FILL_35_1
timestamp 1693479267
transform -1 0 4588 0 -1 3505
box -2 -3 10 103
use FILL  FILL_35_2
timestamp 1693479267
transform -1 0 4596 0 -1 3505
box -2 -3 10 103
use FILL  FILL_35_3
timestamp 1693479267
transform -1 0 4604 0 -1 3505
box -2 -3 10 103
use INVX1  INVX1_165
timestamp 1693479267
transform 1 0 4 0 1 3505
box -2 -3 18 103
use INVX1  INVX1_167
timestamp 1693479267
transform 1 0 20 0 1 3505
box -2 -3 18 103
use NOR3X1  NOR3X1_24
timestamp 1693479267
transform -1 0 100 0 1 3505
box -2 -3 66 103
use DFFPOSX1  DFFPOSX1_417
timestamp 1693479267
transform 1 0 100 0 1 3505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_419
timestamp 1693479267
transform 1 0 196 0 1 3505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_342
timestamp 1693479267
transform 1 0 292 0 1 3505
box -2 -3 98 103
use NOR2X1  NOR2X1_22
timestamp 1693479267
transform 1 0 388 0 1 3505
box -2 -3 26 103
use AOI21X1  AOI21X1_3
timestamp 1693479267
transform -1 0 444 0 1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_23
timestamp 1693479267
transform 1 0 444 0 1 3505
box -2 -3 26 103
use OR2X2  OR2X2_8
timestamp 1693479267
transform -1 0 500 0 1 3505
box -2 -3 34 103
use FILL  FILL_35_0_0
timestamp 1693479267
transform 1 0 500 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_0_1
timestamp 1693479267
transform 1 0 508 0 1 3505
box -2 -3 10 103
use NAND2X1  NAND2X1_923
timestamp 1693479267
transform 1 0 516 0 1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_922
timestamp 1693479267
transform -1 0 564 0 1 3505
box -2 -3 26 103
use CLKBUF1  CLKBUF1_40
timestamp 1693479267
transform 1 0 564 0 1 3505
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_292
timestamp 1693479267
transform 1 0 636 0 1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_889
timestamp 1693479267
transform -1 0 764 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_890
timestamp 1693479267
transform 1 0 764 0 1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_319
timestamp 1693479267
transform 1 0 796 0 1 3505
box -2 -3 98 103
use CLKBUF1  CLKBUF1_42
timestamp 1693479267
transform -1 0 964 0 1 3505
box -2 -3 74 103
use CLKBUF1  CLKBUF1_55
timestamp 1693479267
transform 1 0 964 0 1 3505
box -2 -3 74 103
use FILL  FILL_35_1_0
timestamp 1693479267
transform 1 0 1036 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_1_1
timestamp 1693479267
transform 1 0 1044 0 1 3505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_136
timestamp 1693479267
transform 1 0 1052 0 1 3505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_24
timestamp 1693479267
transform 1 0 1148 0 1 3505
box -2 -3 98 103
use AOI22X1  AOI22X1_11
timestamp 1693479267
transform -1 0 1284 0 1 3505
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_49
timestamp 1693479267
transform -1 0 1380 0 1 3505
box -2 -3 98 103
use INVX1  INVX1_102
timestamp 1693479267
transform 1 0 1380 0 1 3505
box -2 -3 18 103
use AOI22X1  AOI22X1_34
timestamp 1693479267
transform -1 0 1436 0 1 3505
box -2 -3 42 103
use INVX1  INVX1_118
timestamp 1693479267
transform 1 0 1436 0 1 3505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_73
timestamp 1693479267
transform -1 0 1548 0 1 3505
box -2 -3 98 103
use FILL  FILL_35_2_0
timestamp 1693479267
transform 1 0 1548 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_2_1
timestamp 1693479267
transform 1 0 1556 0 1 3505
box -2 -3 10 103
use CLKBUF1  CLKBUF1_30
timestamp 1693479267
transform 1 0 1564 0 1 3505
box -2 -3 74 103
use INVX1  INVX1_218
timestamp 1693479267
transform -1 0 1652 0 1 3505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_53
timestamp 1693479267
transform -1 0 1748 0 1 3505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_105
timestamp 1693479267
transform -1 0 1844 0 1 3505
box -2 -3 98 103
use INVX1  INVX1_105
timestamp 1693479267
transform 1 0 1844 0 1 3505
box -2 -3 18 103
use INVX1  INVX1_106
timestamp 1693479267
transform 1 0 1860 0 1 3505
box -2 -3 18 103
use OAI21X1  OAI21X1_112
timestamp 1693479267
transform 1 0 1876 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_104
timestamp 1693479267
transform 1 0 1908 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_103
timestamp 1693479267
transform -1 0 1972 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_136
timestamp 1693479267
transform 1 0 1972 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_110
timestamp 1693479267
transform -1 0 2036 0 1 3505
box -2 -3 34 103
use FILL  FILL_35_3_0
timestamp 1693479267
transform 1 0 2036 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_3_1
timestamp 1693479267
transform 1 0 2044 0 1 3505
box -2 -3 10 103
use INVX1  INVX1_126
timestamp 1693479267
transform 1 0 2052 0 1 3505
box -2 -3 18 103
use BUFX4  BUFX4_184
timestamp 1693479267
transform 1 0 2068 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_152
timestamp 1693479267
transform 1 0 2100 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_151
timestamp 1693479267
transform 1 0 2132 0 1 3505
box -2 -3 34 103
use BUFX4  BUFX4_269
timestamp 1693479267
transform -1 0 2196 0 1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_240
timestamp 1693479267
transform -1 0 2292 0 1 3505
box -2 -3 98 103
use NAND2X1  NAND2X1_779
timestamp 1693479267
transform -1 0 2316 0 1 3505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_223
timestamp 1693479267
transform -1 0 2412 0 1 3505
box -2 -3 98 103
use NAND2X1  NAND2X1_720
timestamp 1693479267
transform 1 0 2412 0 1 3505
box -2 -3 26 103
use NAND3X1  NAND3X1_197
timestamp 1693479267
transform 1 0 2436 0 1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_716
timestamp 1693479267
transform -1 0 2492 0 1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_878
timestamp 1693479267
transform -1 0 2516 0 1 3505
box -2 -3 26 103
use INVX1  INVX1_549
timestamp 1693479267
transform -1 0 2532 0 1 3505
box -2 -3 18 103
use INVX1  INVX1_507
timestamp 1693479267
transform -1 0 2548 0 1 3505
box -2 -3 18 103
use FILL  FILL_35_4_0
timestamp 1693479267
transform 1 0 2548 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_4_1
timestamp 1693479267
transform 1 0 2556 0 1 3505
box -2 -3 10 103
use INVX1  INVX1_622
timestamp 1693479267
transform 1 0 2564 0 1 3505
box -2 -3 18 103
use NAND2X1  NAND2X1_889
timestamp 1693479267
transform 1 0 2580 0 1 3505
box -2 -3 26 103
use INVX1  INVX1_580
timestamp 1693479267
transform 1 0 2604 0 1 3505
box -2 -3 18 103
use NAND2X1  NAND2X1_826
timestamp 1693479267
transform 1 0 2620 0 1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_765
timestamp 1693479267
transform -1 0 2668 0 1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_763
timestamp 1693479267
transform -1 0 2692 0 1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_755
timestamp 1693479267
transform -1 0 2716 0 1 3505
box -2 -3 26 103
use INVX1  INVX1_533
timestamp 1693479267
transform -1 0 2732 0 1 3505
box -2 -3 18 103
use INVX1  INVX1_606
timestamp 1693479267
transform 1 0 2732 0 1 3505
box -2 -3 18 103
use NAND2X1  NAND2X1_865
timestamp 1693479267
transform 1 0 2748 0 1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_895
timestamp 1693479267
transform -1 0 2796 0 1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_785
timestamp 1693479267
transform 1 0 2796 0 1 3505
box -2 -3 26 103
use INVX1  INVX1_593
timestamp 1693479267
transform 1 0 2820 0 1 3505
box -2 -3 18 103
use NAND3X1  NAND3X1_276
timestamp 1693479267
transform 1 0 2836 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_637
timestamp 1693479267
transform -1 0 2884 0 1 3505
box -2 -3 18 103
use NAND3X1  NAND3X1_320
timestamp 1693479267
transform 1 0 2884 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_522
timestamp 1693479267
transform 1 0 2916 0 1 3505
box -2 -3 18 103
use NAND3X1  NAND3X1_208
timestamp 1693479267
transform 1 0 2932 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_595
timestamp 1693479267
transform 1 0 2964 0 1 3505
box -2 -3 18 103
use NAND3X1  NAND3X1_278
timestamp 1693479267
transform 1 0 2980 0 1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_749
timestamp 1693479267
transform -1 0 3036 0 1 3505
box -2 -3 26 103
use INVX1  INVX1_529
timestamp 1693479267
transform -1 0 3052 0 1 3505
box -2 -3 18 103
use FILL  FILL_35_5_0
timestamp 1693479267
transform 1 0 3052 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_5_1
timestamp 1693479267
transform 1 0 3060 0 1 3505
box -2 -3 10 103
use NAND2X1  NAND2X1_873
timestamp 1693479267
transform 1 0 3068 0 1 3505
box -2 -3 26 103
use INVX1  INVX1_602
timestamp 1693479267
transform 1 0 3092 0 1 3505
box -2 -3 18 103
use NAND2X1  NAND2X1_706
timestamp 1693479267
transform -1 0 3132 0 1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_859
timestamp 1693479267
transform 1 0 3132 0 1 3505
box -2 -3 26 103
use INVX1  INVX1_500
timestamp 1693479267
transform -1 0 3172 0 1 3505
box -2 -3 18 103
use INVX1  INVX1_573
timestamp 1693479267
transform 1 0 3172 0 1 3505
box -2 -3 18 103
use NAND2X1  NAND2X1_791
timestamp 1693479267
transform -1 0 3212 0 1 3505
box -2 -3 26 103
use INVX1  INVX1_557
timestamp 1693479267
transform -1 0 3228 0 1 3505
box -2 -3 18 103
use NAND2X1  NAND2X1_910
timestamp 1693479267
transform -1 0 3252 0 1 3505
box -2 -3 26 103
use INVX1  INVX1_630
timestamp 1693479267
transform 1 0 3252 0 1 3505
box -2 -3 18 103
use NAND2X1  NAND2X1_901
timestamp 1693479267
transform 1 0 3268 0 1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_816
timestamp 1693479267
transform 1 0 3292 0 1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_914
timestamp 1693479267
transform 1 0 3316 0 1 3505
box -2 -3 26 103
use BUFX4  BUFX4_62
timestamp 1693479267
transform 1 0 3340 0 1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_41
timestamp 1693479267
transform -1 0 3396 0 1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_52
timestamp 1693479267
transform -1 0 3420 0 1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_848
timestamp 1693479267
transform 1 0 3420 0 1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_905
timestamp 1693479267
transform 1 0 3444 0 1 3505
box -2 -3 26 103
use INVX1  INVX1_52
timestamp 1693479267
transform 1 0 3468 0 1 3505
box -2 -3 18 103
use OAI21X1  OAI21X1_52
timestamp 1693479267
transform 1 0 3484 0 1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_383
timestamp 1693479267
transform 1 0 3516 0 1 3505
box -2 -3 98 103
use FILL  FILL_35_6_0
timestamp 1693479267
transform 1 0 3612 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_6_1
timestamp 1693479267
transform 1 0 3620 0 1 3505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_395
timestamp 1693479267
transform 1 0 3628 0 1 3505
box -2 -3 98 103
use OAI21X1  OAI21X1_41
timestamp 1693479267
transform -1 0 3756 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_41
timestamp 1693479267
transform -1 0 3772 0 1 3505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_384
timestamp 1693479267
transform 1 0 3772 0 1 3505
box -2 -3 98 103
use NAND2X1  NAND2X1_42
timestamp 1693479267
transform -1 0 3892 0 1 3505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_382
timestamp 1693479267
transform 1 0 3892 0 1 3505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_197
timestamp 1693479267
transform 1 0 3988 0 1 3505
box -2 -3 98 103
use FILL  FILL_35_7_0
timestamp 1693479267
transform 1 0 4084 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_7_1
timestamp 1693479267
transform 1 0 4092 0 1 3505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_213
timestamp 1693479267
transform 1 0 4100 0 1 3505
box -2 -3 98 103
use INVX1  INVX1_725
timestamp 1693479267
transform 1 0 4196 0 1 3505
box -2 -3 18 103
use OAI21X1  OAI21X1_967
timestamp 1693479267
transform 1 0 4212 0 1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_214
timestamp 1693479267
transform 1 0 4244 0 1 3505
box -2 -3 98 103
use INVX4  INVX4_14
timestamp 1693479267
transform 1 0 4340 0 1 3505
box -2 -3 26 103
use BUFX4  BUFX4_106
timestamp 1693479267
transform 1 0 4364 0 1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_198
timestamp 1693479267
transform 1 0 4396 0 1 3505
box -2 -3 98 103
use NAND2X1  NAND2X1_1022
timestamp 1693479267
transform 1 0 4492 0 1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_1001
timestamp 1693479267
transform 1 0 4516 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_952
timestamp 1693479267
transform -1 0 4572 0 1 3505
box -2 -3 34 103
use BUFX4  BUFX4_104
timestamp 1693479267
transform 1 0 4572 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_173
timestamp 1693479267
transform 1 0 4 0 -1 3705
box -2 -3 18 103
use NOR3X1  NOR3X1_32
timestamp 1693479267
transform 1 0 20 0 -1 3705
box -2 -3 66 103
use INVX1  INVX1_166
timestamp 1693479267
transform 1 0 84 0 -1 3705
box -2 -3 18 103
use NOR3X1  NOR3X1_25
timestamp 1693479267
transform -1 0 164 0 -1 3705
box -2 -3 66 103
use DFFPOSX1  DFFPOSX1_418
timestamp 1693479267
transform 1 0 164 0 -1 3705
box -2 -3 98 103
use CLKBUF1  CLKBUF1_59
timestamp 1693479267
transform 1 0 260 0 -1 3705
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_340
timestamp 1693479267
transform 1 0 332 0 -1 3705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_338
timestamp 1693479267
transform 1 0 428 0 -1 3705
box -2 -3 98 103
use FILL  FILL_36_0_0
timestamp 1693479267
transform 1 0 524 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_0_1
timestamp 1693479267
transform 1 0 532 0 -1 3705
box -2 -3 10 103
use BUFX2  BUFX2_87
timestamp 1693479267
transform 1 0 540 0 -1 3705
box -2 -3 26 103
use BUFX2  BUFX2_89
timestamp 1693479267
transform -1 0 588 0 -1 3705
box -2 -3 26 103
use INVX1  INVX1_659
timestamp 1693479267
transform 1 0 588 0 -1 3705
box -2 -3 18 103
use OAI21X1  OAI21X1_888
timestamp 1693479267
transform 1 0 604 0 -1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_320
timestamp 1693479267
transform 1 0 636 0 -1 3705
box -2 -3 98 103
use INVX1  INVX1_661
timestamp 1693479267
transform 1 0 732 0 -1 3705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_141
timestamp 1693479267
transform 1 0 748 0 -1 3705
box -2 -3 98 103
use OAI21X1  OAI21X1_887
timestamp 1693479267
transform -1 0 876 0 -1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_137
timestamp 1693479267
transform 1 0 876 0 -1 3705
box -2 -3 98 103
use BUFX4  BUFX4_4
timestamp 1693479267
transform 1 0 972 0 -1 3705
box -2 -3 34 103
use FILL  FILL_36_1_0
timestamp 1693479267
transform 1 0 1004 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_1_1
timestamp 1693479267
transform 1 0 1012 0 -1 3705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_148
timestamp 1693479267
transform 1 0 1020 0 -1 3705
box -2 -3 98 103
use OAI21X1  OAI21X1_211
timestamp 1693479267
transform -1 0 1148 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_209
timestamp 1693479267
transform -1 0 1164 0 -1 3705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_95
timestamp 1693479267
transform -1 0 1260 0 -1 3705
box -2 -3 98 103
use OAI21X1  OAI21X1_196
timestamp 1693479267
transform -1 0 1292 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_194
timestamp 1693479267
transform -1 0 1308 0 -1 3705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_99
timestamp 1693479267
transform -1 0 1404 0 -1 3705
box -2 -3 98 103
use OAI21X1  OAI21X1_219
timestamp 1693479267
transform -1 0 1436 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_217
timestamp 1693479267
transform -1 0 1452 0 -1 3705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_96
timestamp 1693479267
transform -1 0 1548 0 -1 3705
box -2 -3 98 103
use FILL  FILL_36_2_0
timestamp 1693479267
transform 1 0 1548 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_2_1
timestamp 1693479267
transform 1 0 1556 0 -1 3705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_121
timestamp 1693479267
transform 1 0 1564 0 -1 3705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_72
timestamp 1693479267
transform -1 0 1756 0 -1 3705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_81
timestamp 1693479267
transform -1 0 1852 0 -1 3705
box -2 -3 98 103
use OAI21X1  OAI21X1_139
timestamp 1693479267
transform -1 0 1884 0 -1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_104
timestamp 1693479267
transform -1 0 1980 0 -1 3705
box -2 -3 98 103
use OAI21X1  OAI21X1_149
timestamp 1693479267
transform 1 0 1980 0 -1 3705
box -2 -3 34 103
use FILL  FILL_36_3_0
timestamp 1693479267
transform -1 0 2020 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_3_1
timestamp 1693479267
transform -1 0 2028 0 -1 3705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_239
timestamp 1693479267
transform -1 0 2124 0 -1 3705
box -2 -3 98 103
use NAND3X1  NAND3X1_255
timestamp 1693479267
transform 1 0 2124 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_548
timestamp 1693479267
transform 1 0 2156 0 -1 3705
box -2 -3 18 103
use NAND3X1  NAND3X1_235
timestamp 1693479267
transform -1 0 2204 0 -1 3705
box -2 -3 34 103
use NAND3X1  NAND3X1_234
timestamp 1693479267
transform 1 0 2204 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_552
timestamp 1693479267
transform 1 0 2236 0 -1 3705
box -2 -3 18 103
use NAND3X1  NAND3X1_238
timestamp 1693479267
transform 1 0 2252 0 -1 3705
box -2 -3 34 103
use NAND3X1  NAND3X1_239
timestamp 1693479267
transform -1 0 2316 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_611
timestamp 1693479267
transform 1 0 2316 0 -1 3705
box -2 -3 18 103
use INVX1  INVX1_538
timestamp 1693479267
transform 1 0 2332 0 -1 3705
box -2 -3 18 103
use NAND2X1  NAND2X1_769
timestamp 1693479267
transform 1 0 2348 0 -1 3705
box -2 -3 26 103
use NAND3X1  NAND3X1_224
timestamp 1693479267
transform 1 0 2372 0 -1 3705
box -2 -3 34 103
use NAND3X1  NAND3X1_196
timestamp 1693479267
transform -1 0 2436 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_510
timestamp 1693479267
transform -1 0 2452 0 -1 3705
box -2 -3 18 103
use NAND3X1  NAND3X1_225
timestamp 1693479267
transform 1 0 2452 0 -1 3705
box -2 -3 34 103
use NAND3X1  NAND3X1_199
timestamp 1693479267
transform 1 0 2484 0 -1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_761
timestamp 1693479267
transform -1 0 2540 0 -1 3705
box -2 -3 26 103
use FILL  FILL_36_4_0
timestamp 1693479267
transform 1 0 2540 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_4_1
timestamp 1693479267
transform 1 0 2548 0 -1 3705
box -2 -3 10 103
use NAND3X1  NAND3X1_294
timestamp 1693479267
transform 1 0 2556 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_537
timestamp 1693479267
transform -1 0 2604 0 -1 3705
box -2 -3 18 103
use INVX1  INVX1_610
timestamp 1693479267
transform 1 0 2604 0 -1 3705
box -2 -3 18 103
use NAND2X1  NAND2X1_871
timestamp 1693479267
transform 1 0 2620 0 -1 3705
box -2 -3 26 103
use NAND3X1  NAND3X1_295
timestamp 1693479267
transform 1 0 2644 0 -1 3705
box -2 -3 34 103
use NAND3X1  NAND3X1_269
timestamp 1693479267
transform -1 0 2708 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_583
timestamp 1693479267
transform 1 0 2708 0 -1 3705
box -2 -3 18 103
use BUFX4  BUFX4_120
timestamp 1693479267
transform -1 0 2756 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_553
timestamp 1693479267
transform 1 0 2756 0 -1 3705
box -2 -3 18 103
use INVX1  INVX1_626
timestamp 1693479267
transform 1 0 2772 0 -1 3705
box -2 -3 18 103
use NAND3X1  NAND3X1_266
timestamp 1693479267
transform 1 0 2788 0 -1 3705
box -2 -3 34 103
use NAND3X1  NAND3X1_277
timestamp 1693479267
transform 1 0 2820 0 -1 3705
box -2 -3 34 103
use NAND3X1  NAND3X1_216
timestamp 1693479267
transform -1 0 2884 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_530
timestamp 1693479267
transform -1 0 2900 0 -1 3705
box -2 -3 18 103
use INVX1  INVX1_597
timestamp 1693479267
transform 1 0 2900 0 -1 3705
box -2 -3 18 103
use NAND3X1  NAND3X1_209
timestamp 1693479267
transform -1 0 2948 0 -1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_879
timestamp 1693479267
transform 1 0 2948 0 -1 3705
box -2 -3 26 103
use INVX1  INVX1_603
timestamp 1693479267
transform 1 0 2972 0 -1 3705
box -2 -3 18 103
use NAND3X1  NAND3X1_286
timestamp 1693479267
transform 1 0 2988 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_631
timestamp 1693479267
transform 1 0 3020 0 -1 3705
box -2 -3 18 103
use NAND2X1  NAND2X1_840
timestamp 1693479267
transform 1 0 3036 0 -1 3705
box -2 -3 26 103
use FILL  FILL_36_5_0
timestamp 1693479267
transform 1 0 3060 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_5_1
timestamp 1693479267
transform 1 0 3068 0 -1 3705
box -2 -3 10 103
use NAND3X1  NAND3X1_314
timestamp 1693479267
transform 1 0 3076 0 -1 3705
box -2 -3 34 103
use NAND3X1  NAND3X1_280
timestamp 1693479267
transform 1 0 3108 0 -1 3705
box -2 -3 34 103
use NAND3X1  NAND3X1_281
timestamp 1693479267
transform -1 0 3172 0 -1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_875
timestamp 1693479267
transform 1 0 3172 0 -1 3705
box -2 -3 26 103
use NAND3X1  NAND3X1_267
timestamp 1693479267
transform -1 0 3228 0 -1 3705
box -2 -3 34 103
use NAND3X1  NAND3X1_279
timestamp 1693479267
transform -1 0 3260 0 -1 3705
box -2 -3 34 103
use BUFX4  BUFX4_121
timestamp 1693479267
transform 1 0 3260 0 -1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_51
timestamp 1693479267
transform -1 0 3316 0 -1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_51
timestamp 1693479267
transform -1 0 3348 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_51
timestamp 1693479267
transform -1 0 3364 0 -1 3705
box -2 -3 18 103
use NAND2X1  NAND2X1_830
timestamp 1693479267
transform -1 0 3388 0 -1 3705
box -2 -3 26 103
use NAND2X1  NAND2X1_36
timestamp 1693479267
transform -1 0 3412 0 -1 3705
box -2 -3 26 103
use BUFX4  BUFX4_31
timestamp 1693479267
transform -1 0 3444 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_36
timestamp 1693479267
transform -1 0 3476 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_36
timestamp 1693479267
transform -1 0 3492 0 -1 3705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_115
timestamp 1693479267
transform -1 0 3588 0 -1 3705
box -2 -3 98 103
use FILL  FILL_36_6_0
timestamp 1693479267
transform 1 0 3588 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_6_1
timestamp 1693479267
transform 1 0 3596 0 -1 3705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_379
timestamp 1693479267
transform 1 0 3604 0 -1 3705
box -2 -3 98 103
use BUFX4  BUFX4_32
timestamp 1693479267
transform 1 0 3700 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_39
timestamp 1693479267
transform -1 0 3764 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_39
timestamp 1693479267
transform -1 0 3780 0 -1 3705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_118
timestamp 1693479267
transform -1 0 3876 0 -1 3705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_209
timestamp 1693479267
transform 1 0 3876 0 -1 3705
box -2 -3 98 103
use INVX1  INVX1_721
timestamp 1693479267
transform 1 0 3972 0 -1 3705
box -2 -3 18 103
use OAI21X1  OAI21X1_959
timestamp 1693479267
transform 1 0 3988 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_958
timestamp 1693479267
transform 1 0 4020 0 -1 3705
box -2 -3 34 103
use BUFX2  BUFX2_80
timestamp 1693479267
transform -1 0 4076 0 -1 3705
box -2 -3 26 103
use FILL  FILL_36_7_0
timestamp 1693479267
transform -1 0 4084 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_7_1
timestamp 1693479267
transform -1 0 4092 0 -1 3705
box -2 -3 10 103
use OAI21X1  OAI21X1_1050
timestamp 1693479267
transform -1 0 4124 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1043
timestamp 1693479267
transform -1 0 4156 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1042
timestamp 1693479267
transform -1 0 4188 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1036
timestamp 1693479267
transform -1 0 4220 0 -1 3705
box -2 -3 34 103
use BUFX4  BUFX4_68
timestamp 1693479267
transform -1 0 4252 0 -1 3705
box -2 -3 34 103
use BUFX4  BUFX4_64
timestamp 1693479267
transform -1 0 4284 0 -1 3705
box -2 -3 34 103
use BUFX4  BUFX4_251
timestamp 1693479267
transform -1 0 4316 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_951
timestamp 1693479267
transform 1 0 4316 0 -1 3705
box -2 -3 34 103
use BUFX4  BUFX4_118
timestamp 1693479267
transform -1 0 4380 0 -1 3705
box -2 -3 34 103
use BUFX4  BUFX4_71
timestamp 1693479267
transform 1 0 4380 0 -1 3705
box -2 -3 34 103
use BUFX4  BUFX4_66
timestamp 1693479267
transform 1 0 4412 0 -1 3705
box -2 -3 34 103
use BUFX4  BUFX4_108
timestamp 1693479267
transform 1 0 4444 0 -1 3705
box -2 -3 34 103
use AOI22X1  AOI22X1_167
timestamp 1693479267
transform 1 0 4476 0 -1 3705
box -2 -3 42 103
use OAI21X1  OAI21X1_1051
timestamp 1693479267
transform -1 0 4548 0 -1 3705
box -2 -3 34 103
use BUFX4  BUFX4_250
timestamp 1693479267
transform 1 0 4548 0 -1 3705
box -2 -3 34 103
use FILL  FILL_37_1
timestamp 1693479267
transform -1 0 4588 0 -1 3705
box -2 -3 10 103
use FILL  FILL_37_2
timestamp 1693479267
transform -1 0 4596 0 -1 3705
box -2 -3 10 103
use FILL  FILL_37_3
timestamp 1693479267
transform -1 0 4604 0 -1 3705
box -2 -3 10 103
use INVX1  INVX1_171
timestamp 1693479267
transform 1 0 4 0 1 3705
box -2 -3 18 103
use NOR3X1  NOR3X1_30
timestamp 1693479267
transform -1 0 84 0 1 3705
box -2 -3 66 103
use NOR3X1  NOR3X1_38
timestamp 1693479267
transform -1 0 148 0 1 3705
box -2 -3 66 103
use DFFPOSX1  DFFPOSX1_423
timestamp 1693479267
transform 1 0 148 0 1 3705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_431
timestamp 1693479267
transform 1 0 244 0 1 3705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_341
timestamp 1693479267
transform 1 0 340 0 1 3705
box -2 -3 98 103
use CLKBUF1  CLKBUF1_9
timestamp 1693479267
transform -1 0 508 0 1 3705
box -2 -3 74 103
use FILL  FILL_37_0_0
timestamp 1693479267
transform 1 0 508 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_0_1
timestamp 1693479267
transform 1 0 516 0 1 3705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_154
timestamp 1693479267
transform 1 0 524 0 1 3705
box -2 -3 98 103
use XOR2X1  XOR2X1_11
timestamp 1693479267
transform -1 0 676 0 1 3705
box -2 -3 58 103
use XOR2X1  XOR2X1_10
timestamp 1693479267
transform -1 0 732 0 1 3705
box -2 -3 58 103
use NOR2X1  NOR2X1_399
timestamp 1693479267
transform 1 0 732 0 1 3705
box -2 -3 26 103
use NAND2X1  NAND2X1_703
timestamp 1693479267
transform 1 0 756 0 1 3705
box -2 -3 26 103
use AND2X2  AND2X2_79
timestamp 1693479267
transform 1 0 780 0 1 3705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_29
timestamp 1693479267
transform 1 0 812 0 1 3705
box -2 -3 98 103
use INVX1  INVX1_658
timestamp 1693479267
transform -1 0 924 0 1 3705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_25
timestamp 1693479267
transform 1 0 924 0 1 3705
box -2 -3 98 103
use FILL  FILL_37_1_0
timestamp 1693479267
transform 1 0 1020 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_1_1
timestamp 1693479267
transform 1 0 1028 0 1 3705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_140
timestamp 1693479267
transform 1 0 1036 0 1 3705
box -2 -3 98 103
use AOI22X1  AOI22X1_26
timestamp 1693479267
transform 1 0 1132 0 1 3705
box -2 -3 42 103
use INVX1  INVX1_208
timestamp 1693479267
transform -1 0 1188 0 1 3705
box -2 -3 18 103
use AOI22X1  AOI22X1_25
timestamp 1693479267
transform -1 0 1228 0 1 3705
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_63
timestamp 1693479267
transform -1 0 1324 0 1 3705
box -2 -3 98 103
use OAI21X1  OAI21X1_214
timestamp 1693479267
transform -1 0 1356 0 1 3705
box -2 -3 34 103
use INVX1  INVX1_212
timestamp 1693479267
transform 1 0 1356 0 1 3705
box -2 -3 18 103
use BUFX4  BUFX4_257
timestamp 1693479267
transform -1 0 1404 0 1 3705
box -2 -3 34 103
use AOI22X1  AOI22X1_24
timestamp 1693479267
transform -1 0 1444 0 1 3705
box -2 -3 42 103
use OAI21X1  OAI21X1_209
timestamp 1693479267
transform -1 0 1476 0 1 3705
box -2 -3 34 103
use INVX1  INVX1_116
timestamp 1693479267
transform 1 0 1476 0 1 3705
box -2 -3 18 103
use FILL  FILL_37_2_0
timestamp 1693479267
transform -1 0 1500 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_2_1
timestamp 1693479267
transform -1 0 1508 0 1 3705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_62
timestamp 1693479267
transform -1 0 1604 0 1 3705
box -2 -3 98 103
use CLKBUF1  CLKBUF1_3
timestamp 1693479267
transform 1 0 1604 0 1 3705
box -2 -3 74 103
use INVX1  INVX1_115
timestamp 1693479267
transform 1 0 1676 0 1 3705
box -2 -3 18 103
use INVX1  INVX1_207
timestamp 1693479267
transform -1 0 1708 0 1 3705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_94
timestamp 1693479267
transform -1 0 1804 0 1 3705
box -2 -3 98 103
use OAI21X1  OAI21X1_132
timestamp 1693479267
transform 1 0 1804 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_131
timestamp 1693479267
transform -1 0 1868 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_130
timestamp 1693479267
transform 1 0 1868 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_129
timestamp 1693479267
transform -1 0 1932 0 1 3705
box -2 -3 34 103
use INVX1  INVX1_125
timestamp 1693479267
transform 1 0 1932 0 1 3705
box -2 -3 18 103
use OAI21X1  OAI21X1_150
timestamp 1693479267
transform 1 0 1948 0 1 3705
box -2 -3 34 103
use BUFX4  BUFX4_185
timestamp 1693479267
transform -1 0 2012 0 1 3705
box -2 -3 34 103
use FILL  FILL_37_3_0
timestamp 1693479267
transform 1 0 2012 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_3_1
timestamp 1693479267
transform 1 0 2020 0 1 3705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_110
timestamp 1693479267
transform 1 0 2028 0 1 3705
box -2 -3 98 103
use INVX1  INVX1_621
timestamp 1693479267
transform -1 0 2140 0 1 3705
box -2 -3 18 103
use INVX1  INVX1_625
timestamp 1693479267
transform 1 0 2140 0 1 3705
box -2 -3 18 103
use NAND2X1  NAND2X1_776
timestamp 1693479267
transform 1 0 2156 0 1 3705
box -2 -3 26 103
use INVX1  INVX1_605
timestamp 1693479267
transform 1 0 2180 0 1 3705
box -2 -3 18 103
use BUFX4  BUFX4_219
timestamp 1693479267
transform -1 0 2228 0 1 3705
box -2 -3 34 103
use BUFX4  BUFX4_207
timestamp 1693479267
transform 1 0 2228 0 1 3705
box -2 -3 34 103
use INVX1  INVX1_532
timestamp 1693479267
transform 1 0 2260 0 1 3705
box -2 -3 18 103
use BUFX4  BUFX4_35
timestamp 1693479267
transform 1 0 2276 0 1 3705
box -2 -3 34 103
use NAND3X1  NAND3X1_218
timestamp 1693479267
transform 1 0 2308 0 1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_771
timestamp 1693479267
transform -1 0 2364 0 1 3705
box -2 -3 26 103
use BUFX4  BUFX4_34
timestamp 1693479267
transform -1 0 2396 0 1 3705
box -2 -3 34 103
use BUFX4  BUFX4_218
timestamp 1693479267
transform 1 0 2396 0 1 3705
box -2 -3 34 103
use BUFX4  BUFX4_33
timestamp 1693479267
transform 1 0 2428 0 1 3705
box -2 -3 34 103
use BUFX4  BUFX4_206
timestamp 1693479267
transform 1 0 2460 0 1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_722
timestamp 1693479267
transform -1 0 2516 0 1 3705
box -2 -3 26 103
use NAND2X1  NAND2X1_893
timestamp 1693479267
transform -1 0 2540 0 1 3705
box -2 -3 26 103
use FILL  FILL_37_4_0
timestamp 1693479267
transform -1 0 2548 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_4_1
timestamp 1693479267
transform -1 0 2556 0 1 3705
box -2 -3 10 103
use INVX1  INVX1_511
timestamp 1693479267
transform -1 0 2572 0 1 3705
box -2 -3 18 103
use INVX1  INVX1_584
timestamp 1693479267
transform 1 0 2572 0 1 3705
box -2 -3 18 103
use NAND2X1  NAND2X1_832
timestamp 1693479267
transform 1 0 2588 0 1 3705
box -2 -3 26 103
use NAND2X1  NAND2X1_844
timestamp 1693479267
transform -1 0 2636 0 1 3705
box -2 -3 26 103
use INVX1  INVX1_592
timestamp 1693479267
transform -1 0 2652 0 1 3705
box -2 -3 18 103
use INVX1  INVX1_519
timestamp 1693479267
transform 1 0 2652 0 1 3705
box -2 -3 18 103
use NAND2X1  NAND2X1_734
timestamp 1693479267
transform 1 0 2668 0 1 3705
box -2 -3 26 103
use NAND3X1  NAND3X1_244
timestamp 1693479267
transform -1 0 2724 0 1 3705
box -2 -3 34 103
use INVX1  INVX1_558
timestamp 1693479267
transform -1 0 2740 0 1 3705
box -2 -3 18 103
use INVX1  INVX1_524
timestamp 1693479267
transform 1 0 2740 0 1 3705
box -2 -3 18 103
use NAND3X1  NAND3X1_214
timestamp 1693479267
transform -1 0 2788 0 1 3705
box -2 -3 34 103
use INVX1  INVX1_528
timestamp 1693479267
transform -1 0 2804 0 1 3705
box -2 -3 18 103
use NAND2X1  NAND2X1_719
timestamp 1693479267
transform -1 0 2828 0 1 3705
box -2 -3 26 103
use INVX1  INVX1_601
timestamp 1693479267
transform 1 0 2828 0 1 3705
box -2 -3 18 103
use NAND3X1  NAND3X1_284
timestamp 1693479267
transform 1 0 2844 0 1 3705
box -2 -3 34 103
use INVX1  INVX1_509
timestamp 1693479267
transform -1 0 2892 0 1 3705
box -2 -3 18 103
use NAND2X1  NAND2X1_737
timestamp 1693479267
transform -1 0 2916 0 1 3705
box -2 -3 26 103
use INVX1  INVX1_582
timestamp 1693479267
transform 1 0 2916 0 1 3705
box -2 -3 18 103
use INVX1  INVX1_521
timestamp 1693479267
transform -1 0 2948 0 1 3705
box -2 -3 18 103
use NAND2X1  NAND2X1_881
timestamp 1693479267
transform -1 0 2972 0 1 3705
box -2 -3 26 103
use NAND2X1  NAND2X1_850
timestamp 1693479267
transform 1 0 2972 0 1 3705
box -2 -3 26 103
use NAND2X1  NAND2X1_829
timestamp 1693479267
transform 1 0 2996 0 1 3705
box -2 -3 26 103
use NAND2X1  NAND2X1_839
timestamp 1693479267
transform 1 0 3020 0 1 3705
box -2 -3 26 103
use INVX1  INVX1_594
timestamp 1693479267
transform 1 0 3044 0 1 3705
box -2 -3 18 103
use FILL  FILL_37_5_0
timestamp 1693479267
transform 1 0 3060 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_5_1
timestamp 1693479267
transform 1 0 3068 0 1 3705
box -2 -3 10 103
use NAND2X1  NAND2X1_847
timestamp 1693479267
transform 1 0 3076 0 1 3705
box -2 -3 26 103
use NAND2X1  NAND2X1_842
timestamp 1693479267
transform 1 0 3100 0 1 3705
box -2 -3 26 103
use NAND2X1  NAND2X1_53
timestamp 1693479267
transform -1 0 3148 0 1 3705
box -2 -3 26 103
use NAND2X1  NAND2X1_40
timestamp 1693479267
transform -1 0 3172 0 1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_40
timestamp 1693479267
transform -1 0 3204 0 1 3705
box -2 -3 34 103
use INVX1  INVX1_40
timestamp 1693479267
transform -1 0 3220 0 1 3705
box -2 -3 18 103
use BUFX4  BUFX4_27
timestamp 1693479267
transform 1 0 3220 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_53
timestamp 1693479267
transform -1 0 3284 0 1 3705
box -2 -3 34 103
use INVX1  INVX1_53
timestamp 1693479267
transform -1 0 3300 0 1 3705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_396
timestamp 1693479267
transform 1 0 3300 0 1 3705
box -2 -3 98 103
use NAND2X1  NAND2X1_57
timestamp 1693479267
transform -1 0 3420 0 1 3705
box -2 -3 26 103
use NAND2X1  NAND2X1_39
timestamp 1693479267
transform -1 0 3444 0 1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_57
timestamp 1693479267
transform -1 0 3476 0 1 3705
box -2 -3 34 103
use INVX1  INVX1_57
timestamp 1693479267
transform -1 0 3492 0 1 3705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_400
timestamp 1693479267
transform 1 0 3492 0 1 3705
box -2 -3 98 103
use FILL  FILL_37_6_0
timestamp 1693479267
transform 1 0 3588 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_6_1
timestamp 1693479267
transform 1 0 3596 0 1 3705
box -2 -3 10 103
use CLKBUF1  CLKBUF1_38
timestamp 1693479267
transform 1 0 3604 0 1 3705
box -2 -3 74 103
use INVX8  INVX8_15
timestamp 1693479267
transform -1 0 3716 0 1 3705
box -2 -3 42 103
use NAND2X1  NAND2X1_996
timestamp 1693479267
transform -1 0 3740 0 1 3705
box -2 -3 26 103
use INVX8  INVX8_17
timestamp 1693479267
transform -1 0 3780 0 1 3705
box -2 -3 42 103
use NOR2X1  NOR2X1_473
timestamp 1693479267
transform 1 0 3780 0 1 3705
box -2 -3 26 103
use NOR2X1  NOR2X1_486
timestamp 1693479267
transform -1 0 3828 0 1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_1066
timestamp 1693479267
transform 1 0 3828 0 1 3705
box -2 -3 34 103
use INVX1  INVX1_758
timestamp 1693479267
transform -1 0 3876 0 1 3705
box -2 -3 18 103
use BUFX4  BUFX4_253
timestamp 1693479267
transform 1 0 3876 0 1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_478
timestamp 1693479267
transform 1 0 3908 0 1 3705
box -2 -3 26 103
use AOI22X1  AOI22X1_152
timestamp 1693479267
transform 1 0 3932 0 1 3705
box -2 -3 42 103
use AOI22X1  AOI22X1_159
timestamp 1693479267
transform 1 0 3972 0 1 3705
box -2 -3 42 103
use AOI22X1  AOI22X1_166
timestamp 1693479267
transform 1 0 4012 0 1 3705
box -2 -3 42 103
use AOI22X1  AOI22X1_158
timestamp 1693479267
transform -1 0 4092 0 1 3705
box -2 -3 42 103
use FILL  FILL_37_7_0
timestamp 1693479267
transform -1 0 4100 0 1 3705
box -2 -3 10 103
use FILL  FILL_37_7_1
timestamp 1693479267
transform -1 0 4108 0 1 3705
box -2 -3 10 103
use OAI21X1  OAI21X1_1015
timestamp 1693479267
transform -1 0 4140 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1032
timestamp 1693479267
transform -1 0 4172 0 1 3705
box -2 -3 34 103
use BUFX4  BUFX4_169
timestamp 1693479267
transform 1 0 4172 0 1 3705
box -2 -3 34 103
use BUFX4  BUFX4_109
timestamp 1693479267
transform -1 0 4236 0 1 3705
box -2 -3 34 103
use BUFX4  BUFX4_67
timestamp 1693479267
transform -1 0 4268 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1047
timestamp 1693479267
transform 1 0 4268 0 1 3705
box -2 -3 34 103
use BUFX4  BUFX4_70
timestamp 1693479267
transform -1 0 4332 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1045
timestamp 1693479267
transform 1 0 4332 0 1 3705
box -2 -3 34 103
use AOI22X1  AOI22X1_161
timestamp 1693479267
transform 1 0 4364 0 1 3705
box -2 -3 42 103
use BUFX4  BUFX4_170
timestamp 1693479267
transform 1 0 4404 0 1 3705
box -2 -3 34 103
use INVX1  INVX1_741
timestamp 1693479267
transform -1 0 4452 0 1 3705
box -2 -3 18 103
use OAI21X1  OAI21X1_1037
timestamp 1693479267
transform 1 0 4452 0 1 3705
box -2 -3 34 103
use AOI22X1  AOI22X1_154
timestamp 1693479267
transform 1 0 4484 0 1 3705
box -2 -3 42 103
use OAI21X1  OAI21X1_1038
timestamp 1693479267
transform -1 0 4556 0 1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_1041
timestamp 1693479267
transform 1 0 4556 0 1 3705
box -2 -3 34 103
use FILL  FILL_38_1
timestamp 1693479267
transform 1 0 4588 0 1 3705
box -2 -3 10 103
use FILL  FILL_38_2
timestamp 1693479267
transform 1 0 4596 0 1 3705
box -2 -3 10 103
use INVX1  INVX1_179
timestamp 1693479267
transform 1 0 4 0 -1 3905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_425
timestamp 1693479267
transform 1 0 20 0 -1 3905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_416
timestamp 1693479267
transform 1 0 116 0 -1 3905
box -2 -3 98 103
use XOR2X1  XOR2X1_2
timestamp 1693479267
transform -1 0 268 0 -1 3905
box -2 -3 58 103
use XNOR2X1  XNOR2X1_1
timestamp 1693479267
transform 1 0 268 0 -1 3905
box -2 -3 58 103
use AND2X2  AND2X2_3
timestamp 1693479267
transform -1 0 356 0 -1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_100
timestamp 1693479267
transform 1 0 356 0 -1 3905
box -2 -3 26 103
use AND2X2  AND2X2_4
timestamp 1693479267
transform -1 0 412 0 -1 3905
box -2 -3 34 103
use XNOR2X1  XNOR2X1_3
timestamp 1693479267
transform -1 0 468 0 -1 3905
box -2 -3 58 103
use FILL  FILL_38_0_0
timestamp 1693479267
transform 1 0 468 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_0_1
timestamp 1693479267
transform 1 0 476 0 -1 3905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_339
timestamp 1693479267
transform 1 0 484 0 -1 3905
box -2 -3 98 103
use XOR2X1  XOR2X1_14
timestamp 1693479267
transform 1 0 580 0 -1 3905
box -2 -3 58 103
use XOR2X1  XOR2X1_15
timestamp 1693479267
transform -1 0 692 0 -1 3905
box -2 -3 58 103
use NOR2X1  NOR2X1_405
timestamp 1693479267
transform 1 0 692 0 -1 3905
box -2 -3 26 103
use INVX1  INVX1_499
timestamp 1693479267
transform 1 0 716 0 -1 3905
box -2 -3 18 103
use AOI21X1  AOI21X1_222
timestamp 1693479267
transform -1 0 764 0 -1 3905
box -2 -3 34 103
use INVX1  INVX1_498
timestamp 1693479267
transform -1 0 780 0 -1 3905
box -2 -3 18 103
use INVX1  INVX1_660
timestamp 1693479267
transform -1 0 796 0 -1 3905
box -2 -3 18 103
use INVX1  INVX1_572
timestamp 1693479267
transform 1 0 796 0 -1 3905
box -2 -3 18 103
use AOI21X1  AOI21X1_226
timestamp 1693479267
transform -1 0 844 0 -1 3905
box -2 -3 34 103
use INVX1  INVX1_571
timestamp 1693479267
transform -1 0 860 0 -1 3905
box -2 -3 18 103
use NAND3X1  NAND3X1_257
timestamp 1693479267
transform 1 0 860 0 -1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_406
timestamp 1693479267
transform -1 0 916 0 -1 3905
box -2 -3 26 103
use NAND2X1  NAND2X1_813
timestamp 1693479267
transform 1 0 916 0 -1 3905
box -2 -3 26 103
use AND2X2  AND2X2_80
timestamp 1693479267
transform 1 0 940 0 -1 3905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_19
timestamp 1693479267
transform -1 0 1044 0 -1 3905
box -2 -3 74 103
use FILL  FILL_38_1_0
timestamp 1693479267
transform 1 0 1044 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_1_1
timestamp 1693479267
transform 1 0 1052 0 -1 3905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_28
timestamp 1693479267
transform 1 0 1060 0 -1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_210
timestamp 1693479267
transform 1 0 1156 0 -1 3905
box -2 -3 34 103
use AOI22X1  AOI22X1_28
timestamp 1693479267
transform -1 0 1228 0 -1 3905
box -2 -3 42 103
use OAI21X1  OAI21X1_213
timestamp 1693479267
transform -1 0 1260 0 -1 3905
box -2 -3 34 103
use INVX1  INVX1_211
timestamp 1693479267
transform -1 0 1276 0 -1 3905
box -2 -3 18 103
use AOI22X1  AOI22X1_29
timestamp 1693479267
transform -1 0 1316 0 -1 3905
box -2 -3 42 103
use OR2X2  OR2X2_3
timestamp 1693479267
transform 1 0 1316 0 -1 3905
box -2 -3 34 103
use BUFX4  BUFX4_142
timestamp 1693479267
transform -1 0 1380 0 -1 3905
box -2 -3 34 103
use BUFX4  BUFX4_240
timestamp 1693479267
transform -1 0 1412 0 -1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_19
timestamp 1693479267
transform 1 0 1412 0 -1 3905
box -2 -3 98 103
use FILL  FILL_38_2_0
timestamp 1693479267
transform -1 0 1516 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_2_1
timestamp 1693479267
transform -1 0 1524 0 -1 3905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_67
timestamp 1693479267
transform -1 0 1620 0 -1 3905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_98
timestamp 1693479267
transform -1 0 1716 0 -1 3905
box -2 -3 98 103
use INVX1  INVX1_120
timestamp 1693479267
transform 1 0 1716 0 -1 3905
box -2 -3 18 103
use OAI21X1  OAI21X1_133
timestamp 1693479267
transform -1 0 1764 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_137
timestamp 1693479267
transform 1 0 1764 0 -1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_242
timestamp 1693479267
transform -1 0 1892 0 -1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_140
timestamp 1693479267
transform -1 0 1924 0 -1 3905
box -2 -3 34 103
use BUFX4  BUFX4_270
timestamp 1693479267
transform -1 0 1956 0 -1 3905
box -2 -3 34 103
use INVX1  INVX1_547
timestamp 1693479267
transform 1 0 1956 0 -1 3905
box -2 -3 18 103
use INVX1  INVX1_629
timestamp 1693479267
transform 1 0 1972 0 -1 3905
box -2 -3 18 103
use NAND3X1  NAND3X1_312
timestamp 1693479267
transform 1 0 1988 0 -1 3905
box -2 -3 34 103
use FILL  FILL_38_3_0
timestamp 1693479267
transform -1 0 2028 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_3_1
timestamp 1693479267
transform -1 0 2036 0 -1 3905
box -2 -3 10 103
use NAND3X1  NAND3X1_305
timestamp 1693479267
transform -1 0 2068 0 -1 3905
box -2 -3 34 103
use NAND3X1  NAND3X1_304
timestamp 1693479267
transform -1 0 2100 0 -1 3905
box -2 -3 34 103
use NAND3X1  NAND3X1_308
timestamp 1693479267
transform -1 0 2132 0 -1 3905
box -2 -3 34 103
use NAND3X1  NAND3X1_309
timestamp 1693479267
transform -1 0 2164 0 -1 3905
box -2 -3 34 103
use NAND3X1  NAND3X1_288
timestamp 1693479267
transform -1 0 2196 0 -1 3905
box -2 -3 34 103
use NAND3X1  NAND3X1_271
timestamp 1693479267
transform -1 0 2228 0 -1 3905
box -2 -3 34 103
use NAND3X1  NAND3X1_313
timestamp 1693479267
transform -1 0 2260 0 -1 3905
box -2 -3 34 103
use NAND3X1  NAND3X1_289
timestamp 1693479267
transform 1 0 2260 0 -1 3905
box -2 -3 34 103
use BUFX4  BUFX4_95
timestamp 1693479267
transform 1 0 2292 0 -1 3905
box -2 -3 34 103
use NAND3X1  NAND3X1_219
timestamp 1693479267
transform -1 0 2356 0 -1 3905
box -2 -3 34 103
use BUFX4  BUFX4_209
timestamp 1693479267
transform 1 0 2356 0 -1 3905
box -2 -3 34 103
use INVX1  INVX1_512
timestamp 1693479267
transform 1 0 2388 0 -1 3905
box -2 -3 18 103
use NAND3X1  NAND3X1_198
timestamp 1693479267
transform 1 0 2404 0 -1 3905
box -2 -3 34 103
use INVX1  INVX1_585
timestamp 1693479267
transform 1 0 2436 0 -1 3905
box -2 -3 18 103
use NAND3X1  NAND3X1_204
timestamp 1693479267
transform -1 0 2484 0 -1 3905
box -2 -3 34 103
use INVX1  INVX1_518
timestamp 1693479267
transform -1 0 2500 0 -1 3905
box -2 -3 18 103
use INVX1  INVX1_591
timestamp 1693479267
transform 1 0 2500 0 -1 3905
box -2 -3 18 103
use BUFX4  BUFX4_220
timestamp 1693479267
transform 1 0 2516 0 -1 3905
box -2 -3 34 103
use FILL  FILL_38_4_0
timestamp 1693479267
transform 1 0 2548 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_4_1
timestamp 1693479267
transform 1 0 2556 0 -1 3905
box -2 -3 10 103
use NAND3X1  NAND3X1_268
timestamp 1693479267
transform 1 0 2564 0 -1 3905
box -2 -3 34 103
use NAND3X1  NAND3X1_205
timestamp 1693479267
transform 1 0 2596 0 -1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_731
timestamp 1693479267
transform -1 0 2652 0 -1 3905
box -2 -3 26 103
use NAND3X1  NAND3X1_203
timestamp 1693479267
transform -1 0 2684 0 -1 3905
box -2 -3 34 103
use NAND3X1  NAND3X1_202
timestamp 1693479267
transform -1 0 2716 0 -1 3905
box -2 -3 34 103
use INVX1  INVX1_516
timestamp 1693479267
transform -1 0 2732 0 -1 3905
box -2 -3 18 103
use NAND3X1  NAND3X1_210
timestamp 1693479267
transform -1 0 2764 0 -1 3905
box -2 -3 34 103
use NAND3X1  NAND3X1_215
timestamp 1693479267
transform -1 0 2796 0 -1 3905
box -2 -3 34 103
use NAND3X1  NAND3X1_285
timestamp 1693479267
transform -1 0 2828 0 -1 3905
box -2 -3 34 103
use NAND3X1  NAND3X1_211
timestamp 1693479267
transform 1 0 2828 0 -1 3905
box -2 -3 34 103
use NAND3X1  NAND3X1_283
timestamp 1693479267
transform -1 0 2892 0 -1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_740
timestamp 1693479267
transform -1 0 2916 0 -1 3905
box -2 -3 26 103
use BUFX4  BUFX4_94
timestamp 1693479267
transform 1 0 2916 0 -1 3905
box -2 -3 34 103
use INVX1  INVX1_523
timestamp 1693479267
transform -1 0 2964 0 -1 3905
box -2 -3 18 103
use INVX1  INVX1_596
timestamp 1693479267
transform 1 0 2964 0 -1 3905
box -2 -3 18 103
use INVX1  INVX1_589
timestamp 1693479267
transform 1 0 2980 0 -1 3905
box -2 -3 18 103
use NAND3X1  NAND3X1_272
timestamp 1693479267
transform 1 0 2996 0 -1 3905
box -2 -3 34 103
use NAND3X1  NAND3X1_273
timestamp 1693479267
transform 1 0 3028 0 -1 3905
box -2 -3 34 103
use FILL  FILL_38_5_0
timestamp 1693479267
transform 1 0 3060 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_5_1
timestamp 1693479267
transform 1 0 3068 0 -1 3905
box -2 -3 10 103
use NAND3X1  NAND3X1_274
timestamp 1693479267
transform 1 0 3076 0 -1 3905
box -2 -3 34 103
use NAND3X1  NAND3X1_275
timestamp 1693479267
transform 1 0 3108 0 -1 3905
box -2 -3 34 103
use INVX1  INVX1_517
timestamp 1693479267
transform -1 0 3156 0 -1 3905
box -2 -3 18 103
use INVX1  INVX1_590
timestamp 1693479267
transform 1 0 3156 0 -1 3905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_113
timestamp 1693479267
transform -1 0 3268 0 -1 3905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_116
timestamp 1693479267
transform 1 0 3268 0 -1 3905
box -2 -3 98 103
use INVX1  INVX1_99
timestamp 1693479267
transform 1 0 3364 0 -1 3905
box -2 -3 18 103
use NAND2X1  NAND2X1_99
timestamp 1693479267
transform 1 0 3380 0 -1 3905
box -2 -3 26 103
use NOR2X1  NOR2X1_3
timestamp 1693479267
transform -1 0 3428 0 -1 3905
box -2 -3 26 103
use AND2X2  AND2X2_98
timestamp 1693479267
transform 1 0 3428 0 -1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_114
timestamp 1693479267
transform -1 0 3556 0 -1 3905
box -2 -3 98 103
use FILL  FILL_38_6_0
timestamp 1693479267
transform 1 0 3556 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_6_1
timestamp 1693479267
transform 1 0 3564 0 -1 3905
box -2 -3 10 103
use OAI21X1  OAI21X1_950
timestamp 1693479267
transform 1 0 3572 0 -1 3905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_62
timestamp 1693479267
transform -1 0 3676 0 -1 3905
box -2 -3 74 103
use NOR2X1  NOR2X1_468
timestamp 1693479267
transform -1 0 3700 0 -1 3905
box -2 -3 26 103
use NOR2X1  NOR2X1_470
timestamp 1693479267
transform 1 0 3700 0 -1 3905
box -2 -3 26 103
use AND2X2  AND2X2_99
timestamp 1693479267
transform 1 0 3724 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1012
timestamp 1693479267
transform -1 0 3788 0 -1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_483
timestamp 1693479267
transform 1 0 3788 0 -1 3905
box -2 -3 26 103
use OAI21X1  OAI21X1_978
timestamp 1693479267
transform -1 0 3844 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1067
timestamp 1693479267
transform 1 0 3844 0 -1 3905
box -2 -3 34 103
use INVX1  INVX1_757
timestamp 1693479267
transform 1 0 3876 0 -1 3905
box -2 -3 18 103
use OAI21X1  OAI21X1_1064
timestamp 1693479267
transform -1 0 3924 0 -1 3905
box -2 -3 34 103
use INVX2  INVX2_87
timestamp 1693479267
transform -1 0 3940 0 -1 3905
box -2 -3 18 103
use INVX1  INVX1_753
timestamp 1693479267
transform 1 0 3940 0 -1 3905
box -2 -3 18 103
use NOR2X1  NOR2X1_484
timestamp 1693479267
transform 1 0 3956 0 -1 3905
box -2 -3 26 103
use OAI21X1  OAI21X1_1062
timestamp 1693479267
transform 1 0 3980 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1063
timestamp 1693479267
transform -1 0 4044 0 -1 3905
box -2 -3 34 103
use INVX1  INVX1_754
timestamp 1693479267
transform 1 0 4044 0 -1 3905
box -2 -3 18 103
use NAND2X1  NAND2X1_1020
timestamp 1693479267
transform 1 0 4060 0 -1 3905
box -2 -3 26 103
use FILL  FILL_38_7_0
timestamp 1693479267
transform 1 0 4084 0 -1 3905
box -2 -3 10 103
use FILL  FILL_38_7_1
timestamp 1693479267
transform 1 0 4092 0 -1 3905
box -2 -3 10 103
use OAI21X1  OAI21X1_1031
timestamp 1693479267
transform 1 0 4100 0 -1 3905
box -2 -3 34 103
use AOI22X1  AOI22X1_150
timestamp 1693479267
transform -1 0 4172 0 -1 3905
box -2 -3 42 103
use BUFX4  BUFX4_105
timestamp 1693479267
transform -1 0 4204 0 -1 3905
box -2 -3 34 103
use AOI22X1  AOI22X1_151
timestamp 1693479267
transform -1 0 4244 0 -1 3905
box -2 -3 42 103
use OAI21X1  OAI21X1_1044
timestamp 1693479267
transform -1 0 4276 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1035
timestamp 1693479267
transform -1 0 4308 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1049
timestamp 1693479267
transform -1 0 4340 0 -1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1046
timestamp 1693479267
transform 1 0 4340 0 -1 3905
box -2 -3 34 103
use BUFX4  BUFX4_107
timestamp 1693479267
transform 1 0 4372 0 -1 3905
box -2 -3 34 103
use BUFX4  BUFX4_172
timestamp 1693479267
transform 1 0 4404 0 -1 3905
box -2 -3 34 103
use INVX1  INVX1_736
timestamp 1693479267
transform -1 0 4452 0 -1 3905
box -2 -3 18 103
use AOI22X1  AOI22X1_153
timestamp 1693479267
transform -1 0 4492 0 -1 3905
box -2 -3 42 103
use AOI22X1  AOI22X1_164
timestamp 1693479267
transform 1 0 4492 0 -1 3905
box -2 -3 42 103
use AOI22X1  AOI22X1_157
timestamp 1693479267
transform -1 0 4572 0 -1 3905
box -2 -3 42 103
use FILL  FILL_39_1
timestamp 1693479267
transform -1 0 4580 0 -1 3905
box -2 -3 10 103
use FILL  FILL_39_2
timestamp 1693479267
transform -1 0 4588 0 -1 3905
box -2 -3 10 103
use FILL  FILL_39_3
timestamp 1693479267
transform -1 0 4596 0 -1 3905
box -2 -3 10 103
use FILL  FILL_39_4
timestamp 1693479267
transform -1 0 4604 0 -1 3905
box -2 -3 10 103
use INVX1  INVX1_174
timestamp 1693479267
transform 1 0 4 0 1 3905
box -2 -3 18 103
use NOR3X1  NOR3X1_33
timestamp 1693479267
transform 1 0 20 0 1 3905
box -2 -3 66 103
use INVX1  INVX1_164
timestamp 1693479267
transform 1 0 84 0 1 3905
box -2 -3 18 103
use NOR3X1  NOR3X1_23
timestamp 1693479267
transform 1 0 100 0 1 3905
box -2 -3 66 103
use NOR3X1  NOR3X1_17
timestamp 1693479267
transform -1 0 228 0 1 3905
box -2 -3 66 103
use INVX2  INVX2_3
timestamp 1693479267
transform 1 0 228 0 1 3905
box -2 -3 18 103
use OAI22X1  OAI22X1_5
timestamp 1693479267
transform 1 0 244 0 1 3905
box -2 -3 42 103
use INVX2  INVX2_2
timestamp 1693479267
transform -1 0 300 0 1 3905
box -2 -3 18 103
use AOI22X1  AOI22X1_7
timestamp 1693479267
transform 1 0 300 0 1 3905
box -2 -3 42 103
use INVX1  INVX1_135
timestamp 1693479267
transform 1 0 340 0 1 3905
box -2 -3 18 103
use AOI22X1  AOI22X1_4
timestamp 1693479267
transform -1 0 396 0 1 3905
box -2 -3 42 103
use INVX2  INVX2_1
timestamp 1693479267
transform -1 0 412 0 1 3905
box -2 -3 18 103
use NAND2X1  NAND2X1_101
timestamp 1693479267
transform 1 0 412 0 1 3905
box -2 -3 26 103
use OAI22X1  OAI22X1_1
timestamp 1693479267
transform -1 0 476 0 1 3905
box -2 -3 42 103
use AOI22X1  AOI22X1_2
timestamp 1693479267
transform 1 0 476 0 1 3905
box -2 -3 42 103
use FILL  FILL_39_0_0
timestamp 1693479267
transform -1 0 524 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_0_1
timestamp 1693479267
transform -1 0 532 0 1 3905
box -2 -3 10 103
use INVX1  INVX1_133
timestamp 1693479267
transform -1 0 548 0 1 3905
box -2 -3 18 103
use XNOR2X1  XNOR2X1_4
timestamp 1693479267
transform -1 0 604 0 1 3905
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_155
timestamp 1693479267
transform 1 0 604 0 1 3905
box -2 -3 98 103
use NOR2X1  NOR2X1_400
timestamp 1693479267
transform 1 0 700 0 1 3905
box -2 -3 26 103
use NAND3X1  NAND3X1_187
timestamp 1693479267
transform -1 0 756 0 1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_700
timestamp 1693479267
transform 1 0 756 0 1 3905
box -2 -3 26 103
use INVX1  INVX1_497
timestamp 1693479267
transform -1 0 796 0 1 3905
box -2 -3 18 103
use INVX1  INVX1_570
timestamp 1693479267
transform 1 0 796 0 1 3905
box -2 -3 18 103
use NAND2X1  NAND2X1_810
timestamp 1693479267
transform 1 0 812 0 1 3905
box -2 -3 26 103
use NAND2X1  NAND2X1_701
timestamp 1693479267
transform 1 0 836 0 1 3905
box -2 -3 26 103
use NAND2X1  NAND2X1_811
timestamp 1693479267
transform 1 0 860 0 1 3905
box -2 -3 26 103
use INVX2  INVX2_77
timestamp 1693479267
transform -1 0 900 0 1 3905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_157
timestamp 1693479267
transform 1 0 900 0 1 3905
box -2 -3 98 103
use FILL  FILL_39_1_0
timestamp 1693479267
transform -1 0 1004 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_1_1
timestamp 1693479267
transform -1 0 1012 0 1 3905
box -2 -3 10 103
use BUFX4  BUFX4_1
timestamp 1693479267
transform -1 0 1044 0 1 3905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_43
timestamp 1693479267
transform -1 0 1116 0 1 3905
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_64
timestamp 1693479267
transform -1 0 1212 0 1 3905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_149
timestamp 1693479267
transform -1 0 1308 0 1 3905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_66
timestamp 1693479267
transform -1 0 1404 0 1 3905
box -2 -3 98 103
use INVX1  INVX1_119
timestamp 1693479267
transform 1 0 1404 0 1 3905
box -2 -3 18 103
use CLKBUF1  CLKBUF1_61
timestamp 1693479267
transform -1 0 1492 0 1 3905
box -2 -3 74 103
use INVX1  INVX1_202
timestamp 1693479267
transform -1 0 1508 0 1 3905
box -2 -3 18 103
use INVX1  INVX1_117
timestamp 1693479267
transform 1 0 1508 0 1 3905
box -2 -3 18 103
use FILL  FILL_39_2_0
timestamp 1693479267
transform -1 0 1532 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_2_1
timestamp 1693479267
transform -1 0 1540 0 1 3905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_89
timestamp 1693479267
transform -1 0 1636 0 1 3905
box -2 -3 98 103
use BUFX4  BUFX4_99
timestamp 1693479267
transform -1 0 1668 0 1 3905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_111
timestamp 1693479267
transform 1 0 1668 0 1 3905
box -2 -3 98 103
use OAI21X1  OAI21X1_134
timestamp 1693479267
transform -1 0 1796 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_138
timestamp 1693479267
transform -1 0 1828 0 1 3905
box -2 -3 34 103
use OR2X2  OR2X2_2
timestamp 1693479267
transform 1 0 1828 0 1 3905
box -2 -3 34 103
use BUFX4  BUFX4_271
timestamp 1693479267
transform -1 0 1892 0 1 3905
box -2 -3 34 103
use BUFX4  BUFX4_191
timestamp 1693479267
transform -1 0 1924 0 1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_886
timestamp 1693479267
transform -1 0 1948 0 1 3905
box -2 -3 26 103
use INVX1  INVX1_620
timestamp 1693479267
transform -1 0 1964 0 1 3905
box -2 -3 18 103
use NAND3X1  NAND3X1_299
timestamp 1693479267
transform -1 0 1996 0 1 3905
box -2 -3 34 103
use BUFX4  BUFX4_2
timestamp 1693479267
transform 1 0 1996 0 1 3905
box -2 -3 34 103
use FILL  FILL_39_3_0
timestamp 1693479267
transform 1 0 2028 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_3_1
timestamp 1693479267
transform 1 0 2036 0 1 3905
box -2 -3 10 103
use BUFX4  BUFX4_201
timestamp 1693479267
transform 1 0 2044 0 1 3905
box -2 -3 34 103
use INVX1  INVX1_551
timestamp 1693479267
transform 1 0 2076 0 1 3905
box -2 -3 18 103
use INVX1  INVX1_624
timestamp 1693479267
transform 1 0 2092 0 1 3905
box -2 -3 18 103
use NAND2X1  NAND2X1_892
timestamp 1693479267
transform 1 0 2108 0 1 3905
box -2 -3 26 103
use NAND2X1  NAND2X1_782
timestamp 1693479267
transform 1 0 2132 0 1 3905
box -2 -3 26 103
use BUFX4  BUFX4_123
timestamp 1693479267
transform -1 0 2188 0 1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_835
timestamp 1693479267
transform 1 0 2188 0 1 3905
box -2 -3 26 103
use BUFX4  BUFX4_102
timestamp 1693479267
transform 1 0 2212 0 1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_862
timestamp 1693479267
transform -1 0 2268 0 1 3905
box -2 -3 26 103
use INVX1  INVX1_604
timestamp 1693479267
transform -1 0 2284 0 1 3905
box -2 -3 18 103
use INVX1  INVX1_531
timestamp 1693479267
transform 1 0 2284 0 1 3905
box -2 -3 18 103
use NAND2X1  NAND2X1_752
timestamp 1693479267
transform 1 0 2300 0 1 3905
box -2 -3 26 103
use INVX1  INVX1_546
timestamp 1693479267
transform 1 0 2324 0 1 3905
box -2 -3 18 103
use INVX1  INVX1_619
timestamp 1693479267
transform 1 0 2340 0 1 3905
box -2 -3 18 103
use BUFX4  BUFX4_202
timestamp 1693479267
transform 1 0 2356 0 1 3905
box -2 -3 34 103
use BUFX4  BUFX4_205
timestamp 1693479267
transform 1 0 2388 0 1 3905
box -2 -3 34 103
use BUFX4  BUFX4_100
timestamp 1693479267
transform 1 0 2420 0 1 3905
box -2 -3 34 103
use BUFX4  BUFX4_101
timestamp 1693479267
transform 1 0 2452 0 1 3905
box -2 -3 34 103
use BUFX4  BUFX4_168
timestamp 1693479267
transform -1 0 2516 0 1 3905
box -2 -3 34 103
use BUFX4  BUFX4_165
timestamp 1693479267
transform 1 0 2516 0 1 3905
box -2 -3 34 103
use FILL  FILL_39_4_0
timestamp 1693479267
transform 1 0 2548 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_4_1
timestamp 1693479267
transform 1 0 2556 0 1 3905
box -2 -3 10 103
use BUFX4  BUFX4_166
timestamp 1693479267
transform 1 0 2564 0 1 3905
box -2 -3 34 103
use NAND3X1  NAND3X1_302
timestamp 1693479267
transform 1 0 2596 0 1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_746
timestamp 1693479267
transform -1 0 2652 0 1 3905
box -2 -3 26 103
use INVX1  INVX1_527
timestamp 1693479267
transform -1 0 2668 0 1 3905
box -2 -3 18 103
use NAND2X1  NAND2X1_728
timestamp 1693479267
transform -1 0 2692 0 1 3905
box -2 -3 26 103
use NAND3X1  NAND3X1_282
timestamp 1693479267
transform 1 0 2692 0 1 3905
box -2 -3 34 103
use INVX1  INVX1_600
timestamp 1693479267
transform 1 0 2724 0 1 3905
box -2 -3 18 103
use NAND2X1  NAND2X1_743
timestamp 1693479267
transform -1 0 2764 0 1 3905
box -2 -3 26 103
use INVX1  INVX1_525
timestamp 1693479267
transform -1 0 2780 0 1 3905
box -2 -3 18 103
use NAND2X1  NAND2X1_856
timestamp 1693479267
transform 1 0 2780 0 1 3905
box -2 -3 26 103
use INVX1  INVX1_598
timestamp 1693479267
transform 1 0 2804 0 1 3905
box -2 -3 18 103
use INVX1  INVX1_515
timestamp 1693479267
transform -1 0 2836 0 1 3905
box -2 -3 18 103
use NAND2X1  NAND2X1_853
timestamp 1693479267
transform 1 0 2836 0 1 3905
box -2 -3 26 103
use INVX1  INVX1_588
timestamp 1693479267
transform 1 0 2860 0 1 3905
box -2 -3 18 103
use NAND2X1  NAND2X1_838
timestamp 1693479267
transform 1 0 2876 0 1 3905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_112
timestamp 1693479267
transform 1 0 2900 0 1 3905
box -2 -3 98 103
use BUFX4  BUFX4_119
timestamp 1693479267
transform -1 0 3028 0 1 3905
box -2 -3 34 103
use FILL  FILL_39_5_0
timestamp 1693479267
transform -1 0 3036 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_5_1
timestamp 1693479267
transform -1 0 3044 0 1 3905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_3
timestamp 1693479267
transform -1 0 3140 0 1 3905
box -2 -3 98 103
use NAND2X1  NAND2X1_841
timestamp 1693479267
transform -1 0 3164 0 1 3905
box -2 -3 26 103
use CLKBUF1  CLKBUF1_60
timestamp 1693479267
transform -1 0 3236 0 1 3905
box -2 -3 74 103
use NAND2X1  NAND2X1_997
timestamp 1693479267
transform 1 0 3236 0 1 3905
box -2 -3 26 103
use NOR3X1  NOR3X1_75
timestamp 1693479267
transform -1 0 3324 0 1 3905
box -2 -3 66 103
use NAND3X1  NAND3X1_351
timestamp 1693479267
transform -1 0 3356 0 1 3905
box -2 -3 34 103
use INVX2  INVX2_88
timestamp 1693479267
transform 1 0 3356 0 1 3905
box -2 -3 18 103
use NAND3X1  NAND3X1_348
timestamp 1693479267
transform 1 0 3372 0 1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_999
timestamp 1693479267
transform 1 0 3404 0 1 3905
box -2 -3 26 103
use NAND3X1  NAND3X1_344
timestamp 1693479267
transform 1 0 3428 0 1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_487
timestamp 1693479267
transform 1 0 3460 0 1 3905
box -2 -3 26 103
use BUFX4  BUFX4_11
timestamp 1693479267
transform -1 0 3516 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1059
timestamp 1693479267
transform 1 0 3516 0 1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_1019
timestamp 1693479267
transform 1 0 3548 0 1 3905
box -2 -3 26 103
use FILL  FILL_39_6_0
timestamp 1693479267
transform -1 0 3580 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_6_1
timestamp 1693479267
transform -1 0 3588 0 1 3905
box -2 -3 10 103
use OAI21X1  OAI21X1_1069
timestamp 1693479267
transform -1 0 3620 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1060
timestamp 1693479267
transform 1 0 3620 0 1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_488
timestamp 1693479267
transform -1 0 3676 0 1 3905
box -2 -3 26 103
use OR2X2  OR2X2_70
timestamp 1693479267
transform -1 0 3708 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1061
timestamp 1693479267
transform -1 0 3740 0 1 3905
box -2 -3 34 103
use INVX8  INVX8_16
timestamp 1693479267
transform -1 0 3780 0 1 3905
box -2 -3 42 103
use AND2X2  AND2X2_101
timestamp 1693479267
transform -1 0 3812 0 1 3905
box -2 -3 34 103
use NOR2X1  NOR2X1_472
timestamp 1693479267
transform -1 0 3836 0 1 3905
box -2 -3 26 103
use NOR2X1  NOR2X1_477
timestamp 1693479267
transform 1 0 3836 0 1 3905
box -2 -3 26 103
use OAI22X1  OAI22X1_60
timestamp 1693479267
transform -1 0 3900 0 1 3905
box -2 -3 42 103
use NOR2X1  NOR2X1_485
timestamp 1693479267
transform 1 0 3900 0 1 3905
box -2 -3 26 103
use AOI21X1  AOI21X1_267
timestamp 1693479267
transform 1 0 3924 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_1014
timestamp 1693479267
transform 1 0 3956 0 1 3905
box -2 -3 34 103
use INVX2  INVX2_93
timestamp 1693479267
transform 1 0 3988 0 1 3905
box -2 -3 18 103
use BUFX4  BUFX4_10
timestamp 1693479267
transform 1 0 4004 0 1 3905
box -2 -3 34 103
use INVX1  INVX1_755
timestamp 1693479267
transform 1 0 4036 0 1 3905
box -2 -3 18 103
use OAI21X1  OAI21X1_1034
timestamp 1693479267
transform 1 0 4052 0 1 3905
box -2 -3 34 103
use FILL  FILL_39_7_0
timestamp 1693479267
transform 1 0 4084 0 1 3905
box -2 -3 10 103
use FILL  FILL_39_7_1
timestamp 1693479267
transform 1 0 4092 0 1 3905
box -2 -3 10 103
use BUFX4  BUFX4_171
timestamp 1693479267
transform 1 0 4100 0 1 3905
box -2 -3 34 103
use BUFX4  BUFX4_69
timestamp 1693479267
transform 1 0 4132 0 1 3905
box -2 -3 34 103
use AOI22X1  AOI22X1_160
timestamp 1693479267
transform 1 0 4164 0 1 3905
box -2 -3 42 103
use AOI22X1  AOI22X1_162
timestamp 1693479267
transform 1 0 4204 0 1 3905
box -2 -3 42 103
use AOI22X1  AOI22X1_165
timestamp 1693479267
transform 1 0 4244 0 1 3905
box -2 -3 42 103
use AOI22X1  AOI22X1_163
timestamp 1693479267
transform -1 0 4324 0 1 3905
box -2 -3 42 103
use INVX1  INVX1_738
timestamp 1693479267
transform -1 0 4340 0 1 3905
box -2 -3 18 103
use OAI21X1  OAI21X1_996
timestamp 1693479267
transform -1 0 4372 0 1 3905
box -2 -3 34 103
use AOI21X1  AOI21X1_262
timestamp 1693479267
transform 1 0 4372 0 1 3905
box -2 -3 34 103
use OAI21X1  OAI21X1_998
timestamp 1693479267
transform 1 0 4404 0 1 3905
box -2 -3 34 103
use OAI22X1  OAI22X1_57
timestamp 1693479267
transform -1 0 4476 0 1 3905
box -2 -3 42 103
use INVX1  INVX1_746
timestamp 1693479267
transform -1 0 4492 0 1 3905
box -2 -3 18 103
use AOI22X1  AOI22X1_141
timestamp 1693479267
transform 1 0 4492 0 1 3905
box -2 -3 42 103
use OAI21X1  OAI21X1_997
timestamp 1693479267
transform 1 0 4532 0 1 3905
box -2 -3 34 103
use NAND2X1  NAND2X1_1015
timestamp 1693479267
transform -1 0 4588 0 1 3905
box -2 -3 26 103
use INVX1  INVX1_744
timestamp 1693479267
transform -1 0 4604 0 1 3905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_426
timestamp 1693479267
transform 1 0 4 0 -1 4105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_39
timestamp 1693479267
transform -1 0 172 0 -1 4105
box -2 -3 74 103
use INVX1  INVX1_137
timestamp 1693479267
transform 1 0 172 0 -1 4105
box -2 -3 18 103
use OAI22X1  OAI22X1_4
timestamp 1693479267
transform -1 0 228 0 -1 4105
box -2 -3 42 103
use AOI22X1  AOI22X1_6
timestamp 1693479267
transform -1 0 268 0 -1 4105
box -2 -3 42 103
use AOI22X1  AOI22X1_1
timestamp 1693479267
transform 1 0 268 0 -1 4105
box -2 -3 42 103
use INVX1  INVX1_136
timestamp 1693479267
transform 1 0 308 0 -1 4105
box -2 -3 18 103
use AOI22X1  AOI22X1_5
timestamp 1693479267
transform -1 0 364 0 -1 4105
box -2 -3 42 103
use NAND3X1  NAND3X1_3
timestamp 1693479267
transform 1 0 364 0 -1 4105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_2
timestamp 1693479267
transform 1 0 396 0 -1 4105
box -2 -3 58 103
use NAND3X1  NAND3X1_2
timestamp 1693479267
transform -1 0 484 0 -1 4105
box -2 -3 34 103
use FILL  FILL_40_0_0
timestamp 1693479267
transform 1 0 484 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_0_1
timestamp 1693479267
transform 1 0 492 0 -1 4105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_152
timestamp 1693479267
transform 1 0 500 0 -1 4105
box -2 -3 98 103
use NAND3X1  NAND3X1_186
timestamp 1693479267
transform 1 0 596 0 -1 4105
box -2 -3 34 103
use BUFX2  BUFX2_90
timestamp 1693479267
transform 1 0 628 0 -1 4105
box -2 -3 26 103
use NAND2X1  NAND2X1_807
timestamp 1693479267
transform 1 0 652 0 -1 4105
box -2 -3 26 103
use NAND3X1  NAND3X1_256
timestamp 1693479267
transform 1 0 676 0 -1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_808
timestamp 1693479267
transform -1 0 732 0 -1 4105
box -2 -3 26 103
use AOI21X1  AOI21X1_227
timestamp 1693479267
transform -1 0 764 0 -1 4105
box -2 -3 34 103
use INVX1  INVX1_568
timestamp 1693479267
transform -1 0 780 0 -1 4105
box -2 -3 18 103
use NAND2X1  NAND2X1_818
timestamp 1693479267
transform -1 0 804 0 -1 4105
box -2 -3 26 103
use NAND2X1  NAND2X1_819
timestamp 1693479267
transform -1 0 828 0 -1 4105
box -2 -3 26 103
use NAND2X1  NAND2X1_817
timestamp 1693479267
transform 1 0 828 0 -1 4105
box -2 -3 26 103
use NAND3X1  NAND3X1_259
timestamp 1693479267
transform 1 0 852 0 -1 4105
box -2 -3 34 103
use NOR2X1  NOR2X1_408
timestamp 1693479267
transform -1 0 908 0 -1 4105
box -2 -3 26 103
use OAI22X1  OAI22X1_48
timestamp 1693479267
transform 1 0 908 0 -1 4105
box -2 -3 42 103
use AOI21X1  AOI21X1_228
timestamp 1693479267
transform 1 0 948 0 -1 4105
box -2 -3 34 103
use INVX1  INVX1_575
timestamp 1693479267
transform -1 0 996 0 -1 4105
box -2 -3 18 103
use INVX1  INVX1_577
timestamp 1693479267
transform -1 0 1012 0 -1 4105
box -2 -3 18 103
use FILL  FILL_40_1_0
timestamp 1693479267
transform 1 0 1012 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_1_1
timestamp 1693479267
transform 1 0 1020 0 -1 4105
box -2 -3 10 103
use INVX2  INVX2_74
timestamp 1693479267
transform 1 0 1028 0 -1 4105
box -2 -3 18 103
use NOR2X1  NOR2X1_407
timestamp 1693479267
transform -1 0 1068 0 -1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_873
timestamp 1693479267
transform -1 0 1100 0 -1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_36
timestamp 1693479267
transform 1 0 1100 0 -1 4105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_37
timestamp 1693479267
transform 1 0 1196 0 -1 4105
box -2 -3 98 103
use NAND3X1  NAND3X1_258
timestamp 1693479267
transform -1 0 1324 0 -1 4105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_51
timestamp 1693479267
transform -1 0 1396 0 -1 4105
box -2 -3 74 103
use BUFX4  BUFX4_255
timestamp 1693479267
transform 1 0 1396 0 -1 4105
box -2 -3 34 103
use BUFX4  BUFX4_143
timestamp 1693479267
transform 1 0 1428 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_204
timestamp 1693479267
transform 1 0 1460 0 -1 4105
box -2 -3 34 103
use AOI22X1  AOI22X1_19
timestamp 1693479267
transform -1 0 1532 0 -1 4105
box -2 -3 42 103
use FILL  FILL_40_2_0
timestamp 1693479267
transform -1 0 1540 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_2_1
timestamp 1693479267
transform -1 0 1548 0 -1 4105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_107
timestamp 1693479267
transform -1 0 1644 0 -1 4105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_57
timestamp 1693479267
transform -1 0 1740 0 -1 4105
box -2 -3 98 103
use OAI21X1  OAI21X1_155
timestamp 1693479267
transform -1 0 1772 0 -1 4105
box -2 -3 34 103
use INVX1  INVX1_110
timestamp 1693479267
transform 1 0 1772 0 -1 4105
box -2 -3 18 103
use OAI21X1  OAI21X1_120
timestamp 1693479267
transform 1 0 1788 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_119
timestamp 1693479267
transform -1 0 1852 0 -1 4105
box -2 -3 34 103
use BUFX4  BUFX4_186
timestamp 1693479267
transform -1 0 1884 0 -1 4105
box -2 -3 34 103
use BUFX4  BUFX4_194
timestamp 1693479267
transform -1 0 1916 0 -1 4105
box -2 -3 34 103
use BUFX4  BUFX4_167
timestamp 1693479267
transform 1 0 1916 0 -1 4105
box -2 -3 34 103
use NAND3X1  NAND3X1_298
timestamp 1693479267
transform -1 0 1980 0 -1 4105
box -2 -3 34 103
use INVX1  INVX1_615
timestamp 1693479267
transform -1 0 1996 0 -1 4105
box -2 -3 18 103
use NAND3X1  NAND3X1_270
timestamp 1693479267
transform -1 0 2028 0 -1 4105
box -2 -3 34 103
use FILL  FILL_40_3_0
timestamp 1693479267
transform -1 0 2036 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_3_1
timestamp 1693479267
transform -1 0 2044 0 -1 4105
box -2 -3 10 103
use INVX1  INVX1_587
timestamp 1693479267
transform -1 0 2060 0 -1 4105
box -2 -3 18 103
use BUFX4  BUFX4_221
timestamp 1693479267
transform 1 0 2060 0 -1 4105
box -2 -3 34 103
use NAND3X1  NAND3X1_201
timestamp 1693479267
transform -1 0 2124 0 -1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_725
timestamp 1693479267
transform -1 0 2148 0 -1 4105
box -2 -3 26 103
use INVX1  INVX1_513
timestamp 1693479267
transform -1 0 2164 0 -1 4105
box -2 -3 18 103
use INVX1  INVX1_586
timestamp 1693479267
transform 1 0 2164 0 -1 4105
box -2 -3 18 103
use NAND3X1  NAND3X1_223
timestamp 1693479267
transform 1 0 2180 0 -1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_758
timestamp 1693479267
transform -1 0 2236 0 -1 4105
box -2 -3 26 103
use INVX1  INVX1_535
timestamp 1693479267
transform -1 0 2252 0 -1 4105
box -2 -3 18 103
use NAND3X1  NAND3X1_227
timestamp 1693479267
transform 1 0 2252 0 -1 4105
box -2 -3 34 103
use BUFX4  BUFX4_222
timestamp 1693479267
transform 1 0 2284 0 -1 4105
box -2 -3 34 103
use NAND3X1  NAND3X1_232
timestamp 1693479267
transform -1 0 2348 0 -1 4105
box -2 -3 34 103
use NAND3X1  NAND3X1_233
timestamp 1693479267
transform 1 0 2348 0 -1 4105
box -2 -3 34 103
use INVX1  INVX1_560
timestamp 1693479267
transform 1 0 2380 0 -1 4105
box -2 -3 18 103
use NAND3X1  NAND3X1_246
timestamp 1693479267
transform 1 0 2396 0 -1 4105
box -2 -3 34 103
use NAND3X1  NAND3X1_212
timestamp 1693479267
transform -1 0 2460 0 -1 4105
box -2 -3 34 103
use INVX1  INVX1_526
timestamp 1693479267
transform -1 0 2476 0 -1 4105
box -2 -3 18 103
use NAND3X1  NAND3X1_293
timestamp 1693479267
transform -1 0 2508 0 -1 4105
box -2 -3 34 103
use BUFX4  BUFX4_164
timestamp 1693479267
transform -1 0 2540 0 -1 4105
box -2 -3 34 103
use FILL  FILL_40_4_0
timestamp 1693479267
transform 1 0 2540 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_4_1
timestamp 1693479267
transform 1 0 2548 0 -1 4105
box -2 -3 10 103
use INVX1  INVX1_633
timestamp 1693479267
transform 1 0 2556 0 -1 4105
box -2 -3 18 103
use NAND3X1  NAND3X1_316
timestamp 1693479267
transform 1 0 2572 0 -1 4105
box -2 -3 34 103
use NAND3X1  NAND3X1_247
timestamp 1693479267
transform -1 0 2636 0 -1 4105
box -2 -3 34 103
use INVX1  INVX1_599
timestamp 1693479267
transform 1 0 2636 0 -1 4105
box -2 -3 18 103
use INVX1  INVX1_632
timestamp 1693479267
transform 1 0 2652 0 -1 4105
box -2 -3 18 103
use BUFX4  BUFX4_122
timestamp 1693479267
transform 1 0 2668 0 -1 4105
box -2 -3 34 103
use NAND3X1  NAND3X1_213
timestamp 1693479267
transform 1 0 2700 0 -1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_883
timestamp 1693479267
transform 1 0 2732 0 -1 4105
box -2 -3 26 103
use NAND2X1  NAND2X1_904
timestamp 1693479267
transform 1 0 2756 0 -1 4105
box -2 -3 26 103
use NAND3X1  NAND3X1_303
timestamp 1693479267
transform -1 0 2812 0 -1 4105
box -2 -3 34 103
use NAND3X1  NAND3X1_317
timestamp 1693479267
transform -1 0 2844 0 -1 4105
box -2 -3 34 103
use BUFX4  BUFX4_96
timestamp 1693479267
transform 1 0 2844 0 -1 4105
box -2 -3 34 103
use NAND3X1  NAND3X1_325
timestamp 1693479267
transform -1 0 2908 0 -1 4105
box -2 -3 34 103
use NAND3X1  NAND3X1_1
timestamp 1693479267
transform 1 0 2908 0 -1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_1
timestamp 1693479267
transform -1 0 3036 0 -1 4105
box -2 -3 98 103
use NOR2X1  NOR2X1_4
timestamp 1693479267
transform -1 0 3060 0 -1 4105
box -2 -3 26 103
use FILL  FILL_40_5_0
timestamp 1693479267
transform -1 0 3068 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_5_1
timestamp 1693479267
transform -1 0 3076 0 -1 4105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_4
timestamp 1693479267
transform -1 0 3172 0 -1 4105
box -2 -3 98 103
use NOR2X1  NOR2X1_466
timestamp 1693479267
transform 1 0 3172 0 -1 4105
box -2 -3 26 103
use INVX1  INVX1_716
timestamp 1693479267
transform 1 0 3196 0 -1 4105
box -2 -3 18 103
use NAND3X1  NAND3X1_347
timestamp 1693479267
transform 1 0 3212 0 -1 4105
box -2 -3 34 103
use AND2X2  AND2X2_100
timestamp 1693479267
transform -1 0 3276 0 -1 4105
box -2 -3 34 103
use NOR2X1  NOR2X1_469
timestamp 1693479267
transform 1 0 3276 0 -1 4105
box -2 -3 26 103
use NAND2X1  NAND2X1_994
timestamp 1693479267
transform -1 0 3324 0 -1 4105
box -2 -3 26 103
use INVX2  INVX2_89
timestamp 1693479267
transform 1 0 3324 0 -1 4105
box -2 -3 18 103
use NOR2X1  NOR2X1_474
timestamp 1693479267
transform -1 0 3364 0 -1 4105
box -2 -3 26 103
use NOR2X1  NOR2X1_471
timestamp 1693479267
transform 1 0 3364 0 -1 4105
box -2 -3 26 103
use NAND2X1  NAND2X1_995
timestamp 1693479267
transform -1 0 3412 0 -1 4105
box -2 -3 26 103
use NOR3X1  NOR3X1_74
timestamp 1693479267
transform -1 0 3476 0 -1 4105
box -2 -3 66 103
use NOR3X1  NOR3X1_77
timestamp 1693479267
transform -1 0 3540 0 -1 4105
box -2 -3 66 103
use INVX2  INVX2_90
timestamp 1693479267
transform -1 0 3556 0 -1 4105
box -2 -3 18 103
use FILL  FILL_40_6_0
timestamp 1693479267
transform -1 0 3564 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_6_1
timestamp 1693479267
transform -1 0 3572 0 -1 4105
box -2 -3 10 103
use OAI21X1  OAI21X1_1057
timestamp 1693479267
transform -1 0 3604 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1068
timestamp 1693479267
transform -1 0 3636 0 -1 4105
box -2 -3 34 103
use INVX1  INVX1_759
timestamp 1693479267
transform -1 0 3652 0 -1 4105
box -2 -3 18 103
use OAI21X1  OAI21X1_946
timestamp 1693479267
transform 1 0 3652 0 -1 4105
box -2 -3 34 103
use NOR2X1  NOR2X1_476
timestamp 1693479267
transform 1 0 3684 0 -1 4105
box -2 -3 26 103
use NAND3X1  NAND3X1_346
timestamp 1693479267
transform -1 0 3740 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_975
timestamp 1693479267
transform 1 0 3740 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1007
timestamp 1693479267
transform 1 0 3772 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_947
timestamp 1693479267
transform 1 0 3804 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1065
timestamp 1693479267
transform -1 0 3868 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1008
timestamp 1693479267
transform 1 0 3868 0 -1 4105
box -2 -3 34 103
use NAND3X1  NAND3X1_358
timestamp 1693479267
transform -1 0 3932 0 -1 4105
box -2 -3 34 103
use NAND3X1  NAND3X1_357
timestamp 1693479267
transform -1 0 3964 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1013
timestamp 1693479267
transform -1 0 3996 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1009
timestamp 1693479267
transform 1 0 3996 0 -1 4105
box -2 -3 34 103
use AOI21X1  AOI21X1_265
timestamp 1693479267
transform 1 0 4028 0 -1 4105
box -2 -3 34 103
use AOI21X1  AOI21X1_266
timestamp 1693479267
transform -1 0 4092 0 -1 4105
box -2 -3 34 103
use FILL  FILL_40_7_0
timestamp 1693479267
transform -1 0 4100 0 -1 4105
box -2 -3 10 103
use FILL  FILL_40_7_1
timestamp 1693479267
transform -1 0 4108 0 -1 4105
box -2 -3 10 103
use OAI21X1  OAI21X1_1033
timestamp 1693479267
transform -1 0 4140 0 -1 4105
box -2 -3 34 103
use OAI22X1  OAI22X1_54
timestamp 1693479267
transform 1 0 4140 0 -1 4105
box -2 -3 42 103
use INVX1  INVX1_737
timestamp 1693479267
transform -1 0 4196 0 -1 4105
box -2 -3 18 103
use AOI21X1  AOI21X1_258
timestamp 1693479267
transform -1 0 4228 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_984
timestamp 1693479267
transform 1 0 4228 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_983
timestamp 1693479267
transform 1 0 4260 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_991
timestamp 1693479267
transform 1 0 4292 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_995
timestamp 1693479267
transform 1 0 4324 0 -1 4105
box -2 -3 34 103
use BUFX4  BUFX4_65
timestamp 1693479267
transform -1 0 4388 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1022
timestamp 1693479267
transform 1 0 4388 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1016
timestamp 1693479267
transform 1 0 4420 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1023
timestamp 1693479267
transform -1 0 4484 0 -1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1048
timestamp 1693479267
transform -1 0 4516 0 -1 4105
box -2 -3 34 103
use INVX1  INVX1_745
timestamp 1693479267
transform -1 0 4532 0 -1 4105
box -2 -3 18 103
use AOI22X1  AOI22X1_147
timestamp 1693479267
transform -1 0 4572 0 -1 4105
box -2 -3 42 103
use OAI21X1  OAI21X1_1024
timestamp 1693479267
transform 1 0 4572 0 -1 4105
box -2 -3 34 103
use INVX1  INVX1_172
timestamp 1693479267
transform 1 0 4 0 1 4105
box -2 -3 18 103
use NOR3X1  NOR3X1_31
timestamp 1693479267
transform -1 0 84 0 1 4105
box -2 -3 66 103
use XOR2X1  XOR2X1_1
timestamp 1693479267
transform -1 0 140 0 1 4105
box -2 -3 58 103
use NOR3X1  NOR3X1_16
timestamp 1693479267
transform -1 0 204 0 1 4105
box -2 -3 66 103
use OAI22X1  OAI22X1_2
timestamp 1693479267
transform -1 0 244 0 1 4105
box -2 -3 42 103
use INVX1  INVX1_134
timestamp 1693479267
transform -1 0 260 0 1 4105
box -2 -3 18 103
use OAI22X1  OAI22X1_3
timestamp 1693479267
transform 1 0 260 0 1 4105
box -2 -3 42 103
use INVX1  INVX1_132
timestamp 1693479267
transform -1 0 316 0 1 4105
box -2 -3 18 103
use AOI22X1  AOI22X1_3
timestamp 1693479267
transform -1 0 356 0 1 4105
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_156
timestamp 1693479267
transform 1 0 356 0 1 4105
box -2 -3 98 103
use OR2X2  OR2X2_51
timestamp 1693479267
transform 1 0 452 0 1 4105
box -2 -3 34 103
use INVX1  INVX1_496
timestamp 1693479267
transform 1 0 484 0 1 4105
box -2 -3 18 103
use FILL  FILL_41_0_0
timestamp 1693479267
transform -1 0 508 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_0_1
timestamp 1693479267
transform -1 0 516 0 1 4105
box -2 -3 10 103
use NAND2X1  NAND2X1_699
timestamp 1693479267
transform -1 0 540 0 1 4105
box -2 -3 26 103
use INVX1  INVX1_495
timestamp 1693479267
transform 1 0 540 0 1 4105
box -2 -3 18 103
use NAND2X1  NAND2X1_697
timestamp 1693479267
transform 1 0 556 0 1 4105
box -2 -3 26 103
use NAND2X1  NAND2X1_709
timestamp 1693479267
transform -1 0 604 0 1 4105
box -2 -3 26 103
use NAND2X1  NAND2X1_698
timestamp 1693479267
transform 1 0 604 0 1 4105
box -2 -3 26 103
use INVX2  INVX2_73
timestamp 1693479267
transform -1 0 644 0 1 4105
box -2 -3 18 103
use INVX1  INVX1_569
timestamp 1693479267
transform 1 0 644 0 1 4105
box -2 -3 18 103
use NAND2X1  NAND2X1_809
timestamp 1693479267
transform -1 0 684 0 1 4105
box -2 -3 26 103
use INVX2  INVX2_78
timestamp 1693479267
transform 1 0 684 0 1 4105
box -2 -3 18 103
use INVX2  INVX2_76
timestamp 1693479267
transform 1 0 700 0 1 4105
box -2 -3 18 103
use OAI22X1  OAI22X1_47
timestamp 1693479267
transform 1 0 716 0 1 4105
box -2 -3 42 103
use INVX1  INVX1_574
timestamp 1693479267
transform -1 0 772 0 1 4105
box -2 -3 18 103
use AOI22X1  AOI22X1_113
timestamp 1693479267
transform 1 0 772 0 1 4105
box -2 -3 42 103
use NAND2X1  NAND2X1_820
timestamp 1693479267
transform -1 0 836 0 1 4105
box -2 -3 26 103
use NAND2X1  NAND2X1_708
timestamp 1693479267
transform 1 0 836 0 1 4105
box -2 -3 26 103
use NAND3X1  NAND3X1_189
timestamp 1693479267
transform -1 0 892 0 1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_707
timestamp 1693479267
transform -1 0 916 0 1 4105
box -2 -3 26 103
use OAI22X1  OAI22X1_46
timestamp 1693479267
transform 1 0 916 0 1 4105
box -2 -3 42 103
use INVX1  INVX1_502
timestamp 1693479267
transform 1 0 956 0 1 4105
box -2 -3 18 103
use AOI21X1  AOI21X1_224
timestamp 1693479267
transform 1 0 972 0 1 4105
box -2 -3 34 103
use FILL  FILL_41_1_0
timestamp 1693479267
transform -1 0 1012 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_1_1
timestamp 1693479267
transform -1 0 1020 0 1 4105
box -2 -3 10 103
use INVX1  INVX1_504
timestamp 1693479267
transform -1 0 1036 0 1 4105
box -2 -3 18 103
use NOR2X1  NOR2X1_402
timestamp 1693479267
transform 1 0 1036 0 1 4105
box -2 -3 26 103
use NAND2X1  NAND2X1_710
timestamp 1693479267
transform 1 0 1060 0 1 4105
box -2 -3 26 103
use INVX1  INVX1_501
timestamp 1693479267
transform 1 0 1084 0 1 4105
box -2 -3 18 103
use AOI22X1  AOI22X1_111
timestamp 1693479267
transform 1 0 1100 0 1 4105
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_75
timestamp 1693479267
transform -1 0 1236 0 1 4105
box -2 -3 98 103
use AOI22X1  AOI22X1_37
timestamp 1693479267
transform 1 0 1236 0 1 4105
box -2 -3 42 103
use AOI22X1  AOI22X1_36
timestamp 1693479267
transform -1 0 1316 0 1 4105
box -2 -3 42 103
use INVX1  INVX1_128
timestamp 1693479267
transform 1 0 1316 0 1 4105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_74
timestamp 1693479267
transform -1 0 1428 0 1 4105
box -2 -3 98 103
use INVX1  INVX1_127
timestamp 1693479267
transform 1 0 1428 0 1 4105
box -2 -3 18 103
use OAI21X1  OAI21X1_222
timestamp 1693479267
transform -1 0 1476 0 1 4105
box -2 -3 34 103
use INVX1  INVX1_220
timestamp 1693479267
transform -1 0 1492 0 1 4105
box -2 -3 18 103
use OAI21X1  OAI21X1_221
timestamp 1693479267
transform -1 0 1524 0 1 4105
box -2 -3 34 103
use FILL  FILL_41_2_0
timestamp 1693479267
transform -1 0 1532 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_2_1
timestamp 1693479267
transform -1 0 1540 0 1 4105
box -2 -3 10 103
use INVX1  INVX1_219
timestamp 1693479267
transform -1 0 1556 0 1 4105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_106
timestamp 1693479267
transform -1 0 1652 0 1 4105
box -2 -3 98 103
use BUFX4  BUFX4_239
timestamp 1693479267
transform -1 0 1684 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_156
timestamp 1693479267
transform 1 0 1684 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_154
timestamp 1693479267
transform 1 0 1716 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_153
timestamp 1693479267
transform -1 0 1780 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_99
timestamp 1693479267
transform 1 0 1780 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_107
timestamp 1693479267
transform 1 0 1812 0 1 4105
box -2 -3 34 103
use BUFX4  BUFX4_97
timestamp 1693479267
transform 1 0 1844 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_159
timestamp 1693479267
transform 1 0 1876 0 1 4105
box -2 -3 34 103
use BUFX4  BUFX4_36
timestamp 1693479267
transform 1 0 1908 0 1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_877
timestamp 1693479267
transform -1 0 1964 0 1 4105
box -2 -3 26 103
use INVX1  INVX1_556
timestamp 1693479267
transform 1 0 1964 0 1 4105
box -2 -3 18 103
use INVX1  INVX1_542
timestamp 1693479267
transform 1 0 1980 0 1 4105
box -2 -3 18 103
use NAND3X1  NAND3X1_228
timestamp 1693479267
transform 1 0 1996 0 1 4105
box -2 -3 34 103
use FILL  FILL_41_3_0
timestamp 1693479267
transform -1 0 2036 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_3_1
timestamp 1693479267
transform -1 0 2044 0 1 4105
box -2 -3 10 103
use NAND3X1  NAND3X1_222
timestamp 1693479267
transform -1 0 2076 0 1 4105
box -2 -3 34 103
use INVX1  INVX1_536
timestamp 1693479267
transform -1 0 2092 0 1 4105
box -2 -3 18 103
use BUFX4  BUFX4_208
timestamp 1693479267
transform 1 0 2092 0 1 4105
box -2 -3 34 103
use INVX1  INVX1_609
timestamp 1693479267
transform 1 0 2124 0 1 4105
box -2 -3 18 103
use INVX1  INVX1_540
timestamp 1693479267
transform 1 0 2140 0 1 4105
box -2 -3 18 103
use NAND3X1  NAND3X1_226
timestamp 1693479267
transform 1 0 2156 0 1 4105
box -2 -3 34 103
use INVX1  INVX1_613
timestamp 1693479267
transform 1 0 2188 0 1 4105
box -2 -3 18 103
use NAND2X1  NAND2X1_898
timestamp 1693479267
transform 1 0 2204 0 1 4105
box -2 -3 26 103
use BUFX4  BUFX4_37
timestamp 1693479267
transform 1 0 2228 0 1 4105
box -2 -3 34 103
use INVX1  INVX1_608
timestamp 1693479267
transform 1 0 2260 0 1 4105
box -2 -3 18 103
use NAND2X1  NAND2X1_764
timestamp 1693479267
transform -1 0 2300 0 1 4105
box -2 -3 26 103
use INVX1  INVX1_539
timestamp 1693479267
transform -1 0 2316 0 1 4105
box -2 -3 18 103
use NAND3X1  NAND3X1_248
timestamp 1693479267
transform -1 0 2348 0 1 4105
box -2 -3 34 103
use INVX1  INVX1_562
timestamp 1693479267
transform -1 0 2364 0 1 4105
box -2 -3 18 103
use INVX1  INVX1_612
timestamp 1693479267
transform 1 0 2364 0 1 4105
box -2 -3 18 103
use NAND2X1  NAND2X1_874
timestamp 1693479267
transform 1 0 2380 0 1 4105
box -2 -3 26 103
use NAND2X1  NAND2X1_868
timestamp 1693479267
transform 1 0 2404 0 1 4105
box -2 -3 26 103
use NAND3X1  NAND3X1_292
timestamp 1693479267
transform 1 0 2428 0 1 4105
box -2 -3 34 103
use NAND3X1  NAND3X1_296
timestamp 1693479267
transform 1 0 2460 0 1 4105
box -2 -3 34 103
use NAND3X1  NAND3X1_297
timestamp 1693479267
transform -1 0 2524 0 1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_773
timestamp 1693479267
transform -1 0 2548 0 1 4105
box -2 -3 26 103
use FILL  FILL_41_4_0
timestamp 1693479267
transform -1 0 2556 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_4_1
timestamp 1693479267
transform -1 0 2564 0 1 4105
box -2 -3 10 103
use INVX1  INVX1_545
timestamp 1693479267
transform -1 0 2580 0 1 4105
box -2 -3 18 103
use INVX1  INVX1_635
timestamp 1693479267
transform 1 0 2580 0 1 4105
box -2 -3 18 103
use INVX1  INVX1_618
timestamp 1693479267
transform 1 0 2596 0 1 4105
box -2 -3 18 103
use NAND2X1  NAND2X1_794
timestamp 1693479267
transform -1 0 2636 0 1 4105
box -2 -3 26 103
use INVX1  INVX1_559
timestamp 1693479267
transform -1 0 2652 0 1 4105
box -2 -3 18 103
use BUFX4  BUFX4_98
timestamp 1693479267
transform -1 0 2684 0 1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_250
timestamp 1693479267
transform -1 0 2780 0 1 4105
box -2 -3 98 103
use AND2X2  AND2X2_8
timestamp 1693479267
transform -1 0 2812 0 1 4105
box -2 -3 34 103
use AND2X2  AND2X2_6
timestamp 1693479267
transform -1 0 2844 0 1 4105
box -2 -3 34 103
use AND2X2  AND2X2_7
timestamp 1693479267
transform -1 0 2876 0 1 4105
box -2 -3 34 103
use NOR2X1  NOR2X1_10
timestamp 1693479267
transform 1 0 2876 0 1 4105
box -2 -3 26 103
use NOR2X1  NOR2X1_8
timestamp 1693479267
transform 1 0 2900 0 1 4105
box -2 -3 26 103
use NAND2X1  NAND2X1_104
timestamp 1693479267
transform -1 0 2948 0 1 4105
box -2 -3 26 103
use AND2X2  AND2X2_5
timestamp 1693479267
transform -1 0 2980 0 1 4105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_2
timestamp 1693479267
transform -1 0 3076 0 1 4105
box -2 -3 98 103
use FILL  FILL_41_5_0
timestamp 1693479267
transform 1 0 3076 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_5_1
timestamp 1693479267
transform 1 0 3084 0 1 4105
box -2 -3 10 103
use OR2X2  OR2X2_69
timestamp 1693479267
transform 1 0 3092 0 1 4105
box -2 -3 34 103
use NOR3X1  NOR3X1_76
timestamp 1693479267
transform -1 0 3188 0 1 4105
box -2 -3 66 103
use INVX1  INVX1_715
timestamp 1693479267
transform 1 0 3188 0 1 4105
box -2 -3 18 103
use NOR2X1  NOR2X1_467
timestamp 1693479267
transform -1 0 3228 0 1 4105
box -2 -3 26 103
use NAND3X1  NAND3X1_353
timestamp 1693479267
transform -1 0 3260 0 1 4105
box -2 -3 34 103
use NAND3X1  NAND3X1_350
timestamp 1693479267
transform -1 0 3292 0 1 4105
box -2 -3 34 103
use NAND3X1  NAND3X1_356
timestamp 1693479267
transform -1 0 3324 0 1 4105
box -2 -3 34 103
use NAND3X1  NAND3X1_345
timestamp 1693479267
transform 1 0 3324 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_979
timestamp 1693479267
transform -1 0 3388 0 1 4105
box -2 -3 34 103
use NOR3X1  NOR3X1_73
timestamp 1693479267
transform -1 0 3452 0 1 4105
box -2 -3 66 103
use OAI21X1  OAI21X1_942
timestamp 1693479267
transform -1 0 3484 0 1 4105
box -2 -3 34 103
use NOR2X1  NOR2X1_481
timestamp 1693479267
transform 1 0 3484 0 1 4105
box -2 -3 26 103
use NOR2X1  NOR2X1_480
timestamp 1693479267
transform -1 0 3532 0 1 4105
box -2 -3 26 103
use NOR3X1  NOR3X1_78
timestamp 1693479267
transform -1 0 3596 0 1 4105
box -2 -3 66 103
use FILL  FILL_41_6_0
timestamp 1693479267
transform 1 0 3596 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_6_1
timestamp 1693479267
transform 1 0 3604 0 1 4105
box -2 -3 10 103
use AOI21X1  AOI21X1_256
timestamp 1693479267
transform 1 0 3612 0 1 4105
box -2 -3 34 103
use NOR3X1  NOR3X1_79
timestamp 1693479267
transform -1 0 3708 0 1 4105
box -2 -3 66 103
use NOR3X1  NOR3X1_80
timestamp 1693479267
transform 1 0 3708 0 1 4105
box -2 -3 66 103
use OAI21X1  OAI21X1_949
timestamp 1693479267
transform 1 0 3772 0 1 4105
box -2 -3 34 103
use NOR3X1  NOR3X1_81
timestamp 1693479267
transform 1 0 3804 0 1 4105
box -2 -3 66 103
use INVX1  INVX1_734
timestamp 1693479267
transform 1 0 3868 0 1 4105
box -2 -3 18 103
use OAI21X1  OAI21X1_977
timestamp 1693479267
transform 1 0 3884 0 1 4105
box -2 -3 34 103
use INVX4  INVX4_13
timestamp 1693479267
transform -1 0 3940 0 1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_976
timestamp 1693479267
transform 1 0 3940 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_1011
timestamp 1693479267
transform -1 0 4004 0 1 4105
box -2 -3 34 103
use BUFX4  BUFX4_8
timestamp 1693479267
transform -1 0 4036 0 1 4105
box -2 -3 34 103
use NOR2X1  NOR2X1_482
timestamp 1693479267
transform 1 0 4036 0 1 4105
box -2 -3 26 103
use BUFX4  BUFX4_9
timestamp 1693479267
transform 1 0 4060 0 1 4105
box -2 -3 34 103
use FILL  FILL_41_7_0
timestamp 1693479267
transform 1 0 4092 0 1 4105
box -2 -3 10 103
use FILL  FILL_41_7_1
timestamp 1693479267
transform 1 0 4100 0 1 4105
box -2 -3 10 103
use AOI22X1  AOI22X1_138
timestamp 1693479267
transform 1 0 4108 0 1 4105
box -2 -3 42 103
use OAI21X1  OAI21X1_986
timestamp 1693479267
transform -1 0 4180 0 1 4105
box -2 -3 34 103
use NAND2X1  NAND2X1_1012
timestamp 1693479267
transform 1 0 4180 0 1 4105
box -2 -3 26 103
use OAI21X1  OAI21X1_985
timestamp 1693479267
transform -1 0 4236 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_987
timestamp 1693479267
transform -1 0 4268 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_988
timestamp 1693479267
transform -1 0 4300 0 1 4105
box -2 -3 34 103
use AOI21X1  AOI21X1_260
timestamp 1693479267
transform 1 0 4300 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_990
timestamp 1693479267
transform 1 0 4332 0 1 4105
box -2 -3 34 103
use OAI21X1  OAI21X1_989
timestamp 1693479267
transform 1 0 4364 0 1 4105
box -2 -3 34 103
use AOI22X1  AOI22X1_139
timestamp 1693479267
transform -1 0 4436 0 1 4105
box -2 -3 42 103
use NAND2X1  NAND2X1_1013
timestamp 1693479267
transform -1 0 4460 0 1 4105
box -2 -3 26 103
use INVX1  INVX1_740
timestamp 1693479267
transform 1 0 4460 0 1 4105
box -2 -3 18 103
use OAI22X1  OAI22X1_55
timestamp 1693479267
transform -1 0 4516 0 1 4105
box -2 -3 42 103
use OAI21X1  OAI21X1_1017
timestamp 1693479267
transform -1 0 4548 0 1 4105
box -2 -3 34 103
use INVX1  INVX1_747
timestamp 1693479267
transform -1 0 4564 0 1 4105
box -2 -3 18 103
use AOI22X1  AOI22X1_145
timestamp 1693479267
transform -1 0 4604 0 1 4105
box -2 -3 42 103
use INVX1  INVX1_178
timestamp 1693479267
transform 1 0 4 0 -1 4305
box -2 -3 18 103
use NOR3X1  NOR3X1_37
timestamp 1693479267
transform -1 0 84 0 -1 4305
box -2 -3 66 103
use DFFPOSX1  DFFPOSX1_430
timestamp 1693479267
transform 1 0 84 0 -1 4305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_424
timestamp 1693479267
transform 1 0 180 0 -1 4305
box -2 -3 98 103
use BUFX2  BUFX2_91
timestamp 1693479267
transform -1 0 300 0 -1 4305
box -2 -3 26 103
use XOR2X1  XOR2X1_12
timestamp 1693479267
transform 1 0 300 0 -1 4305
box -2 -3 58 103
use NOR2X1  NOR2X1_403
timestamp 1693479267
transform 1 0 356 0 -1 4305
box -2 -3 26 103
use XOR2X1  XOR2X1_16
timestamp 1693479267
transform -1 0 436 0 -1 4305
box -2 -3 58 103
use NOR2X1  NOR2X1_409
timestamp 1693479267
transform 1 0 436 0 -1 4305
box -2 -3 26 103
use FILL  FILL_42_0_0
timestamp 1693479267
transform -1 0 468 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_0_1
timestamp 1693479267
transform -1 0 476 0 -1 4305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_44
timestamp 1693479267
transform -1 0 572 0 -1 4305
box -2 -3 98 103
use NAND2X1  NAND2X1_814
timestamp 1693479267
transform 1 0 572 0 -1 4305
box -2 -3 26 103
use AOI22X1  AOI22X1_112
timestamp 1693479267
transform 1 0 596 0 -1 4305
box -2 -3 42 103
use OR2X2  OR2X2_52
timestamp 1693479267
transform 1 0 636 0 -1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_704
timestamp 1693479267
transform 1 0 668 0 -1 4305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_153
timestamp 1693479267
transform 1 0 692 0 -1 4305
box -2 -3 98 103
use NAND2X1  NAND2X1_805
timestamp 1693479267
transform -1 0 812 0 -1 4305
box -2 -3 26 103
use NAND3X1  NAND3X1_254
timestamp 1693479267
transform 1 0 812 0 -1 4305
box -2 -3 34 103
use INVX2  INVX2_75
timestamp 1693479267
transform 1 0 844 0 -1 4305
box -2 -3 18 103
use NOR2X1  NOR2X1_404
timestamp 1693479267
transform 1 0 860 0 -1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_871
timestamp 1693479267
transform 1 0 884 0 -1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_915
timestamp 1693479267
transform 1 0 916 0 -1 4305
box -2 -3 26 103
use NAND3X1  NAND3X1_324
timestamp 1693479267
transform 1 0 940 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_875
timestamp 1693479267
transform 1 0 972 0 -1 4305
box -2 -3 34 103
use FILL  FILL_42_1_0
timestamp 1693479267
transform -1 0 1012 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_1_1
timestamp 1693479267
transform -1 0 1020 0 -1 4305
box -2 -3 10 103
use NOR2X1  NOR2X1_410
timestamp 1693479267
transform -1 0 1044 0 -1 4305
box -2 -3 26 103
use NAND2X1  NAND2X1_916
timestamp 1693479267
transform -1 0 1068 0 -1 4305
box -2 -3 26 103
use NAND2X1  NAND2X1_806
timestamp 1693479267
transform -1 0 1092 0 -1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_876
timestamp 1693479267
transform 1 0 1092 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_872
timestamp 1693479267
transform 1 0 1124 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_869
timestamp 1693479267
transform 1 0 1156 0 -1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_401
timestamp 1693479267
transform 1 0 1188 0 -1 4305
box -2 -3 26 103
use OAI22X1  OAI22X1_45
timestamp 1693479267
transform -1 0 1252 0 -1 4305
box -2 -3 42 103
use AOI21X1  AOI21X1_223
timestamp 1693479267
transform -1 0 1284 0 -1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_125
timestamp 1693479267
transform -1 0 1380 0 -1 4305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_151
timestamp 1693479267
transform 1 0 1380 0 -1 4305
box -2 -3 98 103
use INVX1  INVX1_104
timestamp 1693479267
transform 1 0 1476 0 -1 4305
box -2 -3 18 103
use FILL  FILL_42_2_0
timestamp 1693479267
transform 1 0 1492 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_2_1
timestamp 1693479267
transform 1 0 1500 0 -1 4305
box -2 -3 10 103
use CLKBUF1  CLKBUF1_31
timestamp 1693479267
transform 1 0 1508 0 -1 4305
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_39
timestamp 1693479267
transform 1 0 1580 0 -1 4305
box -2 -3 98 103
use AOI22X1  AOI22X1_39
timestamp 1693479267
transform -1 0 1716 0 -1 4305
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_79
timestamp 1693479267
transform -1 0 1812 0 -1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_108
timestamp 1693479267
transform 1 0 1812 0 -1 4305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_77
timestamp 1693479267
transform -1 0 1940 0 -1 4305
box -2 -3 98 103
use OAI21X1  OAI21X1_100
timestamp 1693479267
transform -1 0 1972 0 -1 4305
box -2 -3 34 103
use INVX1  INVX1_100
timestamp 1693479267
transform -1 0 1988 0 -1 4305
box -2 -3 18 103
use NAND3X1  NAND3X1_188
timestamp 1693479267
transform -1 0 2020 0 -1 4305
box -2 -3 34 103
use INVX1  INVX1_130
timestamp 1693479267
transform 1 0 2020 0 -1 4305
box -2 -3 18 103
use FILL  FILL_42_3_0
timestamp 1693479267
transform 1 0 2036 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_3_1
timestamp 1693479267
transform 1 0 2044 0 -1 4305
box -2 -3 10 103
use OAI21X1  OAI21X1_160
timestamp 1693479267
transform 1 0 2052 0 -1 4305
box -2 -3 34 103
use INVX1  INVX1_614
timestamp 1693479267
transform -1 0 2100 0 -1 4305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_227
timestamp 1693479267
transform -1 0 2196 0 -1 4305
box -2 -3 98 103
use NAND3X1  NAND3X1_229
timestamp 1693479267
transform -1 0 2228 0 -1 4305
box -2 -3 34 103
use INVX1  INVX1_514
timestamp 1693479267
transform 1 0 2228 0 -1 4305
box -2 -3 18 103
use NAND3X1  NAND3X1_200
timestamp 1693479267
transform 1 0 2244 0 -1 4305
box -2 -3 34 103
use NAND3X1  NAND3X1_242
timestamp 1693479267
transform 1 0 2276 0 -1 4305
box -2 -3 34 103
use NAND3X1  NAND3X1_243
timestamp 1693479267
transform -1 0 2340 0 -1 4305
box -2 -3 34 103
use NAND3X1  NAND3X1_231
timestamp 1693479267
transform 1 0 2340 0 -1 4305
box -2 -3 34 103
use NAND3X1  NAND3X1_230
timestamp 1693479267
transform -1 0 2404 0 -1 4305
box -2 -3 34 103
use INVX1  INVX1_544
timestamp 1693479267
transform -1 0 2420 0 -1 4305
box -2 -3 18 103
use INVX1  INVX1_617
timestamp 1693479267
transform 1 0 2420 0 -1 4305
box -2 -3 18 103
use INVX1  INVX1_639
timestamp 1693479267
transform 1 0 2436 0 -1 4305
box -2 -3 18 103
use INVX1  INVX1_566
timestamp 1693479267
transform 1 0 2452 0 -1 4305
box -2 -3 18 103
use NAND3X1  NAND3X1_252
timestamp 1693479267
transform 1 0 2468 0 -1 4305
box -2 -3 34 103
use INVX1  INVX1_506
timestamp 1693479267
transform 1 0 2500 0 -1 4305
box -2 -3 18 103
use NAND3X1  NAND3X1_192
timestamp 1693479267
transform 1 0 2516 0 -1 4305
box -2 -3 34 103
use FILL  FILL_42_4_0
timestamp 1693479267
transform -1 0 2556 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_4_1
timestamp 1693479267
transform -1 0 2564 0 -1 4305
box -2 -3 10 103
use NAND3X1  NAND3X1_193
timestamp 1693479267
transform -1 0 2596 0 -1 4305
box -2 -3 34 103
use NAND3X1  NAND3X1_253
timestamp 1693479267
transform -1 0 2628 0 -1 4305
box -2 -3 34 103
use NAND3X1  NAND3X1_249
timestamp 1693479267
transform 1 0 2628 0 -1 4305
box -2 -3 34 103
use NAND3X1  NAND3X1_300
timestamp 1693479267
transform 1 0 2660 0 -1 4305
box -2 -3 34 103
use NAND3X1  NAND3X1_301
timestamp 1693479267
transform -1 0 2724 0 -1 4305
box -2 -3 34 103
use INVX1  INVX1_579
timestamp 1693479267
transform 1 0 2724 0 -1 4305
box -2 -3 18 103
use NAND3X1  NAND3X1_262
timestamp 1693479267
transform 1 0 2740 0 -1 4305
box -2 -3 34 103
use NAND3X1  NAND3X1_263
timestamp 1693479267
transform -1 0 2804 0 -1 4305
box -2 -3 34 103
use NAND3X1  NAND3X1_318
timestamp 1693479267
transform 1 0 2804 0 -1 4305
box -2 -3 34 103
use NAND3X1  NAND3X1_322
timestamp 1693479267
transform 1 0 2836 0 -1 4305
box -2 -3 34 103
use NAND3X1  NAND3X1_319
timestamp 1693479267
transform -1 0 2900 0 -1 4305
box -2 -3 34 103
use NAND3X1  NAND3X1_323
timestamp 1693479267
transform 1 0 2900 0 -1 4305
box -2 -3 34 103
use NAND3X1  NAND3X1_73
timestamp 1693479267
transform -1 0 2964 0 -1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_107
timestamp 1693479267
transform -1 0 2988 0 -1 4305
box -2 -3 26 103
use NOR2X1  NOR2X1_9
timestamp 1693479267
transform -1 0 3012 0 -1 4305
box -2 -3 26 103
use INVX1  INVX1_223
timestamp 1693479267
transform 1 0 3012 0 -1 4305
box -2 -3 18 103
use AOI22X1  AOI22X1_40
timestamp 1693479267
transform -1 0 3068 0 -1 4305
box -2 -3 42 103
use FILL  FILL_42_5_0
timestamp 1693479267
transform -1 0 3076 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_5_1
timestamp 1693479267
transform -1 0 3084 0 -1 4305
box -2 -3 10 103
use INVX1  INVX1_224
timestamp 1693479267
transform -1 0 3100 0 -1 4305
box -2 -3 18 103
use INVX1  INVX1_191
timestamp 1693479267
transform 1 0 3100 0 -1 4305
box -2 -3 18 103
use NOR2X1  NOR2X1_12
timestamp 1693479267
transform -1 0 3140 0 -1 4305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_5
timestamp 1693479267
transform -1 0 3236 0 -1 4305
box -2 -3 98 103
use NAND2X1  NAND2X1_1000
timestamp 1693479267
transform -1 0 3260 0 -1 4305
box -2 -3 26 103
use INVX1  INVX1_717
timestamp 1693479267
transform 1 0 3260 0 -1 4305
box -2 -3 18 103
use NAND3X1  NAND3X1_354
timestamp 1693479267
transform 1 0 3276 0 -1 4305
box -2 -3 34 103
use NAND3X1  NAND3X1_352
timestamp 1693479267
transform 1 0 3308 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_944
timestamp 1693479267
transform -1 0 3372 0 -1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_475
timestamp 1693479267
transform -1 0 3396 0 -1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_943
timestamp 1693479267
transform -1 0 3428 0 -1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_1010
timestamp 1693479267
transform 1 0 3428 0 -1 4305
box -2 -3 26 103
use AOI21X1  AOI21X1_259
timestamp 1693479267
transform 1 0 3452 0 -1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_998
timestamp 1693479267
transform -1 0 3508 0 -1 4305
box -2 -3 26 103
use NAND2X1  NAND2X1_1011
timestamp 1693479267
transform -1 0 3532 0 -1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_1056
timestamp 1693479267
transform 1 0 3532 0 -1 4305
box -2 -3 34 103
use FILL  FILL_42_6_0
timestamp 1693479267
transform -1 0 3572 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_6_1
timestamp 1693479267
transform -1 0 3580 0 -1 4305
box -2 -3 10 103
use AOI21X1  AOI21X1_270
timestamp 1693479267
transform -1 0 3612 0 -1 4305
box -2 -3 34 103
use AOI21X1  AOI21X1_269
timestamp 1693479267
transform -1 0 3644 0 -1 4305
box -2 -3 34 103
use AOI21X1  AOI21X1_268
timestamp 1693479267
transform -1 0 3676 0 -1 4305
box -2 -3 34 103
use AOI21X1  AOI21X1_271
timestamp 1693479267
transform 1 0 3676 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_945
timestamp 1693479267
transform -1 0 3740 0 -1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_1018
timestamp 1693479267
transform -1 0 3764 0 -1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_1010
timestamp 1693479267
transform -1 0 3796 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_982
timestamp 1693479267
transform -1 0 3828 0 -1 4305
box -2 -3 34 103
use AOI21X1  AOI21X1_257
timestamp 1693479267
transform -1 0 3860 0 -1 4305
box -2 -3 34 103
use AOI22X1  AOI22X1_144
timestamp 1693479267
transform -1 0 3900 0 -1 4305
box -2 -3 42 103
use INVX2  INVX2_91
timestamp 1693479267
transform 1 0 3900 0 -1 4305
box -2 -3 18 103
use OAI21X1  OAI21X1_1003
timestamp 1693479267
transform 1 0 3916 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1004
timestamp 1693479267
transform -1 0 3980 0 -1 4305
box -2 -3 34 103
use AOI21X1  AOI21X1_264
timestamp 1693479267
transform -1 0 4012 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1006
timestamp 1693479267
transform -1 0 4044 0 -1 4305
box -2 -3 34 103
use INVX1  INVX1_750
timestamp 1693479267
transform -1 0 4060 0 -1 4305
box -2 -3 18 103
use INVX1  INVX1_743
timestamp 1693479267
transform 1 0 4060 0 -1 4305
box -2 -3 18 103
use FILL  FILL_42_7_0
timestamp 1693479267
transform 1 0 4076 0 -1 4305
box -2 -3 10 103
use FILL  FILL_42_7_1
timestamp 1693479267
transform 1 0 4084 0 -1 4305
box -2 -3 10 103
use OAI22X1  OAI22X1_56
timestamp 1693479267
transform 1 0 4092 0 -1 4305
box -2 -3 42 103
use AOI22X1  AOI22X1_140
timestamp 1693479267
transform 1 0 4132 0 -1 4305
box -2 -3 42 103
use OAI21X1  OAI21X1_993
timestamp 1693479267
transform -1 0 4204 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_994
timestamp 1693479267
transform -1 0 4236 0 -1 4305
box -2 -3 34 103
use AOI21X1  AOI21X1_261
timestamp 1693479267
transform -1 0 4268 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_992
timestamp 1693479267
transform 1 0 4268 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_999
timestamp 1693479267
transform -1 0 4332 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1021
timestamp 1693479267
transform -1 0 4364 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1000
timestamp 1693479267
transform -1 0 4396 0 -1 4305
box -2 -3 34 103
use AOI21X1  AOI21X1_263
timestamp 1693479267
transform 1 0 4396 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1002
timestamp 1693479267
transform 1 0 4428 0 -1 4305
box -2 -3 34 103
use AOI22X1  AOI22X1_142
timestamp 1693479267
transform 1 0 4460 0 -1 4305
box -2 -3 42 103
use NAND2X1  NAND2X1_1016
timestamp 1693479267
transform 1 0 4500 0 -1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_1001
timestamp 1693479267
transform -1 0 4556 0 -1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1018
timestamp 1693479267
transform 1 0 4556 0 -1 4305
box -2 -3 34 103
use FILL  FILL_43_1
timestamp 1693479267
transform -1 0 4596 0 -1 4305
box -2 -3 10 103
use FILL  FILL_43_2
timestamp 1693479267
transform -1 0 4604 0 -1 4305
box -2 -3 10 103
use INVX1  INVX1_175
timestamp 1693479267
transform 1 0 4 0 1 4305
box -2 -3 18 103
use NOR3X1  NOR3X1_34
timestamp 1693479267
transform -1 0 84 0 1 4305
box -2 -3 66 103
use NOR3X1  NOR3X1_35
timestamp 1693479267
transform -1 0 148 0 1 4305
box -2 -3 66 103
use INVX1  INVX1_176
timestamp 1693479267
transform -1 0 164 0 1 4305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_427
timestamp 1693479267
transform 1 0 164 0 1 4305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_428
timestamp 1693479267
transform 1 0 260 0 1 4305
box -2 -3 98 103
use XOR2X1  XOR2X1_13
timestamp 1693479267
transform 1 0 356 0 1 4305
box -2 -3 58 103
use XOR2X1  XOR2X1_17
timestamp 1693479267
transform 1 0 412 0 1 4305
box -2 -3 58 103
use FILL  FILL_43_0_0
timestamp 1693479267
transform -1 0 476 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_0_1
timestamp 1693479267
transform -1 0 484 0 1 4305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_42
timestamp 1693479267
transform -1 0 580 0 1 4305
box -2 -3 98 103
use OR2X2  OR2X2_50
timestamp 1693479267
transform 1 0 580 0 1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_815
timestamp 1693479267
transform 1 0 612 0 1 4305
box -2 -3 26 103
use NAND2X1  NAND2X1_705
timestamp 1693479267
transform 1 0 636 0 1 4305
box -2 -3 26 103
use AOI22X1  AOI22X1_110
timestamp 1693479267
transform -1 0 700 0 1 4305
box -2 -3 42 103
use OR2X2  OR2X2_49
timestamp 1693479267
transform 1 0 700 0 1 4305
box -2 -3 34 103
use AOI21X1  AOI21X1_225
timestamp 1693479267
transform 1 0 732 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_870
timestamp 1693479267
transform 1 0 764 0 1 4305
box -2 -3 34 103
use INVX1  INVX1_567
timestamp 1693479267
transform -1 0 812 0 1 4305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_40
timestamp 1693479267
transform 1 0 812 0 1 4305
box -2 -3 98 103
use INVX1  INVX1_640
timestamp 1693479267
transform 1 0 908 0 1 4305
box -2 -3 18 103
use OAI21X1  OAI21X1_874
timestamp 1693479267
transform -1 0 956 0 1 4305
box -2 -3 34 103
use AOI21X1  AOI21X1_229
timestamp 1693479267
transform -1 0 988 0 1 4305
box -2 -3 34 103
use FILL  FILL_43_1_0
timestamp 1693479267
transform -1 0 996 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_1_1
timestamp 1693479267
transform -1 0 1004 0 1 4305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_41
timestamp 1693479267
transform -1 0 1100 0 1 4305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_43
timestamp 1693479267
transform -1 0 1196 0 1 4305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_45
timestamp 1693479267
transform 1 0 1196 0 1 4305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_13
timestamp 1693479267
transform 1 0 1292 0 1 4305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_51
timestamp 1693479267
transform 1 0 1388 0 1 4305
box -2 -3 98 103
use AOI22X1  AOI22X1_13
timestamp 1693479267
transform 1 0 1484 0 1 4305
box -2 -3 42 103
use FILL  FILL_43_2_0
timestamp 1693479267
transform -1 0 1532 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_2_1
timestamp 1693479267
transform -1 0 1540 0 1 4305
box -2 -3 10 103
use OAI21X1  OAI21X1_198
timestamp 1693479267
transform -1 0 1572 0 1 4305
box -2 -3 34 103
use INVX1  INVX1_196
timestamp 1693479267
transform -1 0 1588 0 1 4305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_9
timestamp 1693479267
transform 1 0 1588 0 1 4305
box -2 -3 98 103
use AOI22X1  AOI22X1_9
timestamp 1693479267
transform -1 0 1724 0 1 4305
box -2 -3 42 103
use INVX1  INVX1_192
timestamp 1693479267
transform 1 0 1724 0 1 4305
box -2 -3 18 103
use OAI21X1  OAI21X1_194
timestamp 1693479267
transform -1 0 1772 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_224
timestamp 1693479267
transform -1 0 1804 0 1 4305
box -2 -3 34 103
use INVX1  INVX1_222
timestamp 1693479267
transform -1 0 1820 0 1 4305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_109
timestamp 1693479267
transform -1 0 1916 0 1 4305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_47
timestamp 1693479267
transform -1 0 2012 0 1 4305
box -2 -3 98 103
use FILL  FILL_43_3_0
timestamp 1693479267
transform -1 0 2020 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_3_1
timestamp 1693479267
transform -1 0 2028 0 1 4305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_83
timestamp 1693479267
transform -1 0 2124 0 1 4305
box -2 -3 98 103
use INVX1  INVX1_541
timestamp 1693479267
transform 1 0 2124 0 1 4305
box -2 -3 18 103
use BUFX4  BUFX4_203
timestamp 1693479267
transform -1 0 2172 0 1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_767
timestamp 1693479267
transform 1 0 2172 0 1 4305
box -2 -3 26 103
use INVX1  INVX1_628
timestamp 1693479267
transform 1 0 2196 0 1 4305
box -2 -3 18 103
use INVX1  INVX1_555
timestamp 1693479267
transform 1 0 2212 0 1 4305
box -2 -3 18 103
use NAND2X1  NAND2X1_788
timestamp 1693479267
transform 1 0 2228 0 1 4305
box -2 -3 26 103
use BUFX2  BUFX2_76
timestamp 1693479267
transform 1 0 2252 0 1 4305
box -2 -3 26 103
use BUFX4  BUFX4_204
timestamp 1693479267
transform -1 0 2308 0 1 4305
box -2 -3 34 103
use BUFX4  BUFX4_210
timestamp 1693479267
transform 1 0 2308 0 1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_770
timestamp 1693479267
transform -1 0 2364 0 1 4305
box -2 -3 26 103
use INVX1  INVX1_543
timestamp 1693479267
transform -1 0 2380 0 1 4305
box -2 -3 18 103
use INVX1  INVX1_616
timestamp 1693479267
transform 1 0 2380 0 1 4305
box -2 -3 18 103
use NAND2X1  NAND2X1_880
timestamp 1693479267
transform 1 0 2396 0 1 4305
box -2 -3 26 103
use BUFX4  BUFX4_103
timestamp 1693479267
transform 1 0 2420 0 1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_823
timestamp 1693479267
transform -1 0 2476 0 1 4305
box -2 -3 26 103
use INVX1  INVX1_578
timestamp 1693479267
transform -1 0 2492 0 1 4305
box -2 -3 18 103
use INVX1  INVX1_505
timestamp 1693479267
transform 1 0 2492 0 1 4305
box -2 -3 18 103
use NAND2X1  NAND2X1_713
timestamp 1693479267
transform 1 0 2508 0 1 4305
box -2 -3 26 103
use NAND2X1  NAND2X1_803
timestamp 1693479267
transform -1 0 2556 0 1 4305
box -2 -3 26 103
use FILL  FILL_43_4_0
timestamp 1693479267
transform -1 0 2564 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_4_1
timestamp 1693479267
transform -1 0 2572 0 1 4305
box -2 -3 10 103
use INVX1  INVX1_565
timestamp 1693479267
transform -1 0 2588 0 1 4305
box -2 -3 18 103
use INVX1  INVX1_638
timestamp 1693479267
transform 1 0 2588 0 1 4305
box -2 -3 18 103
use NAND2X1  NAND2X1_797
timestamp 1693479267
transform -1 0 2628 0 1 4305
box -2 -3 26 103
use INVX1  INVX1_561
timestamp 1693479267
transform -1 0 2644 0 1 4305
box -2 -3 18 103
use INVX1  INVX1_634
timestamp 1693479267
transform 1 0 2644 0 1 4305
box -2 -3 18 103
use NAND2X1  NAND2X1_913
timestamp 1693479267
transform 1 0 2660 0 1 4305
box -2 -3 26 103
use NAND2X1  NAND2X1_907
timestamp 1693479267
transform 1 0 2684 0 1 4305
box -2 -3 26 103
use OR2X2  OR2X2_4
timestamp 1693479267
transform 1 0 2708 0 1 4305
box -2 -3 34 103
use BUFX2  BUFX2_2
timestamp 1693479267
transform -1 0 2764 0 1 4305
box -2 -3 26 103
use BUFX2  BUFX2_1
timestamp 1693479267
transform -1 0 2788 0 1 4305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_7
timestamp 1693479267
transform 1 0 2788 0 1 4305
box -2 -3 98 103
use INVX1  INVX1_190
timestamp 1693479267
transform 1 0 2884 0 1 4305
box -2 -3 18 103
use NAND2X1  NAND2X1_105
timestamp 1693479267
transform -1 0 2924 0 1 4305
box -2 -3 26 103
use NOR2X1  NOR2X1_13
timestamp 1693479267
transform 1 0 2924 0 1 4305
box -2 -3 26 103
use NAND2X1  NAND2X1_106
timestamp 1693479267
transform 1 0 2948 0 1 4305
box -2 -3 26 103
use NOR2X1  NOR2X1_11
timestamp 1693479267
transform 1 0 2972 0 1 4305
box -2 -3 26 103
use INVX1  INVX1_189
timestamp 1693479267
transform 1 0 2996 0 1 4305
box -2 -3 18 103
use FILL  FILL_43_5_0
timestamp 1693479267
transform -1 0 3020 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_5_1
timestamp 1693479267
transform -1 0 3028 0 1 4305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_6
timestamp 1693479267
transform -1 0 3124 0 1 4305
box -2 -3 98 103
use BUFX2  BUFX2_75
timestamp 1693479267
transform -1 0 3148 0 1 4305
box -2 -3 26 103
use BUFX2  BUFX2_74
timestamp 1693479267
transform -1 0 3172 0 1 4305
box -2 -3 26 103
use BUFX2  BUFX2_72
timestamp 1693479267
transform 1 0 3172 0 1 4305
box -2 -3 26 103
use BUFX2  BUFX2_73
timestamp 1693479267
transform 1 0 3196 0 1 4305
box -2 -3 26 103
use INVX4  INVX4_12
timestamp 1693479267
transform -1 0 3244 0 1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_948
timestamp 1693479267
transform -1 0 3276 0 1 4305
box -2 -3 34 103
use BUFX2  BUFX2_33
timestamp 1693479267
transform 1 0 3276 0 1 4305
box -2 -3 26 103
use INVX1  INVX1_756
timestamp 1693479267
transform 1 0 3300 0 1 4305
box -2 -3 18 103
use BUFX2  BUFX2_38
timestamp 1693479267
transform -1 0 3340 0 1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_1058
timestamp 1693479267
transform -1 0 3372 0 1 4305
box -2 -3 34 103
use BUFX2  BUFX2_34
timestamp 1693479267
transform -1 0 3396 0 1 4305
box -2 -3 26 103
use BUFX2  BUFX2_36
timestamp 1693479267
transform -1 0 3420 0 1 4305
box -2 -3 26 103
use NAND3X1  NAND3X1_355
timestamp 1693479267
transform 1 0 3420 0 1 4305
box -2 -3 34 103
use BUFX2  BUFX2_37
timestamp 1693479267
transform -1 0 3476 0 1 4305
box -2 -3 26 103
use NAND3X1  NAND3X1_349
timestamp 1693479267
transform 1 0 3476 0 1 4305
box -2 -3 34 103
use BUFX2  BUFX2_35
timestamp 1693479267
transform 1 0 3508 0 1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_980
timestamp 1693479267
transform 1 0 3532 0 1 4305
box -2 -3 34 103
use FILL  FILL_43_6_0
timestamp 1693479267
transform -1 0 3572 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_6_1
timestamp 1693479267
transform -1 0 3580 0 1 4305
box -2 -3 10 103
use OAI21X1  OAI21X1_981
timestamp 1693479267
transform -1 0 3612 0 1 4305
box -2 -3 34 103
use INVX1  INVX1_735
timestamp 1693479267
transform -1 0 3628 0 1 4305
box -2 -3 18 103
use OAI22X1  OAI22X1_53
timestamp 1693479267
transform -1 0 3668 0 1 4305
box -2 -3 42 103
use AOI22X1  AOI22X1_137
timestamp 1693479267
transform -1 0 3708 0 1 4305
box -2 -3 42 103
use NAND2X1  NAND2X1_1017
timestamp 1693479267
transform -1 0 3732 0 1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_1005
timestamp 1693479267
transform -1 0 3764 0 1 4305
box -2 -3 34 103
use AOI22X1  AOI22X1_143
timestamp 1693479267
transform -1 0 3804 0 1 4305
box -2 -3 42 103
use INVX1  INVX1_752
timestamp 1693479267
transform 1 0 3804 0 1 4305
box -2 -3 18 103
use OAI22X1  OAI22X1_59
timestamp 1693479267
transform -1 0 3860 0 1 4305
box -2 -3 42 103
use INVX1  INVX1_751
timestamp 1693479267
transform -1 0 3876 0 1 4305
box -2 -3 18 103
use INVX2  INVX2_92
timestamp 1693479267
transform 1 0 3876 0 1 4305
box -2 -3 18 103
use AOI22X1  AOI22X1_149
timestamp 1693479267
transform 1 0 3892 0 1 4305
box -2 -3 42 103
use OAI21X1  OAI21X1_1029
timestamp 1693479267
transform 1 0 3932 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1028
timestamp 1693479267
transform 1 0 3964 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1019
timestamp 1693479267
transform 1 0 3996 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1020
timestamp 1693479267
transform -1 0 4060 0 1 4305
box -2 -3 34 103
use NAND2X1  NAND2X1_1014
timestamp 1693479267
transform -1 0 4084 0 1 4305
box -2 -3 26 103
use FILL  FILL_43_7_0
timestamp 1693479267
transform -1 0 4092 0 1 4305
box -2 -3 10 103
use FILL  FILL_43_7_1
timestamp 1693479267
transform -1 0 4100 0 1 4305
box -2 -3 10 103
use INVX1  INVX1_742
timestamp 1693479267
transform -1 0 4116 0 1 4305
box -2 -3 18 103
use AOI22X1  AOI22X1_146
timestamp 1693479267
transform -1 0 4156 0 1 4305
box -2 -3 42 103
use OAI21X1  OAI21X1_1030
timestamp 1693479267
transform -1 0 4188 0 1 4305
box -2 -3 34 103
use OAI21X1  OAI21X1_1025
timestamp 1693479267
transform 1 0 4188 0 1 4305
box -2 -3 34 103
use INVX1  INVX1_749
timestamp 1693479267
transform -1 0 4236 0 1 4305
box -2 -3 18 103
use OAI22X1  OAI22X1_58
timestamp 1693479267
transform -1 0 4276 0 1 4305
box -2 -3 42 103
use OAI21X1  OAI21X1_1026
timestamp 1693479267
transform -1 0 4308 0 1 4305
box -2 -3 34 103
use INVX1  INVX1_748
timestamp 1693479267
transform -1 0 4324 0 1 4305
box -2 -3 18 103
use AOI22X1  AOI22X1_148
timestamp 1693479267
transform -1 0 4364 0 1 4305
box -2 -3 42 103
use OAI21X1  OAI21X1_1027
timestamp 1693479267
transform -1 0 4396 0 1 4305
box -2 -3 34 103
use AOI22X1  AOI22X1_156
timestamp 1693479267
transform -1 0 4436 0 1 4305
box -2 -3 42 103
use OAI21X1  OAI21X1_740
timestamp 1693479267
transform -1 0 4468 0 1 4305
box -2 -3 34 103
use NOR2X1  NOR2X1_365
timestamp 1693479267
transform -1 0 4492 0 1 4305
box -2 -3 26 103
use NOR2X1  NOR2X1_357
timestamp 1693479267
transform -1 0 4516 0 1 4305
box -2 -3 26 103
use NOR2X1  NOR2X1_249
timestamp 1693479267
transform -1 0 4540 0 1 4305
box -2 -3 26 103
use BUFX2  BUFX2_81
timestamp 1693479267
transform 1 0 4540 0 1 4305
box -2 -3 26 103
use OAI21X1  OAI21X1_1040
timestamp 1693479267
transform -1 0 4596 0 1 4305
box -2 -3 34 103
use FILL  FILL_44_1
timestamp 1693479267
transform 1 0 4596 0 1 4305
box -2 -3 10 103
<< labels >>
flabel metal6 s 496 -30 512 -22 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal6 s 1000 -30 1016 -22 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal2 s 1998 4428 2002 4432 3 FreeSans 24 90 0 0 CLK
port 2 nsew
flabel metal3 s -26 2088 -22 2092 7 FreeSans 24 0 0 0 reset
port 3 nsew
flabel metal3 s -26 3148 -22 3152 7 FreeSans 24 0 0 0 instruction_memory_interface_data[0]
port 4 nsew
flabel metal3 s -26 3048 -22 3052 7 FreeSans 24 0 0 0 instruction_memory_interface_data[1]
port 5 nsew
flabel metal3 s -26 3168 -22 3172 7 FreeSans 24 0 0 0 instruction_memory_interface_data[2]
port 6 nsew
flabel metal3 s -26 2868 -22 2872 7 FreeSans 24 0 0 0 instruction_memory_interface_data[3]
port 7 nsew
flabel metal3 s -26 3128 -22 3132 7 FreeSans 24 0 0 0 instruction_memory_interface_data[4]
port 8 nsew
flabel metal3 s -26 3448 -22 3452 7 FreeSans 24 0 0 0 instruction_memory_interface_data[5]
port 9 nsew
flabel metal3 s -26 3348 -22 3352 7 FreeSans 24 0 0 0 instruction_memory_interface_data[6]
port 10 nsew
flabel metal3 s -26 2948 -22 2952 7 FreeSans 24 0 0 0 instruction_memory_interface_data[7]
port 11 nsew
flabel metal3 s -26 3948 -22 3952 7 FreeSans 24 0 0 0 instruction_memory_interface_data[8]
port 12 nsew
flabel metal3 s -26 3548 -22 3552 7 FreeSans 24 0 0 0 instruction_memory_interface_data[9]
port 13 nsew
flabel metal3 s -26 3648 -22 3652 7 FreeSans 24 0 0 0 instruction_memory_interface_data[10]
port 14 nsew
flabel metal3 s -26 3528 -22 3532 7 FreeSans 24 0 0 0 instruction_memory_interface_data[11]
port 15 nsew
flabel metal3 s -26 2148 -22 2152 7 FreeSans 24 0 0 0 instruction_memory_interface_data[12]
port 16 nsew
flabel metal3 s -26 2358 -22 2362 7 FreeSans 24 0 0 0 instruction_memory_interface_data[13]
port 17 nsew
flabel metal3 s -26 2558 -22 2562 7 FreeSans 24 0 0 0 instruction_memory_interface_data[14]
port 18 nsew
flabel metal3 s -26 3748 -22 3752 7 FreeSans 24 0 0 0 instruction_memory_interface_data[15]
port 19 nsew
flabel metal3 s -26 4148 -22 4152 7 FreeSans 24 0 0 0 instruction_memory_interface_data[16]
port 20 nsew
flabel metal3 s -26 3668 -22 3672 7 FreeSans 24 0 0 0 instruction_memory_interface_data[17]
port 21 nsew
flabel metal3 s -26 3968 -22 3972 7 FreeSans 24 0 0 0 instruction_memory_interface_data[18]
port 22 nsew
flabel metal3 s -26 4348 -22 4352 7 FreeSans 24 90 0 0 instruction_memory_interface_data[19]
port 23 nsew
flabel metal2 s 150 4428 154 4432 3 FreeSans 24 90 0 0 instruction_memory_interface_data[20]
port 24 nsew
flabel metal3 s -26 2848 -22 2852 7 FreeSans 24 0 0 0 instruction_memory_interface_data[21]
port 25 nsew
flabel metal3 s -26 4248 -22 4252 7 FreeSans 24 0 0 0 instruction_memory_interface_data[22]
port 26 nsew
flabel metal3 s -26 3848 -22 3852 7 FreeSans 24 0 0 0 instruction_memory_interface_data[23]
port 27 nsew
flabel metal3 s -26 2668 -22 2672 7 FreeSans 24 0 0 0 instruction_memory_interface_data[24]
port 28 nsew
flabel metal3 s -26 2338 -22 2342 7 FreeSans 24 0 0 0 instruction_memory_interface_data[25]
port 29 nsew
flabel metal3 s -26 2728 -22 2732 7 FreeSans 24 0 0 0 instruction_memory_interface_data[26]
port 30 nsew
flabel metal3 s -26 2648 -22 2652 7 FreeSans 24 0 0 0 instruction_memory_interface_data[27]
port 31 nsew
flabel metal3 s -26 2748 -22 2752 7 FreeSans 24 0 0 0 instruction_memory_interface_data[28]
port 32 nsew
flabel metal3 s -26 2448 -22 2452 7 FreeSans 24 0 0 0 instruction_memory_interface_data[29]
port 33 nsew
flabel metal3 s -26 2538 -22 2542 7 FreeSans 24 0 0 0 instruction_memory_interface_data[30]
port 34 nsew
flabel metal3 s -26 2268 -22 2272 7 FreeSans 24 0 0 0 instruction_memory_interface_data[31]
port 35 nsew
flabel metal2 s 3686 4428 3690 4432 3 FreeSans 24 90 0 0 data_memory_interface_data[0]
port 36 nsew
flabel metal2 s 4126 4428 4130 4432 3 FreeSans 24 90 0 0 data_memory_interface_data[1]
port 37 nsew
flabel metal2 s 3750 4428 3754 4432 3 FreeSans 24 90 0 0 data_memory_interface_data[2]
port 38 nsew
flabel metal2 s 4102 4428 4106 4432 3 FreeSans 24 90 0 0 data_memory_interface_data[3]
port 39 nsew
flabel metal3 s 4630 3938 4634 3942 3 FreeSans 24 0 0 0 data_memory_interface_data[4]
port 40 nsew
flabel metal2 s 4230 4428 4234 4432 3 FreeSans 24 90 0 0 data_memory_interface_data[5]
port 41 nsew
flabel metal2 s 3790 4428 3794 4432 3 FreeSans 24 90 0 0 data_memory_interface_data[6]
port 42 nsew
flabel metal2 s 3918 4428 3922 4432 3 FreeSans 24 90 0 0 data_memory_interface_data[7]
port 43 nsew
flabel metal2 s 3878 4428 3882 4432 3 FreeSans 24 90 0 0 data_memory_interface_data[8]
port 44 nsew
flabel metal3 s 4630 4148 4634 4152 3 FreeSans 24 0 0 0 data_memory_interface_data[9]
port 45 nsew
flabel metal2 s 4142 4428 4146 4432 3 FreeSans 24 90 0 0 data_memory_interface_data[10]
port 46 nsew
flabel metal3 s 4630 4048 4634 4052 3 FreeSans 24 0 0 0 data_memory_interface_data[11]
port 47 nsew
flabel metal2 s 4342 4428 4346 4432 3 FreeSans 24 90 0 0 data_memory_interface_data[12]
port 48 nsew
flabel metal2 s 3902 4428 3906 4432 3 FreeSans 24 90 0 0 data_memory_interface_data[13]
port 49 nsew
flabel metal2 s 3982 4428 3986 4432 3 FreeSans 24 90 0 0 data_memory_interface_data[14]
port 50 nsew
flabel metal2 s 3942 4428 3946 4432 3 FreeSans 24 90 0 0 data_memory_interface_data[15]
port 51 nsew
flabel metal2 s 3558 4428 3562 4432 3 FreeSans 24 90 0 0 data_memory_interface_data[16]
port 52 nsew
flabel metal3 s 4630 3848 4634 3852 3 FreeSans 24 0 0 0 data_memory_interface_data[17]
port 53 nsew
flabel metal3 s 4630 3748 4634 3752 3 FreeSans 24 0 0 0 data_memory_interface_data[18]
port 54 nsew
flabel metal3 s 4630 3768 4634 3772 3 FreeSans 24 0 0 0 data_memory_interface_data[19]
port 55 nsew
flabel metal3 s 4630 4168 4634 4172 3 FreeSans 24 0 0 0 data_memory_interface_data[20]
port 56 nsew
flabel metal3 s 4630 3958 4634 3962 3 FreeSans 24 0 0 0 data_memory_interface_data[21]
port 57 nsew
flabel metal2 s 4062 4428 4066 4432 3 FreeSans 24 90 0 0 data_memory_interface_data[22]
port 58 nsew
flabel metal2 s 3766 4428 3770 4432 3 FreeSans 24 90 0 0 data_memory_interface_data[23]
port 59 nsew
flabel metal2 s 4022 4428 4026 4432 3 FreeSans 24 90 0 0 data_memory_interface_data[24]
port 60 nsew
flabel metal2 s 4430 4428 4434 4432 3 FreeSans 24 90 0 0 data_memory_interface_data[25]
port 61 nsew
flabel metal2 s 4046 4428 4050 4432 3 FreeSans 24 90 0 0 data_memory_interface_data[26]
port 62 nsew
flabel metal2 s 4382 4428 4386 4432 3 FreeSans 24 90 0 0 data_memory_interface_data[27]
port 63 nsew
flabel metal2 s 4214 4428 4218 4432 3 FreeSans 24 90 0 0 data_memory_interface_data[28]
port 64 nsew
flabel metal2 s 4006 4428 4010 4432 3 FreeSans 24 90 0 0 data_memory_interface_data[29]
port 65 nsew
flabel metal2 s 3966 4428 3970 4432 3 FreeSans 24 90 0 0 data_memory_interface_data[30]
port 66 nsew
flabel metal2 s 3830 4428 3834 4432 3 FreeSans 24 90 0 0 data_memory_interface_data[31]
port 67 nsew
flabel metal2 s 110 -22 114 -18 7 FreeSans 24 270 0 0 instruction_memory_interface_enable
port 68 nsew
flabel metal2 s 2262 4428 2266 4432 3 FreeSans 24 90 0 0 instruction_memory_interface_state
port 69 nsew
flabel metal3 s -26 2208 -22 2212 7 FreeSans 24 0 0 0 instruction_memory_interface_address[0]
port 70 nsew
flabel metal3 s -26 2048 -22 2052 7 FreeSans 24 0 0 0 instruction_memory_interface_address[1]
port 71 nsew
flabel metal2 s 750 -22 754 -18 7 FreeSans 24 270 0 0 instruction_memory_interface_address[2]
port 72 nsew
flabel metal2 s 766 -22 770 -18 7 FreeSans 24 270 0 0 instruction_memory_interface_address[3]
port 73 nsew
flabel metal2 s 966 -22 970 -18 7 FreeSans 24 270 0 0 instruction_memory_interface_address[4]
port 74 nsew
flabel metal2 s 990 -22 994 -18 7 FreeSans 24 270 0 0 instruction_memory_interface_address[5]
port 75 nsew
flabel metal2 s 470 -22 474 -18 7 FreeSans 24 270 0 0 instruction_memory_interface_address[6]
port 76 nsew
flabel metal2 s 534 -22 538 -18 7 FreeSans 24 270 0 0 instruction_memory_interface_address[7]
port 77 nsew
flabel metal3 s -26 248 -22 252 7 FreeSans 24 0 0 0 instruction_memory_interface_address[8]
port 78 nsew
flabel metal2 s 1350 -22 1354 -18 7 FreeSans 24 270 0 0 instruction_memory_interface_address[9]
port 79 nsew
flabel metal3 s -26 48 -22 52 7 FreeSans 24 270 0 0 instruction_memory_interface_address[10]
port 80 nsew
flabel metal3 s -26 448 -22 452 7 FreeSans 24 0 0 0 instruction_memory_interface_address[11]
port 81 nsew
flabel metal2 s 350 -22 354 -18 7 FreeSans 24 270 0 0 instruction_memory_interface_address[12]
port 82 nsew
flabel metal2 s 630 -22 634 -18 7 FreeSans 24 270 0 0 instruction_memory_interface_address[13]
port 83 nsew
flabel metal2 s 942 -22 946 -18 7 FreeSans 24 270 0 0 instruction_memory_interface_address[14]
port 84 nsew
flabel metal2 s 822 -22 826 -18 7 FreeSans 24 270 0 0 instruction_memory_interface_address[15]
port 85 nsew
flabel metal3 s -26 648 -22 652 7 FreeSans 24 0 0 0 instruction_memory_interface_address[16]
port 86 nsew
flabel metal3 s -26 548 -22 552 7 FreeSans 24 0 0 0 instruction_memory_interface_address[17]
port 87 nsew
flabel metal3 s -26 868 -22 872 7 FreeSans 24 0 0 0 instruction_memory_interface_address[18]
port 88 nsew
flabel metal3 s -26 1148 -22 1152 7 FreeSans 24 0 0 0 instruction_memory_interface_address[19]
port 89 nsew
flabel metal3 s -26 1068 -22 1072 7 FreeSans 24 0 0 0 instruction_memory_interface_address[20]
port 90 nsew
flabel metal3 s -26 1168 -22 1172 7 FreeSans 24 0 0 0 instruction_memory_interface_address[21]
port 91 nsew
flabel metal3 s -26 1468 -22 1472 7 FreeSans 24 0 0 0 instruction_memory_interface_address[22]
port 92 nsew
flabel metal3 s -26 1568 -22 1572 7 FreeSans 24 0 0 0 instruction_memory_interface_address[23]
port 93 nsew
flabel metal3 s -26 1768 -22 1772 7 FreeSans 24 0 0 0 instruction_memory_interface_address[24]
port 94 nsew
flabel metal3 s -26 1968 -22 1972 7 FreeSans 24 0 0 0 instruction_memory_interface_address[25]
port 95 nsew
flabel metal3 s -26 1748 -22 1752 7 FreeSans 24 0 0 0 instruction_memory_interface_address[26]
port 96 nsew
flabel metal3 s -26 1788 -22 1792 7 FreeSans 24 0 0 0 instruction_memory_interface_address[27]
port 97 nsew
flabel metal3 s -26 2228 -22 2232 7 FreeSans 24 0 0 0 instruction_memory_interface_address[28]
port 98 nsew
flabel metal3 s -26 1868 -22 1872 7 FreeSans 24 0 0 0 instruction_memory_interface_address[29]
port 99 nsew
flabel metal3 s -26 1668 -22 1672 7 FreeSans 24 0 0 0 instruction_memory_interface_address[30]
port 100 nsew
flabel metal3 s -26 1548 -22 1552 7 FreeSans 24 0 0 0 instruction_memory_interface_address[31]
port 101 nsew
flabel metal2 s 3182 4428 3186 4432 3 FreeSans 24 90 0 0 instruction_memory_interface_frame_mask[0]
port 102 nsew
flabel metal2 s 3206 4428 3210 4432 3 FreeSans 24 90 0 0 instruction_memory_interface_frame_mask[1]
port 103 nsew
flabel metal2 s 3158 4428 3162 4432 3 FreeSans 24 90 0 0 instruction_memory_interface_frame_mask[2]
port 104 nsew
flabel metal2 s 3134 4428 3138 4432 3 FreeSans 24 90 0 0 instruction_memory_interface_frame_mask[3]
port 105 nsew
flabel metal2 s 3286 4428 3290 4432 3 FreeSans 24 90 0 0 data_memory_interface_enable
port 106 nsew
flabel metal2 s 3326 4428 3330 4432 3 FreeSans 24 90 0 0 data_memory_interface_state
port 107 nsew
flabel metal2 s 2774 4428 2778 4432 3 FreeSans 24 90 0 0 data_memory_interface_address[0]
port 108 nsew
flabel metal2 s 2750 4428 2754 4432 3 FreeSans 24 90 0 0 data_memory_interface_address[1]
port 109 nsew
flabel metal3 s -26 1848 -22 1852 7 FreeSans 24 0 0 0 data_memory_interface_address[2]
port 110 nsew
flabel metal3 s -26 1248 -22 1252 7 FreeSans 24 0 0 0 data_memory_interface_address[3]
port 111 nsew
flabel metal2 s 1382 -22 1386 -18 7 FreeSans 24 270 0 0 data_memory_interface_address[4]
port 112 nsew
flabel metal3 s -26 848 -22 852 7 FreeSans 24 0 0 0 data_memory_interface_address[5]
port 113 nsew
flabel metal3 s -26 948 -22 952 7 FreeSans 24 0 0 0 data_memory_interface_address[6]
port 114 nsew
flabel metal2 s 1398 -22 1402 -18 7 FreeSans 24 270 0 0 data_memory_interface_address[7]
port 115 nsew
flabel metal2 s 1126 -22 1130 -18 7 FreeSans 24 270 0 0 data_memory_interface_address[8]
port 116 nsew
flabel metal2 s 1414 -22 1418 -18 7 FreeSans 24 270 0 0 data_memory_interface_address[9]
port 117 nsew
flabel metal2 s 1246 -22 1250 -18 7 FreeSans 24 270 0 0 data_memory_interface_address[10]
port 118 nsew
flabel metal3 s -26 568 -22 572 7 FreeSans 24 0 0 0 data_memory_interface_address[11]
port 119 nsew
flabel metal2 s 230 -22 234 -18 7 FreeSans 24 270 0 0 data_memory_interface_address[12]
port 120 nsew
flabel metal2 s 1366 -22 1370 -18 7 FreeSans 24 270 0 0 data_memory_interface_address[13]
port 121 nsew
flabel metal2 s 1550 -22 1554 -18 7 FreeSans 24 270 0 0 data_memory_interface_address[14]
port 122 nsew
flabel metal2 s 1574 -22 1578 -18 7 FreeSans 24 270 0 0 data_memory_interface_address[15]
port 123 nsew
flabel metal2 s 518 -22 522 -18 7 FreeSans 24 270 0 0 data_memory_interface_address[16]
port 124 nsew
flabel metal2 s 790 -22 794 -18 7 FreeSans 24 270 0 0 data_memory_interface_address[17]
port 125 nsew
flabel metal3 s -26 1188 -22 1192 7 FreeSans 24 0 0 0 data_memory_interface_address[18]
port 126 nsew
flabel metal2 s 1030 -22 1034 -18 7 FreeSans 24 270 0 0 data_memory_interface_address[19]
port 127 nsew
flabel metal3 s -26 1268 -22 1272 7 FreeSans 24 0 0 0 data_memory_interface_address[20]
port 128 nsew
flabel metal3 s -26 1048 -22 1052 7 FreeSans 24 0 0 0 data_memory_interface_address[21]
port 129 nsew
flabel metal3 s -26 1388 -22 1392 7 FreeSans 24 0 0 0 data_memory_interface_address[22]
port 130 nsew
flabel metal3 s -26 1348 -22 1352 7 FreeSans 24 0 0 0 data_memory_interface_address[23]
port 131 nsew
flabel metal3 s -26 1368 -22 1372 7 FreeSans 24 0 0 0 data_memory_interface_address[24]
port 132 nsew
flabel metal3 s -26 2168 -22 2172 7 FreeSans 24 0 0 0 data_memory_interface_address[25]
port 133 nsew
flabel metal3 s -26 2068 -22 2072 7 FreeSans 24 0 0 0 data_memory_interface_address[26]
port 134 nsew
flabel metal3 s -26 2248 -22 2252 7 FreeSans 24 0 0 0 data_memory_interface_address[27]
port 135 nsew
flabel metal3 s -26 1948 -22 1952 7 FreeSans 24 0 0 0 data_memory_interface_address[28]
port 136 nsew
flabel metal3 s -26 2188 -22 2192 7 FreeSans 24 0 0 0 data_memory_interface_address[29]
port 137 nsew
flabel metal3 s -26 1448 -22 1452 7 FreeSans 24 0 0 0 data_memory_interface_address[30]
port 138 nsew
flabel metal3 s -26 1648 -22 1652 7 FreeSans 24 0 0 0 data_memory_interface_address[31]
port 139 nsew
flabel metal2 s 3382 4428 3386 4432 3 FreeSans 24 90 0 0 data_memory_interface_frame_mask[0]
port 140 nsew
flabel metal2 s 3518 4428 3522 4432 3 FreeSans 24 90 0 0 data_memory_interface_frame_mask[1]
port 141 nsew
flabel metal2 s 3406 4428 3410 4432 3 FreeSans 24 90 0 0 data_memory_interface_frame_mask[2]
port 142 nsew
flabel metal2 s 3462 4428 3466 4432 3 FreeSans 24 90 0 0 data_memory_interface_frame_mask[3]
port 143 nsew
<< end >>
