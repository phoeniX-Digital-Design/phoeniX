module Control_Unit 
(
      input [6 : 0] opcode,
      input [2 : 0] funct3,
      input [6 : 0] funct7,
      input [2 : 0] instruction_type,

      input [4 : 0] read_index_1,
      input [4 : 0] read_index_2,
      input [4 : 0] write_index


      // inputs :)))
);
      
endmodule