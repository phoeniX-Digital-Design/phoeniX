module Register_File
#(
    parameter WIDTH = 32,
    parameter DEPTH = 5
)
(
    input CLK,
    input reset,
    
    input wire read_enable_1,
    input wire read_enable_2,
    input wire write_enable,
    
    input wire [DEPTH - 1 : 0] read_index_1,
    input wire [DEPTH - 1 : 0] read_index_2,
    input wire [DEPTH - 1 : 0] write_index,

    input wire [WIDTH - 1 : 0] write_data,

    output reg [WIDTH - 1 : 0] read_data_1,
    output reg [WIDTH - 1 : 0] read_data_2

);
	reg [WIDTH - 1 : 0] Registers [0 : $pow(2, DEPTH) - 1];      

    integer i;    	
    always @(posedge reset)
    begin
        for (i = 0; i < $pow(2, DEPTH) - 1; i = i + 1)
            Registers[i] = {WIDTH{1'b0}};
    end
	
    always @(negedge CLK)
    begin
        if (write_enable == 1'b1 && write_index != 0)
        begin
            Registers[write_index] <= write_data;
        end
    end

    always @(*) 
    begin
        if (read_enable_1 == 1'b1)
            read_data_1 <= Registers[read_index_1];
        else
            read_data_1 <= {WIDTH{1'bz}};

        if (read_enable_2 == 1'b1)
            read_data_2 <= Registers[read_index_2];
        else
            read_data_2 <= {WIDTH{1'bz}};
    end
    
endmodule