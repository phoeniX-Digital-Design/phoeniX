
module phoeniX ( clk, reset, instruction_memory_interface_enable, 
        instruction_memory_interface_state, 
        instruction_memory_interface_address, 
        instruction_memory_interface_frame_mask, 
        instruction_memory_interface_data, data_memory_interface_enable, 
        data_memory_interface_state, data_memory_interface_address, 
        data_memory_interface_frame_mask, data_memory_interface_data );
  output [31:0] instruction_memory_interface_address;
  output [3:0] instruction_memory_interface_frame_mask;
  input [31:0] instruction_memory_interface_data;
  output [31:0] data_memory_interface_address;
  output [3:0] data_memory_interface_frame_mask;
  inout [31:0] data_memory_interface_data;
  input clk, reset;
  output instruction_memory_interface_enable,
         instruction_memory_interface_state, data_memory_interface_enable,
         data_memory_interface_state;
  wire   _0_net_, jump_branch_enable_EX_wire, N193, N197, N198, N200, N201,
         N203, N204, N206, N207, N209, N210, N212, N213, N215, N216, N218,
         N219, N221, N222, N224, N225, N227, N228, N230, N231, N233, N234,
         N236, N237, N239, N240, N242, N243, N245, N246, N248, N249, N251,
         N252, N254, N255, N257, N258, N260, N261, N263, N264, N266, N267,
         N269, N270, N272, N273, N275, N276, N278, N279, N281, N282, N284,
         N285, N287, N288, N290, N291, read_enable_1_FD_wire,
         read_enable_2_FD_wire, write_enable_FD_wire, read_enable_csr_FD_wire,
         write_enable_csr_FD_wire, FW_enable_1, FW_enable_2,
         write_enable_EX_reg, write_enable_csr_EX_reg, N370, N371, N373, N374,
         N376, N377, N379, N380, N382, N383, N385, N386, N388, N389, N391,
         N392, N394, N395, N397, N398, N400, N401, N403, N404, N406, N407,
         N409, N410, N412, N413, N415, N416, N418, N419, N421, N422, N424,
         N425, N427, N428, N430, N431, N433, N434, N436, N437, N439, N440,
         N442, N443, N445, N446, N448, N449, N451, N452, N454, N455, N457,
         N458, N460, N461, N463, N464, N466, N467, N469, N470, N472, N473,
         N475, N476, N478, N479, N481, N482, N484, N485, N487, N488, N490,
         N491, N493, N494, N496, N497, N499, N500, N502, N503, N505, N506,
         N508, N509, N511, N512, N514, N515, N517, N518, N520, N521, N523,
         N524, N526, N527, N529, N530, N532, N533, N535, N536, N538, N539,
         N541, N542, N544, N545, N547, N548, N550, N551, N553, N554, N556,
         N557, N559, N560, mul_busy_EX_wire, write_enable_MW_reg, N651, N654,
         N655, N656, N657, N658, N659, N660, N661, N662, N663, N664, N665,
         N666, N667, N668, N669, N670, N671, N672, N673, N674, N675, N676,
         N677, N678, N679, N680, N681, N682, N683, N684, N685, N686, N687,
         N688, N689, N690, N691, N692, N693, N694, N695, N696, N697, N698,
         N699, N700, N701, N702, N703, N704, N705, N706, N707, N708, N709,
         N710, N711, N712, N713, N714, N715, N716, N717, \_2_net_[30] ,
         \_2_net_[29] , \_2_net_[28] , \_2_net_[27] , \_2_net_[26] ,
         \_2_net_[25] , \_2_net_[24] , \_2_net_[23] , \_2_net_[22] ,
         \_2_net_[21] , \_2_net_[20] , \_2_net_[19] , \_2_net_[18] ,
         \_2_net_[17] , \_2_net_[16] , \_2_net_[15] , \_2_net_[14] ,
         \_2_net_[13] , \_2_net_[12] , \_2_net_[11] , \_2_net_[10] ,
         \_2_net_[9] , \_2_net_[8] , \_2_net_[7] , \_2_net_[6] , \_2_net_[5] ,
         \_2_net_[4] , \_2_net_[3] , \_2_net_[2] , \_2_net_[1] , \_2_net_[0] ,
         n1, n3, n4, n5, n6, n7, n8, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n22, n23, n25, n26, n27, n28, n29, n30, n31, n32, n36,
         n37, n38, n39, n40, n66, n67, n69, n70, n71, n76, n77, n78, n79, n80,
         n82, n83, n84, n86, n87, n88, n90, n91, n92, n94, n95, n96, n98, n99,
         n100, n102, n103, n104, n106, n107, n108, n110, n111, n112, n114,
         n115, n116, n118, n119, n120, n122, n123, n124, n126, n127, n128,
         n130, n131, n132, n134, n135, n136, n138, n139, n140, n142, n143,
         n144, n146, n147, n148, n150, n151, n152, n154, n155, n156, n158,
         n159, n160, n162, n163, n164, n166, n167, n168, n170, n171, n172,
         n174, n175, n176, n178, n179, n180, n182, n183, n184, n186, n187,
         n188, n190, n191, n192, n194, n195, n196, n198, n199, n200, n201,
         n202, n203, n204, n205, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n595, n596, n597, n599, n601, n603,
         n605, n607, n609, n611, n613, n615, n617, n619, n621, n623, n625,
         n627, n629, n631, n633, n635, n637, n639, n641, n643, n645, n647,
         n649, n651, n653, n655, n657, n787, n788, n789, n790, n792, n795,
         n798, n801, n804, n807, n810, n813, n816, n819, n822, n825, n828,
         n831, n834, n837, n840, n843, n846, n849, n852, n855, n858, n861,
         n864, n867, n870, n873, n876, n879, n882, n885, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1156, n1157, n1158, n1159, n1160,
         n1161, n1163, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1214, n1215, n1216, n1218,
         n1219, n1220, n1221, n1222, n1223, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1234, n1235, n1240, n1241, n1244, n1246, n1247,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1284,
         n1285, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1356, n1360,
         n1361, n1362, n1364, n1366, n1368, n1370, n1372, n1374, n1376, n1378,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1443,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1480, n1481, n1482, n1483, n1484, n1485,
         n1488, n1494, n1559, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1245, n1827,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2004, n2005, n2006, n2007, n2008, n2009, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2055, n2056, n2057, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2077, n2079, n2080, n2081, n2085, n2086, n2087, n2090, n2091, n2092,
         n2093, n2094, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509;
  wire   [31:0] pc_FD_reg;
  wire   [6:0] opcode_EX_reg;
  wire   [2:0] funct3_EX_reg;
  wire   [6:0] funct7_EX_reg;
  wire   [11:0] funct12_EX_reg;
  wire   [31:0] immediate_EX_reg;
  wire   [2:0] instruction_type_EX_reg;
  wire   [4:0] write_index_EX_reg;
  wire   [31:0] pc_EX_reg;
  wire   [31:0] next_pc_EX_reg;
  wire   [11:0] csr_index_EX_reg;
  wire   [31:0] csr_data_EX_reg;
  wire   [4:0] read_index_1_EX_reg;
  wire   [31:0] alucsr_wire;
  wire   [31:0] mulcsr_wire;
  wire   [31:0] divcsr_wire;
  wire   [6:0] opcode_MW_reg;
  wire   [2:0] funct3_MW_reg;
  wire   [6:0] funct7_MW_reg;
  wire   [11:0] funct12_MW_reg;
  wire   [31:0] immediate_MW_reg;
  wire   [4:0] write_index_MW_reg;
  wire   [31:0] address_MW_reg;
  wire   [31:0] rs2_MW_reg;
  wire   [31:0] execution_result_MW_reg;
  wire   [31:0] csr_rd_MW_reg;
  tri   instruction_memory_interface_state;
  tri   [31:0] instruction_memory_interface_address;
  tri   [3:0] instruction_memory_interface_frame_mask;
  tri   data_memory_interface_state;
  tri   [31:0] data_memory_interface_address;
  tri   [3:0] data_memory_interface_frame_mask;
  tri   [31:0] data_memory_interface_data;
  tri   [31:0] next_pc_FD_wire;
  tri   [31:0] address_EX_wire;
  tri   [31:0] instruction_FD_reg;
  tri   [2:0] instruction_type_FD_wire;
  tri   [6:0] opcode_FD_wire;
  tri   [2:0] funct3_FD_wire;
  tri   [6:0] funct7_FD_wire;
  tri   [11:0] funct12_FD_wire;
  tri   [4:0] read_index_1_FD_wire;
  tri   [4:0] read_index_2_FD_wire;
  tri   [4:0] write_index_FD_wire;
  tri   [11:0] csr_index_FD_wire;
  tri   [31:0] immediate_FD_wire;
  tri   [31:0] FW_source_1;
  tri   [31:0] RF_source_1;
  tri   [31:0] FW_source_2;
  tri   [31:0] RF_source_2;
  tri   [31:0] rs1_EX_reg;
  tri   [31:0] rs2_EX_reg;
  tri   [31:0] csr_data_FD_wire;
  tri   [31:0] alu_output_EX_wire;
  tri   [31:0] mul_output_EX_wire;
  tri   [31:0] div_output_EX_wire;
  tri   [31:0] csr_rd_EX_wire;
  tri   [31:0] csr_data_out_EX_wire;
  tri   [31:0] load_data_MW_wire;
  tri   [31:0] write_data_MW_reg;
  tri   n2010;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74;

  Fetch_Unit fetch_unit ( .enable(_0_net_), .pc(pc_FD_reg), .next_pc(
        next_pc_FD_wire), .memory_interface_enable(
        instruction_memory_interface_enable), .memory_interface_state(
        instruction_memory_interface_state), .memory_interface_address(
        instruction_memory_interface_address), .memory_interface_frame_mask(
        instruction_memory_interface_frame_mask) );
  Instruction_Decoder instruction_decoder ( .instruction(instruction_FD_reg), 
        .instruction_type(instruction_type_FD_wire), .opcode(opcode_FD_wire), 
        .funct3(funct3_FD_wire), .funct7(funct7_FD_wire), .funct12(
        funct12_FD_wire), .read_index_1(read_index_1_FD_wire), .read_index_2(
        read_index_2_FD_wire), .write_index(write_index_FD_wire), .csr_index(
        csr_index_FD_wire), .read_enable_1(read_enable_1_FD_wire), 
        .read_enable_2(read_enable_2_FD_wire), .write_enable(
        write_enable_FD_wire), .read_enable_csr(read_enable_csr_FD_wire), 
        .write_enable_csr(write_enable_csr_FD_wire) );
  Immediate_Generator immediate_generator ( .instruction(
        instruction_FD_reg[31:7]), .instruction_type(instruction_type_FD_wire), 
        .immediate(immediate_FD_wire) );
  Arithmetic_Logic_Unit_GENERATE_CIRCUIT_11_GENERATE_CIRCUIT_20_GENERATE_CIRCUIT_30_GENERATE_CIRCUIT_40 arithmetic_logic_unit ( 
        .opcode({n2154, n2414, n2415, n2077, n2072, opcode_EX_reg[1:0]}), 
        .funct3({funct3_EX_reg[2], n2474, funct3_EX_reg[0]}), .funct7(
        funct7_EX_reg), .control_status_register({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, alucsr_wire[10:8], 1'b0, alucsr_wire[6:0]}), 
        .rs1({rs1_EX_reg[31:1], n2062}), .rs2(rs2_EX_reg), .immediate(
        immediate_EX_reg), .alu_output(alu_output_EX_wire) );
  Multiplier_Unit_GENERATE_CIRCUIT_11_GENERATE_CIRCUIT_20_GENERATE_CIRCUIT_30_GENERATE_CIRCUIT_40 \M_EXTENSION_Generate_Block.multiplier_unit  ( 
        .clk(clk), .opcode({n2154, n2414, n2415, opcode_EX_reg[3], n2072, 
        opcode_EX_reg[1:0]}), .funct7(funct7_EX_reg), .funct3({
        funct3_EX_reg[2], n2474, funct3_EX_reg[0]}), .control_status_register(
        {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        mulcsr_wire[9:4], 1'b0, mulcsr_wire[2:0]}), .rs1({rs1_EX_reg[31:1], 
        n2062}), .rs2(rs2_EX_reg), .multiplier_unit_busy(mul_busy_EX_wire), 
        .multiplier_unit_output(mul_output_EX_wire) );
  Divider_Unit_GENERATE_CIRCUIT_11_GENERATE_CIRCUIT_20_GENERATE_CIRCUIT_30_GENERATE_CIRCUIT_40 \M_EXTENSION_Generate_Block.divider_unit  ( 
        .clk(clk), .opcode({n2154, n2414, n2415, n2077, n2072, 
        opcode_EX_reg[1:0]}), .funct7(funct7_EX_reg), .funct3({
        funct3_EX_reg[2], n2474, 1'b0}), .control_status_register({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, divcsr_wire[2:1], 1'b0}), .rs1({rs1_EX_reg[31:1], 
        n2062}), .rs2(rs2_EX_reg), .divider_unit_busy(n2012), 
        .divider_unit_output(div_output_EX_wire) );
  Address_Generator address_generator ( .opcode(opcode_EX_reg), .rs1(
        rs1_EX_reg), .pc(pc_EX_reg), .immediate(immediate_EX_reg), .address({
        address_EX_wire[31:17], n2010, address_EX_wire[15:0]}) );
  Jump_Branch_Unit jump_branch_unit ( .opcode({n2154, n2414, n2415, 1'b0, 
        n2072, opcode_EX_reg[1:0]}), .funct3({funct3_EX_reg[2], n2474, 
        funct3_EX_reg[0]}), .instruction_type(instruction_type_EX_reg), .rs1(
        rs1_EX_reg), .rs2(rs2_EX_reg), .jump_branch_enable(
        jump_branch_enable_EX_wire) );
  Control_Status_Unit control_status_unit ( .opcode({n2154, n2414, n2415, 
        n2077, n2072, opcode_EX_reg[1:0]}), .funct3({funct3_EX_reg[2], n2474, 
        funct3_EX_reg[0]}), .CSR_in(csr_data_EX_reg), .rs1(rs1_EX_reg), 
        .unsigned_immediate(read_index_1_EX_reg), .rd(csr_rd_EX_wire), 
        .CSR_out(csr_data_out_EX_wire) );
  Load_Store_Unit load_store_unit ( .opcode(opcode_MW_reg), .funct3(
        funct3_MW_reg), .address(address_MW_reg), .store_data(rs2_MW_reg), 
        .load_data(load_data_MW_wire), .memory_interface_enable(
        data_memory_interface_enable), .memory_interface_state(
        data_memory_interface_state), .memory_interface_address(
        data_memory_interface_address), .memory_interface_frame_mask(
        data_memory_interface_frame_mask), .memory_interface_data(
        data_memory_interface_data) );
  Hazard_Forward_Unit_1 hazard_forward_unit_source_1 ( .source_index(
        read_index_1_FD_wire), .destination_index_1(write_index_EX_reg), 
        .destination_index_2(write_index_MW_reg), .data_1({n1910, 
        \_2_net_[30] , \_2_net_[29] , \_2_net_[28] , \_2_net_[27] , 
        \_2_net_[26] , \_2_net_[25] , \_2_net_[24] , \_2_net_[23] , n2055, 
        n1832, \_2_net_[20] , \_2_net_[19] , \_2_net_[18] , \_2_net_[17] , 
        \_2_net_[16] , \_2_net_[15] , \_2_net_[14] , \_2_net_[13] , 
        \_2_net_[12] , \_2_net_[11] , \_2_net_[10] , \_2_net_[9] , 
        \_2_net_[8] , \_2_net_[7] , \_2_net_[6] , \_2_net_[5] , \_2_net_[4] , 
        \_2_net_[3] , \_2_net_[2] , \_2_net_[1] , \_2_net_[0] }), .data_2(
        write_data_MW_reg), .enable_1(write_enable_EX_reg), .enable_2(
        write_enable_MW_reg), .forward_enable(FW_enable_1), .forward_data(
        FW_source_1) );
  Hazard_Forward_Unit_0 hazard_forward_unit_source_2 ( .source_index(
        read_index_2_FD_wire), .destination_index_1(write_index_EX_reg), 
        .destination_index_2(write_index_MW_reg), .data_1({n1910, 
        \_2_net_[30] , \_2_net_[29] , \_2_net_[28] , \_2_net_[27] , 
        \_2_net_[26] , \_2_net_[25] , \_2_net_[24] , \_2_net_[23] , 
        \_2_net_[22] , \_2_net_[21] , \_2_net_[20] , \_2_net_[19] , 
        \_2_net_[18] , \_2_net_[17] , \_2_net_[16] , \_2_net_[15] , 
        \_2_net_[14] , \_2_net_[13] , \_2_net_[12] , \_2_net_[11] , 
        \_2_net_[10] , \_2_net_[9] , \_2_net_[8] , \_2_net_[7] , \_2_net_[6] , 
        \_2_net_[5] , \_2_net_[4] , \_2_net_[3] , \_2_net_[2] , \_2_net_[1] , 
        \_2_net_[0] }), .data_2(write_data_MW_reg), .enable_1(
        write_enable_EX_reg), .enable_2(write_enable_MW_reg), .forward_enable(
        FW_enable_2), .forward_data(FW_source_2) );
  Register_File_WIDTH32_DEPTH5 register_file ( .clk(clk), .read_enable_1(
        read_enable_1_FD_wire), .read_enable_2(read_enable_2_FD_wire), 
        .write_enable(write_enable_MW_reg), .read_index_1(read_index_1_FD_wire), .read_index_2(read_index_2_FD_wire), .write_index(write_index_MW_reg), 
        .write_data(write_data_MW_reg), .read_data_1(RF_source_1), 
        .read_data_2(RF_source_2), .reset_BAR(n2475) );
  Control_Status_Register_File control_status_register_file ( .clk(clk), 
        .opcode(opcode_MW_reg), .funct3(funct3_MW_reg), .funct7(funct7_MW_reg), 
        .funct12(funct12_MW_reg), .write_index(write_index_MW_reg), 
        .read_enable_csr(read_enable_csr_FD_wire), .write_enable_csr(
        write_enable_csr_EX_reg), .csr_read_index(csr_index_FD_wire), 
        .csr_write_index(csr_index_EX_reg), .csr_write_data(
        csr_data_out_EX_wire), .csr_read_data(csr_data_FD_wire), .alucsr_wire(
        {SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, alucsr_wire[10:8], SYNOPSYS_UNCONNECTED__21, 
        alucsr_wire[6:0]}), .mulcsr_wire({SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, mulcsr_wire[9:4], SYNOPSYS_UNCONNECTED__44, 
        mulcsr_wire[2:0]}), .divcsr_wire({SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, divcsr_wire[2:1], 
        SYNOPSYS_UNCONNECTED__74}), .reset_BAR(n2475) );
  DFF_X1 \rs2_MW_reg_reg[0]  ( .D(n1123), .CK(clk), .Q(rs2_MW_reg[0]), .QN(
        n211) );
  DFF_X1 \rs2_MW_reg_reg[31]  ( .D(n1122), .CK(clk), .Q(rs2_MW_reg[31]), .QN(
        n212) );
  DFF_X1 \execution_result_MW_reg_reg[31]  ( .D(n1611), .CK(clk), .Q(
        execution_result_MW_reg[31]), .QN(n1176) );
  DFF_X1 \execution_result_MW_reg_reg[0]  ( .D(n1580), .CK(clk), .Q(
        execution_result_MW_reg[0]), .QN(n1207) );
  DFF_X1 \rs1_EX_reg_reg[30]  ( .D(n1418), .CK(clk), .Q(), .QN(N373) );
  DFF_X1 \rs2_EX_reg_reg[0]  ( .D(n1421), .CK(clk), .Q(), .QN(N559) );
  DFF_X1 \rs2_EX_reg_reg[1]  ( .D(n1425), .CK(clk), .Q(), .QN(N556) );
  DFF_X1 \rs2_EX_reg_reg[2]  ( .D(n1427), .CK(clk), .Q(), .QN(N553) );
  DFF_X1 \rs2_EX_reg_reg[3]  ( .D(n1429), .CK(clk), .Q(), .QN(N550) );
  DFF_X1 \rs2_EX_reg_reg[4]  ( .D(n1431), .CK(clk), .Q(), .QN(N547) );
  DFF_X1 \rs2_EX_reg_reg[6]  ( .D(n1435), .CK(clk), .Q(), .QN(N541) );
  DFF_X1 \rs2_EX_reg_reg[7]  ( .D(n1437), .CK(clk), .Q(), .QN(N538) );
  DFF_X1 \rs2_EX_reg_reg[8]  ( .D(n1439), .CK(clk), .Q(), .QN(N535) );
  DFF_X1 \rs2_EX_reg_reg[9]  ( .D(n1441), .CK(clk), .Q(), .QN(N532) );
  DFF_X1 \rs2_EX_reg_reg[11]  ( .D(n1445), .CK(clk), .Q(), .QN(N526) );
  DFF_X1 \rs2_EX_reg_reg[12]  ( .D(n1447), .CK(clk), .Q(), .QN(N523) );
  DFF_X1 \rs2_EX_reg_reg[13]  ( .D(n1449), .CK(clk), .Q(), .QN(N520) );
  DFF_X1 \rs2_EX_reg_reg[14]  ( .D(n1451), .CK(clk), .Q(), .QN(N517) );
  DFF_X1 \rs2_EX_reg_reg[15]  ( .D(n1453), .CK(clk), .Q(), .QN(N514) );
  DFF_X1 \rs2_EX_reg_reg[17]  ( .D(n1457), .CK(clk), .Q(), .QN(N508) );
  DFF_X1 \rs2_EX_reg_reg[18]  ( .D(n1459), .CK(clk), .Q(), .QN(N505) );
  DFF_X1 \rs2_EX_reg_reg[20]  ( .D(n1463), .CK(clk), .Q(), .QN(N499) );
  DFF_X1 \rs2_EX_reg_reg[21]  ( .D(n1465), .CK(clk), .Q(), .QN(N496) );
  DFF_X1 \rs2_EX_reg_reg[22]  ( .D(n1467), .CK(clk), .Q(), .QN(N493) );
  DFF_X1 \rs2_EX_reg_reg[25]  ( .D(n1473), .CK(clk), .Q(), .QN(N484) );
  DFF_X1 \rs2_EX_reg_reg[26]  ( .D(n1475), .CK(clk), .Q(), .QN(N481) );
  DFF_X1 \rs2_EX_reg_reg[27]  ( .D(n1477), .CK(clk), .Q(), .QN(N478) );
  DFF_X1 \rs2_EX_reg_reg[29]  ( .D(n1481), .CK(clk), .Q(), .QN(N472) );
  DFF_X1 \rs2_EX_reg_reg[30]  ( .D(n1483), .CK(clk), .Q(), .QN(N469) );
  DFF_X1 \rs1_EX_reg_reg[0]  ( .D(n1356), .CK(clk), .Q(), .QN(N463) );
  DFF_X1 \rs1_EX_reg_reg[1]  ( .D(n1360), .CK(clk), .Q(), .QN(N460) );
  DFF_X1 \rs1_EX_reg_reg[2]  ( .D(n1362), .CK(clk), .Q(), .QN(N457) );
  DFF_X1 \rs1_EX_reg_reg[4]  ( .D(n1366), .CK(clk), .Q(), .QN(N451) );
  DFF_X1 \rs1_EX_reg_reg[6]  ( .D(n1370), .CK(clk), .Q(), .QN(N445) );
  DFF_X1 \rs1_EX_reg_reg[7]  ( .D(n1372), .CK(clk), .Q(), .QN(N442) );
  DFF_X1 \rs1_EX_reg_reg[8]  ( .D(n1374), .CK(clk), .Q(), .QN(N439) );
  DFF_X1 \rs1_EX_reg_reg[9]  ( .D(n1376), .CK(clk), .Q(), .QN(N436) );
  DFF_X1 \rs1_EX_reg_reg[10]  ( .D(n1378), .CK(clk), .Q(), .QN(N433) );
  DFF_X1 \rs1_EX_reg_reg[11]  ( .D(n1380), .CK(clk), .Q(), .QN(N430) );
  DFF_X1 \rs1_EX_reg_reg[12]  ( .D(n1382), .CK(clk), .Q(), .QN(N427) );
  DFF_X1 \rs1_EX_reg_reg[13]  ( .D(n1384), .CK(clk), .Q(), .QN(N424) );
  DFF_X1 \rs1_EX_reg_reg[14]  ( .D(n1386), .CK(clk), .Q(), .QN(N421) );
  DFF_X1 \rs1_EX_reg_reg[15]  ( .D(n1388), .CK(clk), .Q(), .QN(N418) );
  DFF_X1 \rs1_EX_reg_reg[17]  ( .D(n1392), .CK(clk), .Q(), .QN(N412) );
  DFF_X1 \rs1_EX_reg_reg[18]  ( .D(n1394), .CK(clk), .Q(), .QN(N409) );
  DFF_X1 \rs1_EX_reg_reg[20]  ( .D(n1398), .CK(clk), .Q(), .QN(N403) );
  DFF_X1 \rs1_EX_reg_reg[21]  ( .D(n1400), .CK(clk), .Q(), .QN(N400) );
  DFF_X1 \rs1_EX_reg_reg[22]  ( .D(n1402), .CK(clk), .Q(), .QN(N397) );
  DFF_X1 \rs1_EX_reg_reg[25]  ( .D(n1408), .CK(clk), .Q(), .QN(N388) );
  DFF_X1 \rs1_EX_reg_reg[26]  ( .D(n1410), .CK(clk), .Q(), .QN(N385) );
  DFF_X1 \rs1_EX_reg_reg[27]  ( .D(n1412), .CK(clk), .Q(), .QN(N382) );
  DFF_X1 \rs1_EX_reg_reg[29]  ( .D(n1416), .CK(clk), .Q(), .QN(N376) );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[0]  ( .D(n1762), .CK(clk), .Q(N464), .QN()
         );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[1]  ( .D(n1763), .CK(clk), .Q(N461), .QN()
         );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[2]  ( .D(n1764), .CK(clk), .Q(N458), .QN()
         );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[3]  ( .D(n1765), .CK(clk), .Q(N455), .QN()
         );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[4]  ( .D(n1766), .CK(clk), .Q(N452), .QN()
         );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[5]  ( .D(n1767), .CK(clk), .Q(N449), .QN()
         );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[6]  ( .D(n1768), .CK(clk), .Q(N446), .QN()
         );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[7]  ( .D(n1769), .CK(clk), .Q(N443), .QN()
         );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[8]  ( .D(n1770), .CK(clk), .Q(N440), .QN()
         );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[9]  ( .D(n1771), .CK(clk), .Q(N437), .QN()
         );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[10]  ( .D(n1772), .CK(clk), .Q(N434), .QN(
        n2085) );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[11]  ( .D(n1773), .CK(clk), .Q(N431), 
        .QN() );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[12]  ( .D(n1774), .CK(clk), .Q(N428), 
        .QN() );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[13]  ( .D(n1775), .CK(clk), .Q(N425), 
        .QN() );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[14]  ( .D(n1776), .CK(clk), .Q(N422), 
        .QN() );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[15]  ( .D(n1777), .CK(clk), .Q(N419), 
        .QN() );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[16]  ( .D(n1778), .CK(clk), .Q(N416), 
        .QN() );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[17]  ( .D(n1779), .CK(clk), .Q(N413), 
        .QN() );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[18]  ( .D(n1780), .CK(clk), .Q(N410), 
        .QN() );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[19]  ( .D(n1781), .CK(clk), .Q(N407), 
        .QN() );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[20]  ( .D(n1782), .CK(clk), .Q(N404), 
        .QN() );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[21]  ( .D(n1783), .CK(clk), .Q(N401), 
        .QN() );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[22]  ( .D(n1784), .CK(clk), .Q(N398), 
        .QN() );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[23]  ( .D(n1785), .CK(clk), .Q(N395), 
        .QN() );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[24]  ( .D(n1786), .CK(clk), .Q(N392), 
        .QN() );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[25]  ( .D(n1787), .CK(clk), .Q(N389), 
        .QN() );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[26]  ( .D(n1788), .CK(clk), .Q(N386), 
        .QN() );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[27]  ( .D(n1789), .CK(clk), .Q(N383), 
        .QN() );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[28]  ( .D(n1790), .CK(clk), .Q(N380), 
        .QN() );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[29]  ( .D(n1791), .CK(clk), .Q(N377), 
        .QN() );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[30]  ( .D(n1792), .CK(clk), .Q(N374), 
        .QN() );
  DFF_X1 \rs1_EX_reg_tri_enable_reg[31]  ( .D(n1793), .CK(clk), .Q(N371), 
        .QN() );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[0]  ( .D(n1794), .CK(clk), .Q(N560), .QN()
         );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[1]  ( .D(n1795), .CK(clk), .Q(N557), .QN()
         );
  DFF_X1 \rs2_MW_reg_reg[1]  ( .D(n1121), .CK(clk), .Q(rs2_MW_reg[1]), .QN(
        n213) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[2]  ( .D(n1796), .CK(clk), .Q(N554), .QN()
         );
  DFF_X1 \rs2_MW_reg_reg[2]  ( .D(n1120), .CK(clk), .Q(rs2_MW_reg[2]), .QN(
        n214) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[3]  ( .D(n1797), .CK(clk), .Q(N551), .QN()
         );
  DFF_X1 \rs2_MW_reg_reg[3]  ( .D(n1119), .CK(clk), .Q(rs2_MW_reg[3]), .QN(
        n215) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[4]  ( .D(n1798), .CK(clk), .Q(N548), .QN()
         );
  DFF_X1 \rs2_MW_reg_reg[4]  ( .D(n1118), .CK(clk), .Q(rs2_MW_reg[4]), .QN(
        n216) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[5]  ( .D(n1799), .CK(clk), .Q(N545), .QN()
         );
  DFF_X1 \rs2_MW_reg_reg[5]  ( .D(n1117), .CK(clk), .Q(rs2_MW_reg[5]), .QN(
        n217) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[6]  ( .D(n1800), .CK(clk), .Q(N542), .QN()
         );
  DFF_X1 \rs2_MW_reg_reg[6]  ( .D(n1116), .CK(clk), .Q(rs2_MW_reg[6]), .QN(
        n218) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[7]  ( .D(n1801), .CK(clk), .Q(N539), .QN()
         );
  DFF_X1 \rs2_MW_reg_reg[7]  ( .D(n1115), .CK(clk), .Q(rs2_MW_reg[7]), .QN(
        n219) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[8]  ( .D(n1802), .CK(clk), .Q(N536), .QN()
         );
  DFF_X1 \rs2_MW_reg_reg[8]  ( .D(n1114), .CK(clk), .Q(rs2_MW_reg[8]), .QN(
        n220) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[9]  ( .D(n1803), .CK(clk), .Q(N533), .QN()
         );
  DFF_X1 \rs2_MW_reg_reg[9]  ( .D(n1113), .CK(clk), .Q(rs2_MW_reg[9]), .QN(
        n221) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[10]  ( .D(n1804), .CK(clk), .Q(N530), 
        .QN() );
  DFF_X1 \rs2_MW_reg_reg[10]  ( .D(n1112), .CK(clk), .Q(rs2_MW_reg[10]), .QN(
        n222) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[11]  ( .D(n1805), .CK(clk), .Q(N527), 
        .QN() );
  DFF_X1 \rs2_MW_reg_reg[11]  ( .D(n1111), .CK(clk), .Q(rs2_MW_reg[11]), .QN(
        n223) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[12]  ( .D(n1806), .CK(clk), .Q(N524), 
        .QN() );
  DFF_X1 \rs2_MW_reg_reg[12]  ( .D(n1110), .CK(clk), .Q(rs2_MW_reg[12]), .QN(
        n224) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[13]  ( .D(n1807), .CK(clk), .Q(N521), 
        .QN() );
  DFF_X1 \rs2_MW_reg_reg[13]  ( .D(n1109), .CK(clk), .Q(rs2_MW_reg[13]), .QN(
        n225) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[14]  ( .D(n1808), .CK(clk), .Q(N518), 
        .QN() );
  DFF_X1 \rs2_MW_reg_reg[14]  ( .D(n1108), .CK(clk), .Q(rs2_MW_reg[14]), .QN(
        n226) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[15]  ( .D(n1809), .CK(clk), .Q(N515), 
        .QN() );
  DFF_X1 \rs2_MW_reg_reg[15]  ( .D(n1107), .CK(clk), .Q(rs2_MW_reg[15]), .QN(
        n227) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[16]  ( .D(n1810), .CK(clk), .Q(N512), 
        .QN() );
  DFF_X1 \rs2_MW_reg_reg[16]  ( .D(n1106), .CK(clk), .Q(rs2_MW_reg[16]), .QN(
        n228) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[17]  ( .D(n1811), .CK(clk), .Q(N509), 
        .QN() );
  DFF_X1 \rs2_MW_reg_reg[17]  ( .D(n1105), .CK(clk), .Q(rs2_MW_reg[17]), .QN(
        n229) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[18]  ( .D(n1812), .CK(clk), .Q(N506), 
        .QN() );
  DFF_X1 \rs2_MW_reg_reg[18]  ( .D(n1104), .CK(clk), .Q(rs2_MW_reg[18]), .QN(
        n230) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[19]  ( .D(n1813), .CK(clk), .Q(N503), 
        .QN() );
  DFF_X1 \rs2_MW_reg_reg[19]  ( .D(n1103), .CK(clk), .Q(rs2_MW_reg[19]), .QN(
        n231) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[20]  ( .D(n1814), .CK(clk), .Q(N500), 
        .QN() );
  DFF_X1 \rs2_MW_reg_reg[20]  ( .D(n1102), .CK(clk), .Q(rs2_MW_reg[20]), .QN(
        n232) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[21]  ( .D(n1815), .CK(clk), .Q(N497), 
        .QN() );
  DFF_X1 \rs2_MW_reg_reg[21]  ( .D(n1101), .CK(clk), .Q(rs2_MW_reg[21]), .QN(
        n233) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[22]  ( .D(n1816), .CK(clk), .Q(N494), 
        .QN() );
  DFF_X1 \rs2_MW_reg_reg[22]  ( .D(n1100), .CK(clk), .Q(rs2_MW_reg[22]), .QN(
        n234) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[23]  ( .D(n1817), .CK(clk), .Q(N491), 
        .QN() );
  DFF_X1 \rs2_MW_reg_reg[23]  ( .D(n1099), .CK(clk), .Q(rs2_MW_reg[23]), .QN(
        n235) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[24]  ( .D(n1818), .CK(clk), .Q(N488), 
        .QN() );
  DFF_X1 \rs2_MW_reg_reg[24]  ( .D(n1098), .CK(clk), .Q(rs2_MW_reg[24]), .QN(
        n236) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[25]  ( .D(n1819), .CK(clk), .Q(N485), 
        .QN() );
  DFF_X1 \rs2_MW_reg_reg[25]  ( .D(n1097), .CK(clk), .Q(rs2_MW_reg[25]), .QN(
        n237) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[26]  ( .D(n1820), .CK(clk), .Q(N482), 
        .QN() );
  DFF_X1 \rs2_MW_reg_reg[26]  ( .D(n1096), .CK(clk), .Q(rs2_MW_reg[26]), .QN(
        n238) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[27]  ( .D(n1821), .CK(clk), .Q(N479), 
        .QN() );
  DFF_X1 \rs2_MW_reg_reg[27]  ( .D(n1095), .CK(clk), .Q(rs2_MW_reg[27]), .QN(
        n239) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[28]  ( .D(n1822), .CK(clk), .Q(N476), 
        .QN() );
  DFF_X1 \rs2_MW_reg_reg[28]  ( .D(n1094), .CK(clk), .Q(rs2_MW_reg[28]), .QN(
        n240) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[29]  ( .D(n1823), .CK(clk), .Q(N473), 
        .QN() );
  DFF_X1 \rs2_MW_reg_reg[29]  ( .D(n1093), .CK(clk), .Q(rs2_MW_reg[29]), .QN(
        n241) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[30]  ( .D(n1824), .CK(clk), .Q(N470), 
        .QN() );
  DFF_X1 \rs2_MW_reg_reg[30]  ( .D(n1092), .CK(clk), .Q(rs2_MW_reg[30]), .QN(
        n242) );
  DFF_X1 \rs2_EX_reg_tri_enable_reg[31]  ( .D(n1825), .CK(clk), .Q(N467), 
        .QN() );
  DLH_X1 \instruction_FD_reg_reg[31]  ( .G(N193), .D(
        instruction_memory_interface_data[31]), .Q(N197) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[31]  ( .G(N193), .D(reset), .Q(
        N198) );
  DLH_X1 \instruction_FD_reg_reg[30]  ( .G(N193), .D(
        instruction_memory_interface_data[30]), .Q(N200) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[30]  ( .G(N193), .D(reset), .Q(
        N201) );
  DLH_X1 \instruction_FD_reg_reg[29]  ( .G(N193), .D(
        instruction_memory_interface_data[29]), .Q(N203) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[29]  ( .G(N193), .D(reset), .Q(
        N204) );
  DLH_X1 \instruction_FD_reg_reg[28]  ( .G(N193), .D(
        instruction_memory_interface_data[28]), .Q(N206) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[28]  ( .G(N193), .D(reset), .Q(
        N207) );
  DLH_X1 \instruction_FD_reg_reg[27]  ( .G(N193), .D(
        instruction_memory_interface_data[27]), .Q(N209) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[27]  ( .G(N193), .D(n2476), .Q(
        N210) );
  DLH_X1 \instruction_FD_reg_reg[26]  ( .G(N193), .D(
        instruction_memory_interface_data[26]), .Q(N212) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[26]  ( .G(N193), .D(n2476), .Q(
        N213) );
  DLH_X1 \instruction_FD_reg_reg[25]  ( .G(N193), .D(
        instruction_memory_interface_data[25]), .Q(N215) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[25]  ( .G(N193), .D(n2476), .Q(
        N216) );
  DLH_X1 \instruction_FD_reg_reg[24]  ( .G(N193), .D(
        instruction_memory_interface_data[24]), .Q(N218) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[24]  ( .G(N193), .D(n2476), .Q(
        N219) );
  DLH_X1 \instruction_FD_reg_reg[23]  ( .G(N193), .D(
        instruction_memory_interface_data[23]), .Q(N221) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[23]  ( .G(N193), .D(n2476), .Q(
        N222) );
  DLH_X1 \instruction_FD_reg_reg[22]  ( .G(N193), .D(
        instruction_memory_interface_data[22]), .Q(N224) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[22]  ( .G(N193), .D(n2476), .Q(
        N225) );
  DLH_X1 \instruction_FD_reg_reg[21]  ( .G(N193), .D(
        instruction_memory_interface_data[21]), .Q(N227) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[21]  ( .G(N193), .D(n2476), .Q(
        N228) );
  DLH_X1 \instruction_FD_reg_reg[20]  ( .G(N193), .D(
        instruction_memory_interface_data[20]), .Q(N230) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[20]  ( .G(N193), .D(n2476), .Q(
        N231) );
  DLH_X1 \instruction_FD_reg_reg[19]  ( .G(N193), .D(
        instruction_memory_interface_data[19]), .Q(N233) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[19]  ( .G(N193), .D(n2476), .Q(
        N234) );
  DLH_X1 \instruction_FD_reg_reg[18]  ( .G(N193), .D(
        instruction_memory_interface_data[18]), .Q(N236) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[18]  ( .G(N193), .D(n2476), .Q(
        N237) );
  DLH_X1 \instruction_FD_reg_reg[17]  ( .G(N193), .D(
        instruction_memory_interface_data[17]), .Q(N239) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[17]  ( .G(N193), .D(n2476), .Q(
        N240) );
  DLH_X1 \instruction_FD_reg_reg[16]  ( .G(N193), .D(
        instruction_memory_interface_data[16]), .Q(N242) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[16]  ( .G(N193), .D(reset), .Q(
        N243) );
  DLH_X1 \instruction_FD_reg_reg[15]  ( .G(N193), .D(
        instruction_memory_interface_data[15]), .Q(N245) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[15]  ( .G(N193), .D(reset), .Q(
        N246) );
  DLH_X1 \instruction_FD_reg_reg[14]  ( .G(N193), .D(
        instruction_memory_interface_data[14]), .Q(N248) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[14]  ( .G(N193), .D(reset), .Q(
        N249) );
  DLH_X1 \instruction_FD_reg_reg[13]  ( .G(N193), .D(
        instruction_memory_interface_data[13]), .Q(N251) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[13]  ( .G(N193), .D(reset), .Q(
        N252) );
  DLH_X1 \instruction_FD_reg_reg[12]  ( .G(N193), .D(
        instruction_memory_interface_data[12]), .Q(N254) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[12]  ( .G(N193), .D(reset), .Q(
        N255) );
  DLH_X1 \instruction_FD_reg_reg[11]  ( .G(N193), .D(
        instruction_memory_interface_data[11]), .Q(N257) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[11]  ( .G(N193), .D(reset), .Q(
        N258) );
  DLH_X1 \instruction_FD_reg_reg[10]  ( .G(N193), .D(
        instruction_memory_interface_data[10]), .Q(N260) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[10]  ( .G(N193), .D(reset), .Q(
        N261) );
  DLH_X1 \instruction_FD_reg_reg[9]  ( .G(N193), .D(
        instruction_memory_interface_data[9]), .Q(N263) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[9]  ( .G(N193), .D(reset), .Q(N264) );
  DLH_X1 \instruction_FD_reg_reg[8]  ( .G(N193), .D(
        instruction_memory_interface_data[8]), .Q(N266) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[8]  ( .G(N193), .D(reset), .Q(N267) );
  DLH_X1 \instruction_FD_reg_reg[7]  ( .G(N193), .D(
        instruction_memory_interface_data[7]), .Q(N269) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[7]  ( .G(N193), .D(reset), .Q(N270) );
  DLH_X1 \instruction_FD_reg_reg[6]  ( .G(N193), .D(
        instruction_memory_interface_data[6]), .Q(N272) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[6]  ( .G(N193), .D(reset), .Q(N273) );
  DLH_X1 \instruction_FD_reg_reg[5]  ( .G(N193), .D(
        instruction_memory_interface_data[5]), .Q(N275) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[5]  ( .G(N193), .D(reset), .Q(N276) );
  DLH_X1 \instruction_FD_reg_reg[4]  ( .G(N193), .D(
        instruction_memory_interface_data[4]), .Q(N278) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[4]  ( .G(N193), .D(reset), .Q(N279) );
  DLH_X1 \instruction_FD_reg_reg[3]  ( .G(N193), .D(
        instruction_memory_interface_data[3]), .Q(N281) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[3]  ( .G(N193), .D(reset), .Q(N282) );
  DLH_X1 \instruction_FD_reg_reg[2]  ( .G(N193), .D(
        instruction_memory_interface_data[2]), .Q(N284) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[2]  ( .G(N193), .D(reset), .Q(N285) );
  DLH_X1 \instruction_FD_reg_reg[1]  ( .G(N193), .D(
        instruction_memory_interface_data[1]), .Q(N287) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[1]  ( .G(N193), .D(reset), .Q(N288) );
  DLH_X1 \instruction_FD_reg_reg[0]  ( .G(N193), .D(
        instruction_memory_interface_data[0]), .Q(N290) );
  DLH_X1 \instruction_FD_reg_tri_enable_reg[0]  ( .G(N193), .D(reset), .Q(N291) );
  DFF_X1 write_enable_csr_EX_reg_reg ( .D(n1761), .CK(clk), .Q(
        write_enable_csr_EX_reg), .QN() );
  DFF_X1 write_enable_EX_reg_reg ( .D(n1353), .CK(clk), .Q(), .QN(
        write_enable_EX_reg) );
  DFF_X1 write_enable_MW_reg_reg ( .D(N651), .CK(clk), .Q(write_enable_MW_reg), 
        .QN() );
  DFF_X1 \csr_index_EX_reg_reg[0]  ( .D(n1760), .CK(clk), .Q(
        csr_index_EX_reg[0]), .QN() );
  DFF_X1 \csr_index_EX_reg_reg[1]  ( .D(n1759), .CK(clk), .Q(
        csr_index_EX_reg[1]), .QN() );
  DFF_X1 \csr_index_EX_reg_reg[2]  ( .D(n1758), .CK(clk), .Q(
        csr_index_EX_reg[2]), .QN() );
  DFF_X1 \csr_index_EX_reg_reg[3]  ( .D(n1757), .CK(clk), .Q(
        csr_index_EX_reg[3]), .QN() );
  DFF_X1 \csr_index_EX_reg_reg[4]  ( .D(n1756), .CK(clk), .Q(
        csr_index_EX_reg[4]), .QN() );
  DFF_X1 \csr_index_EX_reg_reg[5]  ( .D(n1755), .CK(clk), .Q(
        csr_index_EX_reg[5]), .QN() );
  DFF_X1 \csr_index_EX_reg_reg[6]  ( .D(n1754), .CK(clk), .Q(
        csr_index_EX_reg[6]), .QN() );
  DFF_X1 \csr_index_EX_reg_reg[7]  ( .D(n1753), .CK(clk), .Q(
        csr_index_EX_reg[7]), .QN() );
  DFF_X1 \csr_index_EX_reg_reg[8]  ( .D(n1752), .CK(clk), .Q(
        csr_index_EX_reg[8]), .QN() );
  DFF_X1 \csr_index_EX_reg_reg[9]  ( .D(n1751), .CK(clk), .Q(
        csr_index_EX_reg[9]), .QN() );
  DFF_X1 \csr_index_EX_reg_reg[10]  ( .D(n1750), .CK(clk), .Q(
        csr_index_EX_reg[10]), .QN() );
  DFF_X1 \csr_index_EX_reg_reg[11]  ( .D(n1749), .CK(clk), .Q(
        csr_index_EX_reg[11]), .QN() );
  DFF_X1 \write_index_EX_reg_reg[0]  ( .D(n1156), .CK(clk), .Q(
        write_index_EX_reg[0]), .QN(n1173) );
  DFF_X1 \write_index_MW_reg_reg[0]  ( .D(N713), .CK(clk), .Q(
        write_index_MW_reg[0]), .QN() );
  DFF_X1 \write_index_EX_reg_reg[1]  ( .D(n1351), .CK(clk), .Q(), .QN(
        write_index_EX_reg[1]) );
  DFF_X1 \write_index_MW_reg_reg[1]  ( .D(N714), .CK(clk), .Q(
        write_index_MW_reg[1]), .QN() );
  DFF_X1 \write_index_EX_reg_reg[2]  ( .D(n1157), .CK(clk), .Q(
        write_index_EX_reg[2]), .QN(n1172) );
  DFF_X1 \write_index_MW_reg_reg[2]  ( .D(N715), .CK(clk), .Q(
        write_index_MW_reg[2]), .QN() );
  DFF_X1 \write_index_EX_reg_reg[3]  ( .D(n1158), .CK(clk), .Q(
        write_index_EX_reg[3]), .QN(n1171) );
  DFF_X1 \write_index_MW_reg_reg[3]  ( .D(N716), .CK(clk), .Q(
        write_index_MW_reg[3]), .QN() );
  DFF_X1 \write_index_EX_reg_reg[4]  ( .D(n1159), .CK(clk), .Q(
        write_index_EX_reg[4]), .QN(n1170) );
  DFF_X1 \write_index_MW_reg_reg[4]  ( .D(N717), .CK(clk), .Q(
        write_index_MW_reg[4]), .QN() );
  DFF_X1 \read_index_1_EX_reg_reg[0]  ( .D(n1748), .CK(clk), .Q(
        read_index_1_EX_reg[0]), .QN() );
  DFF_X1 \read_index_1_EX_reg_reg[1]  ( .D(n1747), .CK(clk), .Q(
        read_index_1_EX_reg[1]), .QN() );
  DFF_X1 \read_index_1_EX_reg_reg[2]  ( .D(n1746), .CK(clk), .Q(
        read_index_1_EX_reg[2]), .QN() );
  DFF_X1 \read_index_1_EX_reg_reg[3]  ( .D(n1745), .CK(clk), .Q(
        read_index_1_EX_reg[3]), .QN() );
  DFF_X1 \read_index_1_EX_reg_reg[4]  ( .D(n1744), .CK(clk), .Q(
        read_index_1_EX_reg[4]), .QN() );
  DFF_X1 \funct12_EX_reg_reg[0]  ( .D(n1347), .CK(clk), .Q(), .QN(
        funct12_EX_reg[0]) );
  DFF_X1 \funct12_MW_reg_reg[0]  ( .D(N669), .CK(clk), .Q(funct12_MW_reg[0]), 
        .QN() );
  DFF_X1 \funct12_EX_reg_reg[1]  ( .D(n1346), .CK(clk), .Q(), .QN(
        funct12_EX_reg[1]) );
  DFF_X1 \funct12_MW_reg_reg[1]  ( .D(N670), .CK(clk), .Q(funct12_MW_reg[1]), 
        .QN() );
  DFF_X1 \funct12_EX_reg_reg[2]  ( .D(n1345), .CK(clk), .Q(), .QN(
        funct12_EX_reg[2]) );
  DFF_X1 \funct12_MW_reg_reg[2]  ( .D(N671), .CK(clk), .Q(funct12_MW_reg[2]), 
        .QN() );
  DFF_X1 \funct12_EX_reg_reg[3]  ( .D(n1344), .CK(clk), .Q(), .QN(
        funct12_EX_reg[3]) );
  DFF_X1 \funct12_MW_reg_reg[3]  ( .D(N672), .CK(clk), .Q(funct12_MW_reg[3]), 
        .QN() );
  DFF_X1 \funct12_EX_reg_reg[4]  ( .D(n1343), .CK(clk), .Q(), .QN(
        funct12_EX_reg[4]) );
  DFF_X1 \funct12_MW_reg_reg[4]  ( .D(N673), .CK(clk), .Q(funct12_MW_reg[4]), 
        .QN() );
  DFF_X1 \funct12_EX_reg_reg[5]  ( .D(n1342), .CK(clk), .Q(), .QN(
        funct12_EX_reg[5]) );
  DFF_X1 \funct12_MW_reg_reg[5]  ( .D(N674), .CK(clk), .Q(funct12_MW_reg[5]), 
        .QN() );
  DFF_X1 \funct12_EX_reg_reg[6]  ( .D(n1341), .CK(clk), .Q(), .QN(
        funct12_EX_reg[6]) );
  DFF_X1 \funct12_MW_reg_reg[6]  ( .D(N675), .CK(clk), .Q(funct12_MW_reg[6]), 
        .QN() );
  DFF_X1 \funct12_EX_reg_reg[7]  ( .D(n1340), .CK(clk), .Q(), .QN(
        funct12_EX_reg[7]) );
  DFF_X1 \funct12_MW_reg_reg[7]  ( .D(N676), .CK(clk), .Q(funct12_MW_reg[7]), 
        .QN() );
  DFF_X1 \funct12_EX_reg_reg[8]  ( .D(n1339), .CK(clk), .Q(), .QN(
        funct12_EX_reg[8]) );
  DFF_X1 \funct12_MW_reg_reg[8]  ( .D(N677), .CK(clk), .Q(funct12_MW_reg[8]), 
        .QN() );
  DFF_X1 \funct12_EX_reg_reg[9]  ( .D(n1338), .CK(clk), .Q(), .QN(
        funct12_EX_reg[9]) );
  DFF_X1 \funct12_MW_reg_reg[9]  ( .D(N678), .CK(clk), .Q(funct12_MW_reg[9]), 
        .QN() );
  DFF_X1 \funct12_EX_reg_reg[10]  ( .D(n1337), .CK(clk), .Q(), .QN(
        funct12_EX_reg[10]) );
  DFF_X1 \funct12_MW_reg_reg[10]  ( .D(N679), .CK(clk), .Q(funct12_MW_reg[10]), 
        .QN() );
  DFF_X1 \funct12_EX_reg_reg[11]  ( .D(n1336), .CK(clk), .Q(), .QN(
        funct12_EX_reg[11]) );
  DFF_X1 \funct12_MW_reg_reg[11]  ( .D(N680), .CK(clk), .Q(funct12_MW_reg[11]), 
        .QN() );
  DFF_X1 \funct7_EX_reg_reg[0]  ( .D(n1335), .CK(clk), .Q(), .QN(
        funct7_EX_reg[0]) );
  DFF_X1 \funct7_MW_reg_reg[0]  ( .D(N662), .CK(clk), .Q(funct7_MW_reg[0]), 
        .QN() );
  DFF_X1 \funct7_EX_reg_reg[1]  ( .D(n1334), .CK(clk), .Q(), .QN(
        funct7_EX_reg[1]) );
  DFF_X1 \funct7_MW_reg_reg[1]  ( .D(N663), .CK(clk), .Q(funct7_MW_reg[1]), 
        .QN() );
  DFF_X1 \funct7_EX_reg_reg[2]  ( .D(n1333), .CK(clk), .Q(), .QN(
        funct7_EX_reg[2]) );
  DFF_X1 \funct7_MW_reg_reg[2]  ( .D(N664), .CK(clk), .Q(funct7_MW_reg[2]), 
        .QN() );
  DFF_X1 \funct7_EX_reg_reg[3]  ( .D(n1332), .CK(clk), .Q(), .QN(
        funct7_EX_reg[3]) );
  DFF_X1 \funct7_MW_reg_reg[3]  ( .D(N665), .CK(clk), .Q(funct7_MW_reg[3]), 
        .QN() );
  DFF_X1 \funct7_EX_reg_reg[4]  ( .D(n1331), .CK(clk), .Q(), .QN(
        funct7_EX_reg[4]) );
  DFF_X1 \funct7_MW_reg_reg[4]  ( .D(N666), .CK(clk), .Q(funct7_MW_reg[4]), 
        .QN() );
  DFF_X1 \funct7_EX_reg_reg[5]  ( .D(n1330), .CK(clk), .Q(), .QN(
        funct7_EX_reg[5]) );
  DFF_X1 \funct7_MW_reg_reg[5]  ( .D(N667), .CK(clk), .Q(funct7_MW_reg[5]), 
        .QN() );
  DFF_X1 \funct7_EX_reg_reg[6]  ( .D(n1329), .CK(clk), .Q(), .QN(
        funct7_EX_reg[6]) );
  DFF_X1 \funct7_MW_reg_reg[6]  ( .D(N668), .CK(clk), .Q(funct7_MW_reg[6]), 
        .QN() );
  DFF_X1 \funct3_EX_reg_reg[0]  ( .D(n1328), .CK(clk), .Q(), .QN(
        funct3_EX_reg[0]) );
  DFF_X1 \funct3_MW_reg_reg[0]  ( .D(N659), .CK(clk), .Q(funct3_MW_reg[0]), 
        .QN() );
  DFF_X1 \funct3_EX_reg_reg[1]  ( .D(n1327), .CK(clk), .Q(), .QN(
        funct3_EX_reg[1]) );
  DFF_X1 \funct3_MW_reg_reg[1]  ( .D(N660), .CK(clk), .Q(funct3_MW_reg[1]), 
        .QN() );
  DFF_X1 \funct3_EX_reg_reg[2]  ( .D(n1160), .CK(clk), .Q(funct3_EX_reg[2]), 
        .QN(n1169) );
  DFF_X1 \funct3_MW_reg_reg[2]  ( .D(N661), .CK(clk), .Q(funct3_MW_reg[2]), 
        .QN() );
  DFF_X1 \opcode_MW_reg_reg[2]  ( .D(N654), .CK(clk), .Q(opcode_MW_reg[2]), 
        .QN(n1210) );
  DFF_X1 \opcode_MW_reg_reg[3]  ( .D(N655), .CK(clk), .Q(opcode_MW_reg[3]), 
        .QN(n789) );
  DFF_X1 \opcode_MW_reg_reg[5]  ( .D(N657), .CK(clk), .Q(opcode_MW_reg[5]), 
        .QN(n1208) );
  DFF_X1 \opcode_MW_reg_reg[6]  ( .D(N658), .CK(clk), .Q(opcode_MW_reg[6]), 
        .QN(n790) );
  DFF_X1 \instruction_type_EX_reg_reg[0]  ( .D(n1708), .CK(clk), .Q(
        instruction_type_EX_reg[0]), .QN() );
  DFF_X1 \instruction_type_EX_reg_reg[1]  ( .D(n1284), .CK(clk), .Q(), .QN(
        instruction_type_EX_reg[1]) );
  DFF_X1 \immediate_EX_reg_reg[0]  ( .D(n1318), .CK(clk), .Q(), .QN(
        immediate_EX_reg[0]) );
  DFF_X1 \immediate_MW_reg_reg[0]  ( .D(N681), .CK(clk), .Q(
        immediate_MW_reg[0]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[1]  ( .D(n1317), .CK(clk), .Q(), .QN(
        immediate_EX_reg[1]) );
  DFF_X1 \immediate_MW_reg_reg[1]  ( .D(N682), .CK(clk), .Q(
        immediate_MW_reg[1]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[2]  ( .D(n1316), .CK(clk), .Q(), .QN(
        immediate_EX_reg[2]) );
  DFF_X1 \immediate_MW_reg_reg[2]  ( .D(N683), .CK(clk), .Q(
        immediate_MW_reg[2]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[3]  ( .D(n1315), .CK(clk), .Q(), .QN(
        immediate_EX_reg[3]) );
  DFF_X1 \immediate_MW_reg_reg[3]  ( .D(N684), .CK(clk), .Q(
        immediate_MW_reg[3]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[4]  ( .D(n1314), .CK(clk), .Q(), .QN(
        immediate_EX_reg[4]) );
  DFF_X1 \immediate_MW_reg_reg[4]  ( .D(N685), .CK(clk), .Q(
        immediate_MW_reg[4]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[5]  ( .D(n1313), .CK(clk), .Q(), .QN(
        immediate_EX_reg[5]) );
  DFF_X1 \immediate_MW_reg_reg[5]  ( .D(N686), .CK(clk), .Q(
        immediate_MW_reg[5]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[6]  ( .D(n1312), .CK(clk), .Q(n2168), .QN(
        immediate_EX_reg[6]) );
  DFF_X1 \immediate_MW_reg_reg[6]  ( .D(N687), .CK(clk), .Q(
        immediate_MW_reg[6]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[7]  ( .D(n1311), .CK(clk), .Q(n2169), .QN(
        immediate_EX_reg[7]) );
  DFF_X1 \immediate_MW_reg_reg[7]  ( .D(N688), .CK(clk), .Q(
        immediate_MW_reg[7]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[8]  ( .D(n1310), .CK(clk), .Q(n2170), .QN(
        immediate_EX_reg[8]) );
  DFF_X1 \immediate_MW_reg_reg[8]  ( .D(N689), .CK(clk), .Q(
        immediate_MW_reg[8]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[9]  ( .D(n1309), .CK(clk), .Q(n2175), .QN(
        immediate_EX_reg[9]) );
  DFF_X1 \immediate_MW_reg_reg[9]  ( .D(N690), .CK(clk), .Q(
        immediate_MW_reg[9]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[10]  ( .D(n1308), .CK(clk), .Q(n2171), .QN(
        immediate_EX_reg[10]) );
  DFF_X1 \immediate_MW_reg_reg[10]  ( .D(N691), .CK(clk), .Q(
        immediate_MW_reg[10]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[11]  ( .D(n1307), .CK(clk), .Q(n2172), .QN(
        immediate_EX_reg[11]) );
  DFF_X1 \immediate_MW_reg_reg[11]  ( .D(N692), .CK(clk), .Q(
        immediate_MW_reg[11]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[12]  ( .D(n1306), .CK(clk), .Q(n2173), .QN(
        immediate_EX_reg[12]) );
  DFF_X1 \immediate_MW_reg_reg[12]  ( .D(N693), .CK(clk), .Q(
        immediate_MW_reg[12]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[13]  ( .D(n1305), .CK(clk), .Q(n2176), .QN(
        immediate_EX_reg[13]) );
  DFF_X1 \immediate_MW_reg_reg[13]  ( .D(N694), .CK(clk), .Q(
        immediate_MW_reg[13]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[14]  ( .D(n1304), .CK(clk), .Q(n2177), .QN(
        immediate_EX_reg[14]) );
  DFF_X1 \immediate_MW_reg_reg[14]  ( .D(N695), .CK(clk), .Q(
        immediate_MW_reg[14]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[15]  ( .D(n1303), .CK(clk), .Q(n2178), .QN(
        immediate_EX_reg[15]) );
  DFF_X1 \immediate_MW_reg_reg[15]  ( .D(N696), .CK(clk), .Q(
        immediate_MW_reg[15]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[16]  ( .D(n1302), .CK(clk), .Q(n2174), .QN(
        immediate_EX_reg[16]) );
  DFF_X1 \immediate_MW_reg_reg[16]  ( .D(N697), .CK(clk), .Q(
        immediate_MW_reg[16]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[17]  ( .D(n1301), .CK(clk), .Q(n2179), .QN(
        immediate_EX_reg[17]) );
  DFF_X1 \immediate_MW_reg_reg[17]  ( .D(N698), .CK(clk), .Q(
        immediate_MW_reg[17]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[18]  ( .D(n1300), .CK(clk), .Q(n2160), .QN(
        immediate_EX_reg[18]) );
  DFF_X1 \immediate_MW_reg_reg[18]  ( .D(N699), .CK(clk), .Q(
        immediate_MW_reg[18]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[19]  ( .D(n1299), .CK(clk), .Q(n2157), .QN(
        immediate_EX_reg[19]) );
  DFF_X1 \immediate_MW_reg_reg[19]  ( .D(N700), .CK(clk), .Q(
        immediate_MW_reg[19]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[20]  ( .D(n1298), .CK(clk), .Q(n2167), .QN(
        immediate_EX_reg[20]) );
  DFF_X1 \immediate_MW_reg_reg[20]  ( .D(N701), .CK(clk), .Q(
        immediate_MW_reg[20]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[21]  ( .D(n1297), .CK(clk), .Q(n2162), .QN(
        immediate_EX_reg[21]) );
  DFF_X1 \immediate_MW_reg_reg[21]  ( .D(N702), .CK(clk), .Q(
        immediate_MW_reg[21]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[22]  ( .D(n1296), .CK(clk), .Q(n2166), .QN(
        immediate_EX_reg[22]) );
  DFF_X1 \immediate_MW_reg_reg[22]  ( .D(N703), .CK(clk), .Q(
        immediate_MW_reg[22]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[23]  ( .D(n1295), .CK(clk), .Q(), .QN(
        immediate_EX_reg[23]) );
  DFF_X1 \immediate_MW_reg_reg[23]  ( .D(N704), .CK(clk), .Q(
        immediate_MW_reg[23]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[24]  ( .D(n1294), .CK(clk), .Q(n2158), .QN(
        immediate_EX_reg[24]) );
  DFF_X1 \immediate_MW_reg_reg[24]  ( .D(N705), .CK(clk), .Q(
        immediate_MW_reg[24]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[25]  ( .D(n1293), .CK(clk), .Q(n2159), .QN(
        immediate_EX_reg[25]) );
  DFF_X1 \immediate_MW_reg_reg[25]  ( .D(N706), .CK(clk), .Q(
        immediate_MW_reg[25]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[26]  ( .D(n1292), .CK(clk), .Q(n2163), .QN(
        immediate_EX_reg[26]) );
  DFF_X1 \immediate_MW_reg_reg[26]  ( .D(N707), .CK(clk), .Q(
        immediate_MW_reg[26]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[27]  ( .D(n1291), .CK(clk), .Q(n2164), .QN(
        immediate_EX_reg[27]) );
  DFF_X1 \immediate_MW_reg_reg[27]  ( .D(N708), .CK(clk), .Q(
        immediate_MW_reg[27]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[28]  ( .D(n1290), .CK(clk), .Q(), .QN(
        immediate_EX_reg[28]) );
  DFF_X1 \immediate_MW_reg_reg[28]  ( .D(N709), .CK(clk), .Q(
        immediate_MW_reg[28]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[29]  ( .D(n1289), .CK(clk), .Q(n2165), .QN(
        immediate_EX_reg[29]) );
  DFF_X1 \immediate_MW_reg_reg[29]  ( .D(N710), .CK(clk), .Q(
        immediate_MW_reg[29]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[30]  ( .D(n1288), .CK(clk), .Q(n2161), .QN(
        immediate_EX_reg[30]) );
  DFF_X1 \immediate_MW_reg_reg[30]  ( .D(N711), .CK(clk), .Q(
        immediate_MW_reg[30]), .QN() );
  DFF_X1 \immediate_EX_reg_reg[31]  ( .D(n1287), .CK(clk), .Q(), .QN(
        immediate_EX_reg[31]) );
  DFF_X1 \immediate_MW_reg_reg[31]  ( .D(N712), .CK(clk), .Q(
        immediate_MW_reg[31]), .QN() );
  DFF_X1 \instruction_type_EX_reg_reg[2]  ( .D(n1282), .CK(clk), .Q(), .QN(
        instruction_type_EX_reg[2]) );
  DFF_X1 \opcode_MW_reg_reg[4]  ( .D(N656), .CK(clk), .Q(opcode_MW_reg[4]), 
        .QN(n1209) );
  DFF_X1 \csr_data_EX_reg_reg[0]  ( .D(n1740), .CK(clk), .Q(csr_data_EX_reg[0]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[1]  ( .D(n1739), .CK(clk), .Q(csr_data_EX_reg[1]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[2]  ( .D(n1738), .CK(clk), .Q(csr_data_EX_reg[2]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[3]  ( .D(n1737), .CK(clk), .Q(csr_data_EX_reg[3]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[4]  ( .D(n1736), .CK(clk), .Q(csr_data_EX_reg[4]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[5]  ( .D(n1735), .CK(clk), .Q(csr_data_EX_reg[5]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[6]  ( .D(n1734), .CK(clk), .Q(csr_data_EX_reg[6]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[7]  ( .D(n1733), .CK(clk), .Q(csr_data_EX_reg[7]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[8]  ( .D(n1732), .CK(clk), .Q(csr_data_EX_reg[8]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[9]  ( .D(n1731), .CK(clk), .Q(csr_data_EX_reg[9]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[10]  ( .D(n1730), .CK(clk), .Q(
        csr_data_EX_reg[10]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[11]  ( .D(n1729), .CK(clk), .Q(
        csr_data_EX_reg[11]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[12]  ( .D(n1728), .CK(clk), .Q(
        csr_data_EX_reg[12]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[13]  ( .D(n1727), .CK(clk), .Q(
        csr_data_EX_reg[13]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[14]  ( .D(n1726), .CK(clk), .Q(
        csr_data_EX_reg[14]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[15]  ( .D(n1725), .CK(clk), .Q(
        csr_data_EX_reg[15]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[16]  ( .D(n1724), .CK(clk), .Q(
        csr_data_EX_reg[16]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[17]  ( .D(n1723), .CK(clk), .Q(
        csr_data_EX_reg[17]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[18]  ( .D(n1722), .CK(clk), .Q(
        csr_data_EX_reg[18]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[19]  ( .D(n1721), .CK(clk), .Q(
        csr_data_EX_reg[19]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[20]  ( .D(n1720), .CK(clk), .Q(
        csr_data_EX_reg[20]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[21]  ( .D(n1719), .CK(clk), .Q(
        csr_data_EX_reg[21]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[22]  ( .D(n1718), .CK(clk), .Q(
        csr_data_EX_reg[22]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[23]  ( .D(n1717), .CK(clk), .Q(
        csr_data_EX_reg[23]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[24]  ( .D(n1716), .CK(clk), .Q(
        csr_data_EX_reg[24]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[25]  ( .D(n1715), .CK(clk), .Q(
        csr_data_EX_reg[25]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[26]  ( .D(n1714), .CK(clk), .Q(
        csr_data_EX_reg[26]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[27]  ( .D(n1713), .CK(clk), .Q(
        csr_data_EX_reg[27]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[28]  ( .D(n1712), .CK(clk), .Q(
        csr_data_EX_reg[28]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[29]  ( .D(n1711), .CK(clk), .Q(
        csr_data_EX_reg[29]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[30]  ( .D(n1710), .CK(clk), .Q(
        csr_data_EX_reg[30]), .QN() );
  DFF_X1 \csr_data_EX_reg_reg[31]  ( .D(n1709), .CK(clk), .Q(
        csr_data_EX_reg[31]), .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[0]  ( .D(n950), .CK(clk), .Q(csr_rd_MW_reg[0]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[1]  ( .D(n949), .CK(clk), .Q(csr_rd_MW_reg[1]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[2]  ( .D(n948), .CK(clk), .Q(csr_rd_MW_reg[2]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[3]  ( .D(n947), .CK(clk), .Q(csr_rd_MW_reg[3]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[4]  ( .D(n946), .CK(clk), .Q(csr_rd_MW_reg[4]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[5]  ( .D(n945), .CK(clk), .Q(csr_rd_MW_reg[5]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[6]  ( .D(n944), .CK(clk), .Q(csr_rd_MW_reg[6]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[7]  ( .D(n943), .CK(clk), .Q(csr_rd_MW_reg[7]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[8]  ( .D(n942), .CK(clk), .Q(csr_rd_MW_reg[8]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[9]  ( .D(n941), .CK(clk), .Q(csr_rd_MW_reg[9]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[10]  ( .D(n940), .CK(clk), .Q(csr_rd_MW_reg[10]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[11]  ( .D(n939), .CK(clk), .Q(csr_rd_MW_reg[11]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[12]  ( .D(n938), .CK(clk), .Q(csr_rd_MW_reg[12]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[13]  ( .D(n937), .CK(clk), .Q(csr_rd_MW_reg[13]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[14]  ( .D(n936), .CK(clk), .Q(csr_rd_MW_reg[14]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[15]  ( .D(n935), .CK(clk), .Q(csr_rd_MW_reg[15]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[16]  ( .D(n934), .CK(clk), .Q(csr_rd_MW_reg[16]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[17]  ( .D(n933), .CK(clk), .Q(csr_rd_MW_reg[17]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[18]  ( .D(n932), .CK(clk), .Q(csr_rd_MW_reg[18]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[19]  ( .D(n931), .CK(clk), .Q(csr_rd_MW_reg[19]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[20]  ( .D(n930), .CK(clk), .Q(csr_rd_MW_reg[20]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[21]  ( .D(n929), .CK(clk), .Q(csr_rd_MW_reg[21]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[22]  ( .D(n928), .CK(clk), .Q(csr_rd_MW_reg[22]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[23]  ( .D(n927), .CK(clk), .Q(csr_rd_MW_reg[23]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[24]  ( .D(n926), .CK(clk), .Q(csr_rd_MW_reg[24]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[25]  ( .D(n925), .CK(clk), .Q(csr_rd_MW_reg[25]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[26]  ( .D(n924), .CK(clk), .Q(csr_rd_MW_reg[26]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[27]  ( .D(n923), .CK(clk), .Q(csr_rd_MW_reg[27]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[28]  ( .D(n922), .CK(clk), .Q(csr_rd_MW_reg[28]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[29]  ( .D(n921), .CK(clk), .Q(csr_rd_MW_reg[29]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[30]  ( .D(n920), .CK(clk), .Q(csr_rd_MW_reg[30]), 
        .QN() );
  DFF_X1 \csr_rd_MW_reg_reg[31]  ( .D(n919), .CK(clk), .Q(csr_rd_MW_reg[31]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[0]  ( .D(n918), .CK(clk), .Q(address_MW_reg[0]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[1]  ( .D(n917), .CK(clk), .Q(address_MW_reg[1]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[2]  ( .D(n916), .CK(clk), .Q(address_MW_reg[2]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[3]  ( .D(n915), .CK(clk), .Q(address_MW_reg[3]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[4]  ( .D(n914), .CK(clk), .Q(address_MW_reg[4]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[5]  ( .D(n913), .CK(clk), .Q(address_MW_reg[5]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[6]  ( .D(n912), .CK(clk), .Q(address_MW_reg[6]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[7]  ( .D(n911), .CK(clk), .Q(address_MW_reg[7]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[8]  ( .D(n910), .CK(clk), .Q(address_MW_reg[8]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[9]  ( .D(n909), .CK(clk), .Q(address_MW_reg[9]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[10]  ( .D(n908), .CK(clk), .Q(address_MW_reg[10]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[11]  ( .D(n907), .CK(clk), .Q(address_MW_reg[11]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[12]  ( .D(n906), .CK(clk), .Q(address_MW_reg[12]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[13]  ( .D(n905), .CK(clk), .Q(address_MW_reg[13]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[14]  ( .D(n904), .CK(clk), .Q(address_MW_reg[14]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[15]  ( .D(n903), .CK(clk), .Q(address_MW_reg[15]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[16]  ( .D(n902), .CK(clk), .Q(address_MW_reg[16]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[17]  ( .D(n901), .CK(clk), .Q(address_MW_reg[17]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[18]  ( .D(n900), .CK(clk), .Q(address_MW_reg[18]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[19]  ( .D(n899), .CK(clk), .Q(address_MW_reg[19]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[20]  ( .D(n898), .CK(clk), .Q(address_MW_reg[20]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[21]  ( .D(n897), .CK(clk), .Q(address_MW_reg[21]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[22]  ( .D(n896), .CK(clk), .Q(address_MW_reg[22]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[23]  ( .D(n895), .CK(clk), .Q(address_MW_reg[23]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[24]  ( .D(n894), .CK(clk), .Q(address_MW_reg[24]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[25]  ( .D(n893), .CK(clk), .Q(address_MW_reg[25]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[26]  ( .D(n892), .CK(clk), .Q(address_MW_reg[26]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[27]  ( .D(n891), .CK(clk), .Q(address_MW_reg[27]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[28]  ( .D(n890), .CK(clk), .Q(address_MW_reg[28]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[29]  ( .D(n889), .CK(clk), .Q(address_MW_reg[29]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[30]  ( .D(n888), .CK(clk), .Q(address_MW_reg[30]), 
        .QN() );
  DFF_X1 \address_MW_reg_reg[31]  ( .D(n887), .CK(clk), .Q(address_MW_reg[31]), 
        .QN() );
  DFF_X1 \pc_FD_reg_reg[31]  ( .D(n1613), .CK(clk), .Q(pc_FD_reg[31]), .QN()
         );
  DFF_X1 \next_pc_EX_reg_reg[0]  ( .D(n1707), .CK(clk), .Q(next_pc_EX_reg[0]), 
        .QN(n244) );
  DFF_X1 \next_pc_MW_reg_reg[0]  ( .D(n885), .CK(clk), .Q(n2180), .QN(n243) );
  DFF_X1 \pc_FD_reg_reg[0]  ( .D(n1675), .CK(clk), .Q(pc_FD_reg[0]), .QN() );
  DFF_X1 \pc_EX_reg_reg[0]  ( .D(n1674), .CK(clk), .Q(pc_EX_reg[0]), .QN() );
  DFF_X1 \next_pc_EX_reg_reg[1]  ( .D(n1706), .CK(clk), .Q(next_pc_EX_reg[1]), 
        .QN(n246) );
  DFF_X1 \next_pc_MW_reg_reg[1]  ( .D(n882), .CK(clk), .Q(n2181), .QN(n245) );
  DFF_X1 \pc_FD_reg_reg[1]  ( .D(n1673), .CK(clk), .Q(pc_FD_reg[1]), .QN() );
  DFF_X1 \pc_EX_reg_reg[1]  ( .D(n1672), .CK(clk), .Q(pc_EX_reg[1]), .QN() );
  DFF_X1 \next_pc_EX_reg_reg[2]  ( .D(n1705), .CK(clk), .Q(next_pc_EX_reg[2]), 
        .QN(n248) );
  DFF_X1 \next_pc_MW_reg_reg[2]  ( .D(n879), .CK(clk), .Q(n2182), .QN(n247) );
  DFF_X1 \pc_FD_reg_reg[2]  ( .D(n1671), .CK(clk), .Q(pc_FD_reg[2]), .QN() );
  DFF_X1 \pc_EX_reg_reg[2]  ( .D(n1670), .CK(clk), .Q(pc_EX_reg[2]), .QN() );
  DFF_X1 \next_pc_EX_reg_reg[3]  ( .D(n1704), .CK(clk), .Q(next_pc_EX_reg[3]), 
        .QN(n250) );
  DFF_X1 \next_pc_MW_reg_reg[3]  ( .D(n876), .CK(clk), .Q(n2183), .QN(n249) );
  DFF_X1 \pc_FD_reg_reg[3]  ( .D(n1669), .CK(clk), .Q(pc_FD_reg[3]), .QN() );
  DFF_X1 \pc_EX_reg_reg[3]  ( .D(n1668), .CK(clk), .Q(pc_EX_reg[3]), .QN() );
  DFF_X1 \next_pc_EX_reg_reg[4]  ( .D(n1703), .CK(clk), .Q(next_pc_EX_reg[4]), 
        .QN(n252) );
  DFF_X1 \next_pc_MW_reg_reg[4]  ( .D(n873), .CK(clk), .Q(n2184), .QN(n251) );
  DFF_X1 \pc_FD_reg_reg[4]  ( .D(n1667), .CK(clk), .Q(pc_FD_reg[4]), .QN() );
  DFF_X1 \pc_EX_reg_reg[4]  ( .D(n1666), .CK(clk), .Q(pc_EX_reg[4]), .QN() );
  DFF_X1 \next_pc_EX_reg_reg[5]  ( .D(n1702), .CK(clk), .Q(next_pc_EX_reg[5]), 
        .QN(n254) );
  DFF_X1 \next_pc_MW_reg_reg[5]  ( .D(n870), .CK(clk), .Q(n2185), .QN(n253) );
  DFF_X1 \pc_FD_reg_reg[5]  ( .D(n1665), .CK(clk), .Q(pc_FD_reg[5]), .QN() );
  DFF_X1 \pc_EX_reg_reg[5]  ( .D(n1664), .CK(clk), .Q(pc_EX_reg[5]), .QN() );
  DFF_X1 \next_pc_EX_reg_reg[6]  ( .D(n1701), .CK(clk), .Q(next_pc_EX_reg[6]), 
        .QN(n256) );
  DFF_X1 \next_pc_MW_reg_reg[6]  ( .D(n867), .CK(clk), .Q(n2186), .QN(n255) );
  DFF_X1 \pc_FD_reg_reg[6]  ( .D(n1663), .CK(clk), .Q(pc_FD_reg[6]), .QN() );
  DFF_X1 \pc_EX_reg_reg[6]  ( .D(n1662), .CK(clk), .Q(pc_EX_reg[6]), .QN() );
  DFF_X1 \next_pc_EX_reg_reg[7]  ( .D(n1700), .CK(clk), .Q(next_pc_EX_reg[7]), 
        .QN(n258) );
  DFF_X1 \next_pc_MW_reg_reg[7]  ( .D(n864), .CK(clk), .Q(n2187), .QN(n257) );
  DFF_X1 \pc_FD_reg_reg[7]  ( .D(n1661), .CK(clk), .Q(pc_FD_reg[7]), .QN() );
  DFF_X1 \pc_EX_reg_reg[7]  ( .D(n1660), .CK(clk), .Q(pc_EX_reg[7]), .QN() );
  DFF_X1 \next_pc_EX_reg_reg[8]  ( .D(n1699), .CK(clk), .Q(next_pc_EX_reg[8]), 
        .QN(n260) );
  DFF_X1 \next_pc_MW_reg_reg[8]  ( .D(n861), .CK(clk), .Q(n2188), .QN(n259) );
  DFF_X1 \pc_FD_reg_reg[8]  ( .D(n1659), .CK(clk), .Q(pc_FD_reg[8]), .QN() );
  DFF_X1 \pc_EX_reg_reg[8]  ( .D(n1658), .CK(clk), .Q(pc_EX_reg[8]), .QN() );
  DFF_X1 \next_pc_EX_reg_reg[9]  ( .D(n1698), .CK(clk), .Q(next_pc_EX_reg[9]), 
        .QN(n262) );
  DFF_X1 \next_pc_MW_reg_reg[9]  ( .D(n858), .CK(clk), .Q(n2189), .QN(n261) );
  DFF_X1 \pc_FD_reg_reg[9]  ( .D(n1657), .CK(clk), .Q(pc_FD_reg[9]), .QN() );
  DFF_X1 \pc_EX_reg_reg[9]  ( .D(n1656), .CK(clk), .Q(pc_EX_reg[9]), .QN() );
  DFF_X1 \next_pc_EX_reg_reg[10]  ( .D(n1697), .CK(clk), .Q(next_pc_EX_reg[10]), .QN(n264) );
  DFF_X1 \next_pc_MW_reg_reg[10]  ( .D(n855), .CK(clk), .Q(n2190), .QN(n263)
         );
  DFF_X1 \pc_FD_reg_reg[10]  ( .D(n1655), .CK(clk), .Q(pc_FD_reg[10]), .QN()
         );
  DFF_X1 \pc_EX_reg_reg[10]  ( .D(n1654), .CK(clk), .Q(pc_EX_reg[10]), .QN()
         );
  DFF_X1 \next_pc_EX_reg_reg[11]  ( .D(n1696), .CK(clk), .Q(next_pc_EX_reg[11]), .QN(n266) );
  DFF_X1 \next_pc_MW_reg_reg[11]  ( .D(n852), .CK(clk), .Q(n2191), .QN(n265)
         );
  DFF_X1 \pc_FD_reg_reg[11]  ( .D(n1653), .CK(clk), .Q(pc_FD_reg[11]), .QN()
         );
  DFF_X1 \pc_EX_reg_reg[11]  ( .D(n1652), .CK(clk), .Q(pc_EX_reg[11]), .QN()
         );
  DFF_X1 \next_pc_EX_reg_reg[12]  ( .D(n1695), .CK(clk), .Q(next_pc_EX_reg[12]), .QN(n268) );
  DFF_X1 \next_pc_MW_reg_reg[12]  ( .D(n849), .CK(clk), .Q(n2192), .QN(n267)
         );
  DFF_X1 \pc_FD_reg_reg[12]  ( .D(n1651), .CK(clk), .Q(pc_FD_reg[12]), .QN()
         );
  DFF_X1 \pc_EX_reg_reg[12]  ( .D(n1650), .CK(clk), .Q(pc_EX_reg[12]), .QN()
         );
  DFF_X1 \next_pc_EX_reg_reg[13]  ( .D(n1694), .CK(clk), .Q(next_pc_EX_reg[13]), .QN(n270) );
  DFF_X1 \next_pc_MW_reg_reg[13]  ( .D(n846), .CK(clk), .Q(n2193), .QN(n269)
         );
  DFF_X1 \pc_FD_reg_reg[13]  ( .D(n1649), .CK(clk), .Q(pc_FD_reg[13]), .QN()
         );
  DFF_X1 \pc_EX_reg_reg[13]  ( .D(n1648), .CK(clk), .Q(pc_EX_reg[13]), .QN()
         );
  DFF_X1 \next_pc_EX_reg_reg[14]  ( .D(n1693), .CK(clk), .Q(next_pc_EX_reg[14]), .QN(n272) );
  DFF_X1 \next_pc_MW_reg_reg[14]  ( .D(n843), .CK(clk), .Q(n2194), .QN(n271)
         );
  DFF_X1 \pc_FD_reg_reg[14]  ( .D(n1647), .CK(clk), .Q(pc_FD_reg[14]), .QN()
         );
  DFF_X1 \pc_EX_reg_reg[14]  ( .D(n1646), .CK(clk), .Q(pc_EX_reg[14]), .QN()
         );
  DFF_X1 \next_pc_EX_reg_reg[15]  ( .D(n1692), .CK(clk), .Q(next_pc_EX_reg[15]), .QN(n274) );
  DFF_X1 \next_pc_MW_reg_reg[15]  ( .D(n840), .CK(clk), .Q(n2195), .QN(n273)
         );
  DFF_X1 \pc_FD_reg_reg[15]  ( .D(n1645), .CK(clk), .Q(pc_FD_reg[15]), .QN()
         );
  DFF_X1 \pc_EX_reg_reg[15]  ( .D(n1644), .CK(clk), .Q(pc_EX_reg[15]), .QN()
         );
  DFF_X1 \next_pc_EX_reg_reg[16]  ( .D(n1691), .CK(clk), .Q(next_pc_EX_reg[16]), .QN(n276) );
  DFF_X1 \next_pc_MW_reg_reg[16]  ( .D(n837), .CK(clk), .Q(n2196), .QN(n275)
         );
  DFF_X1 \pc_FD_reg_reg[16]  ( .D(n1643), .CK(clk), .Q(pc_FD_reg[16]), .QN()
         );
  DFF_X1 \pc_EX_reg_reg[16]  ( .D(n1642), .CK(clk), .Q(pc_EX_reg[16]), .QN()
         );
  DFF_X1 \next_pc_EX_reg_reg[17]  ( .D(n1690), .CK(clk), .Q(next_pc_EX_reg[17]), .QN(n278) );
  DFF_X1 \next_pc_MW_reg_reg[17]  ( .D(n834), .CK(clk), .Q(n2197), .QN(n277)
         );
  DFF_X1 \pc_FD_reg_reg[17]  ( .D(n1641), .CK(clk), .Q(pc_FD_reg[17]), .QN()
         );
  DFF_X1 \pc_EX_reg_reg[17]  ( .D(n1640), .CK(clk), .Q(pc_EX_reg[17]), .QN()
         );
  DFF_X1 \next_pc_EX_reg_reg[18]  ( .D(n1689), .CK(clk), .Q(next_pc_EX_reg[18]), .QN(n280) );
  DFF_X1 \next_pc_MW_reg_reg[18]  ( .D(n831), .CK(clk), .Q(n2198), .QN(n279)
         );
  DFF_X1 \pc_FD_reg_reg[18]  ( .D(n1639), .CK(clk), .Q(pc_FD_reg[18]), .QN()
         );
  DFF_X1 \pc_EX_reg_reg[18]  ( .D(n1638), .CK(clk), .Q(pc_EX_reg[18]), .QN()
         );
  DFF_X1 \next_pc_EX_reg_reg[19]  ( .D(n1688), .CK(clk), .Q(next_pc_EX_reg[19]), .QN(n282) );
  DFF_X1 \next_pc_MW_reg_reg[19]  ( .D(n828), .CK(clk), .Q(n2199), .QN(n281)
         );
  DFF_X1 \pc_FD_reg_reg[19]  ( .D(n1637), .CK(clk), .Q(pc_FD_reg[19]), .QN()
         );
  DFF_X1 \pc_EX_reg_reg[19]  ( .D(n1636), .CK(clk), .Q(pc_EX_reg[19]), .QN()
         );
  DFF_X1 \next_pc_EX_reg_reg[20]  ( .D(n1687), .CK(clk), .Q(next_pc_EX_reg[20]), .QN(n284) );
  DFF_X1 \next_pc_MW_reg_reg[20]  ( .D(n825), .CK(clk), .Q(n2200), .QN(n283)
         );
  DFF_X1 \pc_FD_reg_reg[20]  ( .D(n1635), .CK(clk), .Q(pc_FD_reg[20]), .QN()
         );
  DFF_X1 \pc_EX_reg_reg[20]  ( .D(n1634), .CK(clk), .Q(pc_EX_reg[20]), .QN()
         );
  DFF_X1 \next_pc_EX_reg_reg[21]  ( .D(n1686), .CK(clk), .Q(next_pc_EX_reg[21]), .QN(n286) );
  DFF_X1 \next_pc_MW_reg_reg[21]  ( .D(n822), .CK(clk), .Q(n2201), .QN(n285)
         );
  DFF_X1 \pc_FD_reg_reg[21]  ( .D(n1633), .CK(clk), .Q(pc_FD_reg[21]), .QN()
         );
  DFF_X1 \pc_EX_reg_reg[21]  ( .D(n1632), .CK(clk), .Q(pc_EX_reg[21]), .QN()
         );
  DFF_X1 \next_pc_EX_reg_reg[22]  ( .D(n1685), .CK(clk), .Q(next_pc_EX_reg[22]), .QN(n288) );
  DFF_X1 \next_pc_MW_reg_reg[22]  ( .D(n819), .CK(clk), .Q(n2202), .QN(n287)
         );
  DFF_X1 \pc_FD_reg_reg[22]  ( .D(n1631), .CK(clk), .Q(pc_FD_reg[22]), .QN()
         );
  DFF_X1 \pc_EX_reg_reg[22]  ( .D(n1630), .CK(clk), .Q(pc_EX_reg[22]), .QN()
         );
  DFF_X1 \next_pc_EX_reg_reg[23]  ( .D(n1684), .CK(clk), .Q(next_pc_EX_reg[23]), .QN(n290) );
  DFF_X1 \next_pc_MW_reg_reg[23]  ( .D(n816), .CK(clk), .Q(n2203), .QN(n289)
         );
  DFF_X1 \pc_FD_reg_reg[23]  ( .D(n1629), .CK(clk), .Q(pc_FD_reg[23]), .QN()
         );
  DFF_X1 \pc_EX_reg_reg[23]  ( .D(n1628), .CK(clk), .Q(pc_EX_reg[23]), .QN()
         );
  DFF_X1 \next_pc_EX_reg_reg[24]  ( .D(n1683), .CK(clk), .Q(next_pc_EX_reg[24]), .QN(n292) );
  DFF_X1 \next_pc_MW_reg_reg[24]  ( .D(n813), .CK(clk), .Q(n2204), .QN(n291)
         );
  DFF_X1 \pc_FD_reg_reg[24]  ( .D(n1627), .CK(clk), .Q(pc_FD_reg[24]), .QN()
         );
  DFF_X1 \pc_EX_reg_reg[24]  ( .D(n1626), .CK(clk), .Q(pc_EX_reg[24]), .QN()
         );
  DFF_X1 \next_pc_EX_reg_reg[25]  ( .D(n1682), .CK(clk), .Q(next_pc_EX_reg[25]), .QN(n294) );
  DFF_X1 \next_pc_MW_reg_reg[25]  ( .D(n810), .CK(clk), .Q(n2205), .QN(n293)
         );
  DFF_X1 \pc_FD_reg_reg[25]  ( .D(n1625), .CK(clk), .Q(pc_FD_reg[25]), .QN()
         );
  DFF_X1 \pc_EX_reg_reg[25]  ( .D(n1624), .CK(clk), .Q(pc_EX_reg[25]), .QN()
         );
  DFF_X1 \next_pc_EX_reg_reg[26]  ( .D(n1681), .CK(clk), .Q(next_pc_EX_reg[26]), .QN(n296) );
  DFF_X1 \next_pc_MW_reg_reg[26]  ( .D(n807), .CK(clk), .Q(n2206), .QN(n295)
         );
  DFF_X1 \pc_FD_reg_reg[26]  ( .D(n1623), .CK(clk), .Q(pc_FD_reg[26]), .QN()
         );
  DFF_X1 \pc_EX_reg_reg[26]  ( .D(n1622), .CK(clk), .Q(pc_EX_reg[26]), .QN()
         );
  DFF_X1 \next_pc_EX_reg_reg[27]  ( .D(n1680), .CK(clk), .Q(next_pc_EX_reg[27]), .QN(n298) );
  DFF_X1 \next_pc_MW_reg_reg[27]  ( .D(n804), .CK(clk), .Q(n2207), .QN(n297)
         );
  DFF_X1 \pc_FD_reg_reg[27]  ( .D(n1621), .CK(clk), .Q(pc_FD_reg[27]), .QN()
         );
  DFF_X1 \pc_EX_reg_reg[27]  ( .D(n1620), .CK(clk), .Q(pc_EX_reg[27]), .QN()
         );
  DFF_X1 \next_pc_EX_reg_reg[28]  ( .D(n1679), .CK(clk), .Q(next_pc_EX_reg[28]), .QN(n300) );
  DFF_X1 \next_pc_MW_reg_reg[28]  ( .D(n801), .CK(clk), .Q(n2208), .QN(n299)
         );
  DFF_X1 \pc_FD_reg_reg[28]  ( .D(n1619), .CK(clk), .Q(pc_FD_reg[28]), .QN()
         );
  DFF_X1 \pc_EX_reg_reg[28]  ( .D(n1618), .CK(clk), .Q(pc_EX_reg[28]), .QN()
         );
  DFF_X1 \next_pc_EX_reg_reg[29]  ( .D(n1678), .CK(clk), .Q(next_pc_EX_reg[29]), .QN(n302) );
  DFF_X1 \next_pc_MW_reg_reg[29]  ( .D(n798), .CK(clk), .Q(n2209), .QN(n301)
         );
  DFF_X1 \pc_FD_reg_reg[29]  ( .D(n1617), .CK(clk), .Q(pc_FD_reg[29]), .QN()
         );
  DFF_X1 \pc_EX_reg_reg[29]  ( .D(n1616), .CK(clk), .Q(pc_EX_reg[29]), .QN()
         );
  DFF_X1 \next_pc_EX_reg_reg[30]  ( .D(n1677), .CK(clk), .Q(next_pc_EX_reg[30]), .QN(n304) );
  DFF_X1 \next_pc_MW_reg_reg[30]  ( .D(n795), .CK(clk), .Q(n2210), .QN(n303)
         );
  DFF_X1 \pc_FD_reg_reg[30]  ( .D(n1615), .CK(clk), .Q(pc_FD_reg[30]), .QN()
         );
  DFF_X1 \pc_EX_reg_reg[30]  ( .D(n1614), .CK(clk), .Q(pc_EX_reg[30]), .QN()
         );
  DFF_X1 \next_pc_EX_reg_reg[31]  ( .D(n1676), .CK(clk), .Q(next_pc_EX_reg[31]), .QN(n306) );
  DFF_X1 \next_pc_MW_reg_reg[31]  ( .D(n792), .CK(clk), .Q(n2211), .QN(n305)
         );
  DFF_X1 \pc_EX_reg_reg[31]  ( .D(n1612), .CK(clk), .Q(pc_EX_reg[31]), .QN()
         );
  DFF_X1 \execution_result_MW_reg_reg[1]  ( .D(n1581), .CK(clk), .Q(
        execution_result_MW_reg[1]), .QN(n1206) );
  DFF_X1 \execution_result_MW_reg_reg[2]  ( .D(n1582), .CK(clk), .Q(
        execution_result_MW_reg[2]), .QN(n1205) );
  DFF_X1 \execution_result_MW_reg_reg[3]  ( .D(n1583), .CK(clk), .Q(
        execution_result_MW_reg[3]), .QN(n1204) );
  DFF_X1 \execution_result_MW_reg_reg[4]  ( .D(n1584), .CK(clk), .Q(
        execution_result_MW_reg[4]), .QN(n1203) );
  DFF_X1 \execution_result_MW_reg_reg[5]  ( .D(n1585), .CK(clk), .Q(
        execution_result_MW_reg[5]), .QN(n1202) );
  DFF_X1 \execution_result_MW_reg_reg[6]  ( .D(n1586), .CK(clk), .Q(
        execution_result_MW_reg[6]), .QN(n1201) );
  DFF_X1 \execution_result_MW_reg_reg[7]  ( .D(n1587), .CK(clk), .Q(
        execution_result_MW_reg[7]), .QN(n1200) );
  DFF_X1 \execution_result_MW_reg_reg[8]  ( .D(n1588), .CK(clk), .Q(
        execution_result_MW_reg[8]), .QN(n1199) );
  DFF_X1 \execution_result_MW_reg_reg[9]  ( .D(n1589), .CK(clk), .Q(
        execution_result_MW_reg[9]), .QN(n1198) );
  DFF_X1 \execution_result_MW_reg_reg[10]  ( .D(n1590), .CK(clk), .Q(
        execution_result_MW_reg[10]), .QN(n1197) );
  DFF_X1 \execution_result_MW_reg_reg[11]  ( .D(n1591), .CK(clk), .Q(
        execution_result_MW_reg[11]), .QN(n1196) );
  DFF_X1 \execution_result_MW_reg_reg[12]  ( .D(n1592), .CK(clk), .Q(
        execution_result_MW_reg[12]), .QN(n1195) );
  DFF_X1 \execution_result_MW_reg_reg[13]  ( .D(n1593), .CK(clk), .Q(
        execution_result_MW_reg[13]), .QN(n1194) );
  DFF_X1 \execution_result_MW_reg_reg[14]  ( .D(n1594), .CK(clk), .Q(
        execution_result_MW_reg[14]), .QN(n1193) );
  DFF_X1 \execution_result_MW_reg_reg[15]  ( .D(n1595), .CK(clk), .Q(
        execution_result_MW_reg[15]), .QN(n1192) );
  DFF_X1 \execution_result_MW_reg_reg[16]  ( .D(n1596), .CK(clk), .Q(
        execution_result_MW_reg[16]), .QN(n1191) );
  DFF_X1 \execution_result_MW_reg_reg[17]  ( .D(n1597), .CK(clk), .Q(
        execution_result_MW_reg[17]), .QN(n1190) );
  DFF_X1 \execution_result_MW_reg_reg[18]  ( .D(n1598), .CK(clk), .Q(
        execution_result_MW_reg[18]), .QN(n1189) );
  DFF_X1 \execution_result_MW_reg_reg[19]  ( .D(n1599), .CK(clk), .Q(
        execution_result_MW_reg[19]), .QN(n1188) );
  DFF_X1 \execution_result_MW_reg_reg[20]  ( .D(n1600), .CK(clk), .Q(
        execution_result_MW_reg[20]), .QN(n1187) );
  DFF_X1 \execution_result_MW_reg_reg[21]  ( .D(n1601), .CK(clk), .Q(
        execution_result_MW_reg[21]), .QN(n1186) );
  DFF_X1 \execution_result_MW_reg_reg[22]  ( .D(n1602), .CK(clk), .Q(
        execution_result_MW_reg[22]), .QN(n1185) );
  DFF_X1 \execution_result_MW_reg_reg[23]  ( .D(n1603), .CK(clk), .Q(
        execution_result_MW_reg[23]), .QN(n1184) );
  DFF_X1 \execution_result_MW_reg_reg[24]  ( .D(n1604), .CK(clk), .Q(
        execution_result_MW_reg[24]), .QN(n1183) );
  DFF_X1 \execution_result_MW_reg_reg[25]  ( .D(n1605), .CK(clk), .Q(
        execution_result_MW_reg[25]), .QN(n1182) );
  DFF_X1 \execution_result_MW_reg_reg[26]  ( .D(n1606), .CK(clk), .Q(
        execution_result_MW_reg[26]), .QN(n1181) );
  DFF_X1 \execution_result_MW_reg_reg[27]  ( .D(n1607), .CK(clk), .Q(
        execution_result_MW_reg[27]), .QN(n1180) );
  DFF_X1 \execution_result_MW_reg_reg[28]  ( .D(n1608), .CK(clk), .Q(
        execution_result_MW_reg[28]), .QN(n1179) );
  DFF_X1 \execution_result_MW_reg_reg[29]  ( .D(n1609), .CK(clk), .Q(
        execution_result_MW_reg[29]), .QN(n1178) );
  DFF_X1 \execution_result_MW_reg_reg[30]  ( .D(n1610), .CK(clk), .Q(
        execution_result_MW_reg[30]), .QN(n1177) );
  TBUF_X2 \write_data_MW_reg_tri[0]  ( .A(n657), .EN(n2471), .Z(
        write_data_MW_reg[0]) );
  TBUF_X2 \write_data_MW_reg_tri[1]  ( .A(n655), .EN(n2471), .Z(
        write_data_MW_reg[1]) );
  TBUF_X2 \write_data_MW_reg_tri[2]  ( .A(n653), .EN(n596), .Z(
        write_data_MW_reg[2]) );
  TBUF_X2 \write_data_MW_reg_tri[3]  ( .A(n651), .EN(n2471), .Z(
        write_data_MW_reg[3]) );
  TBUF_X2 \write_data_MW_reg_tri[4]  ( .A(n649), .EN(n596), .Z(
        write_data_MW_reg[4]) );
  TBUF_X2 \write_data_MW_reg_tri[5]  ( .A(n647), .EN(n596), .Z(
        write_data_MW_reg[5]) );
  TBUF_X2 \write_data_MW_reg_tri[6]  ( .A(n645), .EN(n596), .Z(
        write_data_MW_reg[6]) );
  TBUF_X2 \write_data_MW_reg_tri[7]  ( .A(n643), .EN(n596), .Z(
        write_data_MW_reg[7]) );
  TBUF_X2 \write_data_MW_reg_tri[8]  ( .A(n641), .EN(n596), .Z(
        write_data_MW_reg[8]) );
  TBUF_X2 \write_data_MW_reg_tri[9]  ( .A(n639), .EN(n596), .Z(
        write_data_MW_reg[9]) );
  TBUF_X2 \write_data_MW_reg_tri[10]  ( .A(n637), .EN(n596), .Z(
        write_data_MW_reg[10]) );
  TBUF_X2 \write_data_MW_reg_tri[11]  ( .A(n635), .EN(n2471), .Z(
        write_data_MW_reg[11]) );
  TBUF_X2 \write_data_MW_reg_tri[12]  ( .A(n633), .EN(n2471), .Z(
        write_data_MW_reg[12]) );
  TBUF_X2 \write_data_MW_reg_tri[13]  ( .A(n631), .EN(n2471), .Z(
        write_data_MW_reg[13]) );
  TBUF_X2 \write_data_MW_reg_tri[14]  ( .A(n629), .EN(n2471), .Z(
        write_data_MW_reg[14]) );
  TBUF_X2 \write_data_MW_reg_tri[15]  ( .A(n627), .EN(n2471), .Z(
        write_data_MW_reg[15]) );
  TBUF_X2 \write_data_MW_reg_tri[16]  ( .A(n625), .EN(n2471), .Z(
        write_data_MW_reg[16]) );
  TBUF_X2 \write_data_MW_reg_tri[17]  ( .A(n623), .EN(n2471), .Z(
        write_data_MW_reg[17]) );
  TBUF_X2 \write_data_MW_reg_tri[18]  ( .A(n621), .EN(n2471), .Z(
        write_data_MW_reg[18]) );
  TBUF_X2 \write_data_MW_reg_tri[19]  ( .A(n619), .EN(n2471), .Z(
        write_data_MW_reg[19]) );
  TBUF_X2 \write_data_MW_reg_tri[20]  ( .A(n617), .EN(n2471), .Z(
        write_data_MW_reg[20]) );
  TBUF_X2 \write_data_MW_reg_tri[21]  ( .A(n615), .EN(n2471), .Z(
        write_data_MW_reg[21]) );
  TBUF_X2 \write_data_MW_reg_tri[22]  ( .A(n613), .EN(n2471), .Z(
        write_data_MW_reg[22]) );
  TBUF_X2 \write_data_MW_reg_tri[23]  ( .A(n611), .EN(n2471), .Z(
        write_data_MW_reg[23]) );
  TBUF_X2 \write_data_MW_reg_tri[24]  ( .A(n609), .EN(n596), .Z(
        write_data_MW_reg[24]) );
  TBUF_X2 \write_data_MW_reg_tri[25]  ( .A(n607), .EN(n596), .Z(
        write_data_MW_reg[25]) );
  TBUF_X2 \write_data_MW_reg_tri[26]  ( .A(n605), .EN(n2471), .Z(
        write_data_MW_reg[26]) );
  TBUF_X2 \write_data_MW_reg_tri[27]  ( .A(n603), .EN(n596), .Z(
        write_data_MW_reg[27]) );
  TBUF_X2 \write_data_MW_reg_tri[28]  ( .A(n601), .EN(n596), .Z(
        write_data_MW_reg[28]) );
  TBUF_X2 \write_data_MW_reg_tri[29]  ( .A(n599), .EN(n2471), .Z(
        write_data_MW_reg[29]) );
  TBUF_X2 \write_data_MW_reg_tri[30]  ( .A(n597), .EN(n596), .Z(
        write_data_MW_reg[30]) );
  TBUF_X2 \write_data_MW_reg_tri[31]  ( .A(n595), .EN(n596), .Z(
        write_data_MW_reg[31]) );
  TBUF_X2 \rs2_EX_reg_tri[0]  ( .A(N559), .EN(N560), .Z(rs2_EX_reg[0]) );
  TBUF_X2 \rs2_EX_reg_tri[1]  ( .A(N556), .EN(N557), .Z(rs2_EX_reg[1]) );
  TBUF_X2 \rs2_EX_reg_tri[2]  ( .A(N553), .EN(N554), .Z(rs2_EX_reg[2]) );
  TBUF_X2 \rs2_EX_reg_tri[3]  ( .A(N550), .EN(N551), .Z(rs2_EX_reg[3]) );
  TBUF_X2 \rs2_EX_reg_tri[4]  ( .A(N547), .EN(N548), .Z(rs2_EX_reg[4]) );
  TBUF_X2 \rs2_EX_reg_tri[5]  ( .A(N544), .EN(N545), .Z(rs2_EX_reg[5]) );
  TBUF_X2 \rs2_EX_reg_tri[6]  ( .A(N541), .EN(N542), .Z(rs2_EX_reg[6]) );
  TBUF_X2 \rs2_EX_reg_tri[7]  ( .A(N538), .EN(N539), .Z(rs2_EX_reg[7]) );
  TBUF_X2 \rs2_EX_reg_tri[8]  ( .A(N535), .EN(N536), .Z(rs2_EX_reg[8]) );
  TBUF_X2 \rs2_EX_reg_tri[9]  ( .A(N532), .EN(N533), .Z(rs2_EX_reg[9]) );
  TBUF_X2 \rs2_EX_reg_tri[10]  ( .A(N529), .EN(N530), .Z(rs2_EX_reg[10]) );
  TBUF_X2 \rs2_EX_reg_tri[11]  ( .A(N526), .EN(N527), .Z(rs2_EX_reg[11]) );
  TBUF_X2 \rs2_EX_reg_tri[12]  ( .A(N523), .EN(N524), .Z(rs2_EX_reg[12]) );
  TBUF_X2 \rs2_EX_reg_tri[13]  ( .A(N520), .EN(N521), .Z(rs2_EX_reg[13]) );
  TBUF_X2 \rs2_EX_reg_tri[14]  ( .A(N517), .EN(N518), .Z(rs2_EX_reg[14]) );
  TBUF_X2 \rs2_EX_reg_tri[15]  ( .A(N514), .EN(N515), .Z(rs2_EX_reg[15]) );
  TBUF_X2 \rs2_EX_reg_tri[16]  ( .A(N511), .EN(N512), .Z(rs2_EX_reg[16]) );
  TBUF_X2 \rs2_EX_reg_tri[17]  ( .A(N508), .EN(N509), .Z(rs2_EX_reg[17]) );
  TBUF_X2 \rs2_EX_reg_tri[18]  ( .A(N505), .EN(N506), .Z(rs2_EX_reg[18]) );
  TBUF_X2 \rs2_EX_reg_tri[19]  ( .A(N502), .EN(N503), .Z(rs2_EX_reg[19]) );
  TBUF_X2 \rs2_EX_reg_tri[20]  ( .A(N499), .EN(N500), .Z(rs2_EX_reg[20]) );
  TBUF_X2 \rs2_EX_reg_tri[21]  ( .A(N496), .EN(N497), .Z(rs2_EX_reg[21]) );
  TBUF_X2 \rs2_EX_reg_tri[22]  ( .A(N493), .EN(N494), .Z(rs2_EX_reg[22]) );
  TBUF_X2 \rs2_EX_reg_tri[23]  ( .A(N490), .EN(N491), .Z(rs2_EX_reg[23]) );
  TBUF_X2 \rs2_EX_reg_tri[24]  ( .A(N487), .EN(N488), .Z(rs2_EX_reg[24]) );
  TBUF_X2 \rs2_EX_reg_tri[25]  ( .A(N484), .EN(N485), .Z(rs2_EX_reg[25]) );
  TBUF_X2 \rs2_EX_reg_tri[26]  ( .A(N481), .EN(N482), .Z(rs2_EX_reg[26]) );
  TBUF_X2 \rs2_EX_reg_tri[27]  ( .A(N478), .EN(N479), .Z(rs2_EX_reg[27]) );
  TBUF_X2 \rs2_EX_reg_tri[28]  ( .A(N475), .EN(N476), .Z(rs2_EX_reg[28]) );
  TBUF_X2 \rs2_EX_reg_tri[29]  ( .A(N472), .EN(N473), .Z(rs2_EX_reg[29]) );
  TBUF_X2 \rs2_EX_reg_tri[30]  ( .A(N469), .EN(N470), .Z(rs2_EX_reg[30]) );
  TBUF_X2 \rs2_EX_reg_tri[31]  ( .A(N466), .EN(N467), .Z(rs2_EX_reg[31]) );
  TBUF_X2 \rs1_EX_reg_tri[2]  ( .A(N457), .EN(N458), .Z(rs1_EX_reg[2]) );
  TBUF_X2 \rs1_EX_reg_tri[3]  ( .A(N454), .EN(N455), .Z(rs1_EX_reg[3]) );
  TBUF_X2 \rs1_EX_reg_tri[4]  ( .A(N451), .EN(N452), .Z(rs1_EX_reg[4]) );
  TBUF_X2 \rs1_EX_reg_tri[5]  ( .A(N448), .EN(N449), .Z(rs1_EX_reg[5]) );
  TBUF_X2 \rs1_EX_reg_tri[6]  ( .A(N445), .EN(N446), .Z(rs1_EX_reg[6]) );
  TBUF_X2 \rs1_EX_reg_tri[7]  ( .A(N442), .EN(N443), .Z(rs1_EX_reg[7]) );
  TBUF_X2 \rs1_EX_reg_tri[8]  ( .A(N439), .EN(N440), .Z(rs1_EX_reg[8]) );
  TBUF_X2 \rs1_EX_reg_tri[9]  ( .A(N436), .EN(N437), .Z(rs1_EX_reg[9]) );
  TBUF_X2 \rs1_EX_reg_tri[11]  ( .A(N430), .EN(N431), .Z(rs1_EX_reg[11]) );
  TBUF_X2 \rs1_EX_reg_tri[12]  ( .A(N427), .EN(N428), .Z(rs1_EX_reg[12]) );
  TBUF_X2 \rs1_EX_reg_tri[13]  ( .A(N424), .EN(N425), .Z(rs1_EX_reg[13]) );
  TBUF_X2 \rs1_EX_reg_tri[14]  ( .A(N421), .EN(N422), .Z(rs1_EX_reg[14]) );
  TBUF_X2 \rs1_EX_reg_tri[15]  ( .A(N418), .EN(N419), .Z(rs1_EX_reg[15]) );
  TBUF_X2 \rs1_EX_reg_tri[16]  ( .A(N415), .EN(N416), .Z(rs1_EX_reg[16]) );
  TBUF_X2 \rs1_EX_reg_tri[17]  ( .A(N412), .EN(N413), .Z(rs1_EX_reg[17]) );
  TBUF_X2 \rs1_EX_reg_tri[18]  ( .A(N409), .EN(N410), .Z(rs1_EX_reg[18]) );
  TBUF_X2 \rs1_EX_reg_tri[19]  ( .A(N406), .EN(N407), .Z(rs1_EX_reg[19]) );
  TBUF_X2 \rs1_EX_reg_tri[20]  ( .A(N403), .EN(N404), .Z(rs1_EX_reg[20]) );
  TBUF_X2 \rs1_EX_reg_tri[21]  ( .A(N400), .EN(N401), .Z(rs1_EX_reg[21]) );
  TBUF_X2 \rs1_EX_reg_tri[22]  ( .A(N397), .EN(N398), .Z(rs1_EX_reg[22]) );
  TBUF_X2 \rs1_EX_reg_tri[23]  ( .A(N394), .EN(N395), .Z(rs1_EX_reg[23]) );
  TBUF_X2 \rs1_EX_reg_tri[24]  ( .A(N391), .EN(N392), .Z(rs1_EX_reg[24]) );
  TBUF_X2 \rs1_EX_reg_tri[25]  ( .A(N388), .EN(N389), .Z(rs1_EX_reg[25]) );
  TBUF_X2 \rs1_EX_reg_tri[26]  ( .A(N385), .EN(N386), .Z(rs1_EX_reg[26]) );
  TBUF_X2 \rs1_EX_reg_tri[27]  ( .A(N382), .EN(N383), .Z(rs1_EX_reg[27]) );
  TBUF_X2 \rs1_EX_reg_tri[28]  ( .A(N379), .EN(N380), .Z(rs1_EX_reg[28]) );
  TBUF_X2 \rs1_EX_reg_tri[29]  ( .A(N376), .EN(N377), .Z(rs1_EX_reg[29]) );
  TBUF_X2 \rs1_EX_reg_tri[30]  ( .A(N373), .EN(N374), .Z(rs1_EX_reg[30]) );
  TBUF_X2 \rs1_EX_reg_tri[31]  ( .A(N370), .EN(N371), .Z(rs1_EX_reg[31]) );
  AOI22_X1 U6 ( .A1(n2447), .A2(n1), .B1(n211), .B2(n2441), .ZN(n1123) );
  AOI22_X1 U10 ( .A1(n2447), .A2(n3), .B1(n213), .B2(n2437), .ZN(n1121) );
  AOI22_X1 U12 ( .A1(n2447), .A2(n4), .B1(n214), .B2(n2441), .ZN(n1120) );
  AOI22_X1 U14 ( .A1(n2447), .A2(n5), .B1(n215), .B2(n2439), .ZN(n1119) );
  AOI22_X1 U16 ( .A1(n2445), .A2(n6), .B1(n216), .B2(n2437), .ZN(n1118) );
  AOI22_X1 U18 ( .A1(n2446), .A2(n7), .B1(n217), .B2(n2441), .ZN(n1117) );
  AOI22_X1 U20 ( .A1(n2447), .A2(n8), .B1(n218), .B2(n2441), .ZN(n1116) );
  AOI22_X1 U24 ( .A1(n2446), .A2(n10), .B1(n220), .B2(n2441), .ZN(n1114) );
  AOI22_X1 U26 ( .A1(n2447), .A2(n11), .B1(n221), .B2(n2441), .ZN(n1113) );
  AOI22_X1 U28 ( .A1(n2447), .A2(n12), .B1(n222), .B2(n2441), .ZN(n1112) );
  AOI22_X1 U30 ( .A1(n2447), .A2(n13), .B1(n223), .B2(n2438), .ZN(n1111) );
  AOI22_X1 U32 ( .A1(n2447), .A2(n14), .B1(n224), .B2(n2441), .ZN(n1110) );
  AOI22_X1 U34 ( .A1(n2446), .A2(n15), .B1(n225), .B2(n2438), .ZN(n1109) );
  AOI22_X1 U38 ( .A1(n2446), .A2(n17), .B1(n227), .B2(n2441), .ZN(n1107) );
  AOI22_X1 U40 ( .A1(n2446), .A2(n18), .B1(n228), .B2(n2443), .ZN(n1106) );
  AOI22_X1 U42 ( .A1(n2445), .A2(n19), .B1(n229), .B2(n2441), .ZN(n1105) );
  AOI22_X1 U44 ( .A1(n2446), .A2(n20), .B1(n230), .B2(n2441), .ZN(n1104) );
  AOI22_X1 U46 ( .A1(n2446), .A2(n21), .B1(n231), .B2(n2441), .ZN(n1103) );
  AOI22_X1 U48 ( .A1(n2446), .A2(n22), .B1(n232), .B2(n2440), .ZN(n1102) );
  AOI22_X1 U50 ( .A1(n2445), .A2(n23), .B1(n233), .B2(n2443), .ZN(n1101) );
  AOI22_X1 U54 ( .A1(n2445), .A2(n25), .B1(n235), .B2(n2439), .ZN(n1099) );
  AOI22_X1 U56 ( .A1(n2445), .A2(n26), .B1(n236), .B2(n2440), .ZN(n1098) );
  AOI22_X1 U58 ( .A1(n2445), .A2(n27), .B1(n237), .B2(n2441), .ZN(n1097) );
  AOI22_X1 U60 ( .A1(n2445), .A2(n28), .B1(n238), .B2(n2441), .ZN(n1096) );
  AOI22_X1 U62 ( .A1(n2445), .A2(n29), .B1(n239), .B2(n2440), .ZN(n1095) );
  AOI22_X1 U64 ( .A1(n2445), .A2(n30), .B1(n240), .B2(n2441), .ZN(n1094) );
  AOI22_X1 U66 ( .A1(n2445), .A2(n31), .B1(n241), .B2(n2437), .ZN(n1093) );
  AOI22_X1 U68 ( .A1(n2445), .A2(n32), .B1(n242), .B2(n2441), .ZN(n1092) );
  MUX2_X1 U69 ( .A(csr_rd_EX_wire[0]), .B(csr_rd_MW_reg[0]), .S(n2442), .Z(
        n950) );
  MUX2_X1 U70 ( .A(csr_rd_EX_wire[1]), .B(csr_rd_MW_reg[1]), .S(n2440), .Z(
        n949) );
  MUX2_X1 U71 ( .A(csr_rd_EX_wire[2]), .B(csr_rd_MW_reg[2]), .S(n2442), .Z(
        n948) );
  MUX2_X1 U72 ( .A(csr_rd_EX_wire[3]), .B(csr_rd_MW_reg[3]), .S(n2440), .Z(
        n947) );
  MUX2_X1 U73 ( .A(csr_rd_EX_wire[4]), .B(csr_rd_MW_reg[4]), .S(n2439), .Z(
        n946) );
  MUX2_X1 U74 ( .A(csr_rd_EX_wire[5]), .B(csr_rd_MW_reg[5]), .S(n2437), .Z(
        n945) );
  MUX2_X1 U75 ( .A(csr_rd_EX_wire[6]), .B(csr_rd_MW_reg[6]), .S(n2438), .Z(
        n944) );
  MUX2_X1 U76 ( .A(csr_rd_EX_wire[7]), .B(csr_rd_MW_reg[7]), .S(n2442), .Z(
        n943) );
  MUX2_X1 U77 ( .A(csr_rd_EX_wire[8]), .B(csr_rd_MW_reg[8]), .S(n2440), .Z(
        n942) );
  MUX2_X1 U78 ( .A(csr_rd_EX_wire[9]), .B(csr_rd_MW_reg[9]), .S(n2440), .Z(
        n941) );
  MUX2_X1 U79 ( .A(csr_rd_EX_wire[10]), .B(csr_rd_MW_reg[10]), .S(n2440), .Z(
        n940) );
  MUX2_X1 U80 ( .A(csr_rd_EX_wire[11]), .B(csr_rd_MW_reg[11]), .S(n2440), .Z(
        n939) );
  MUX2_X1 U81 ( .A(csr_rd_EX_wire[12]), .B(csr_rd_MW_reg[12]), .S(n2440), .Z(
        n938) );
  MUX2_X1 U82 ( .A(csr_rd_EX_wire[13]), .B(csr_rd_MW_reg[13]), .S(n2440), .Z(
        n937) );
  MUX2_X1 U83 ( .A(csr_rd_EX_wire[14]), .B(csr_rd_MW_reg[14]), .S(n2440), .Z(
        n936) );
  MUX2_X1 U84 ( .A(csr_rd_EX_wire[15]), .B(csr_rd_MW_reg[15]), .S(n2440), .Z(
        n935) );
  MUX2_X1 U85 ( .A(csr_rd_EX_wire[16]), .B(csr_rd_MW_reg[16]), .S(n2440), .Z(
        n934) );
  MUX2_X1 U86 ( .A(csr_rd_EX_wire[17]), .B(csr_rd_MW_reg[17]), .S(n2440), .Z(
        n933) );
  MUX2_X1 U87 ( .A(csr_rd_EX_wire[18]), .B(csr_rd_MW_reg[18]), .S(n2440), .Z(
        n932) );
  MUX2_X1 U88 ( .A(csr_rd_EX_wire[19]), .B(csr_rd_MW_reg[19]), .S(n2440), .Z(
        n931) );
  MUX2_X1 U89 ( .A(csr_rd_EX_wire[20]), .B(csr_rd_MW_reg[20]), .S(n2439), .Z(
        n930) );
  MUX2_X1 U90 ( .A(csr_rd_EX_wire[21]), .B(csr_rd_MW_reg[21]), .S(n2439), .Z(
        n929) );
  MUX2_X1 U91 ( .A(csr_rd_EX_wire[22]), .B(csr_rd_MW_reg[22]), .S(n2439), .Z(
        n928) );
  MUX2_X1 U92 ( .A(csr_rd_EX_wire[23]), .B(csr_rd_MW_reg[23]), .S(n2439), .Z(
        n927) );
  MUX2_X1 U93 ( .A(csr_rd_EX_wire[24]), .B(csr_rd_MW_reg[24]), .S(n2439), .Z(
        n926) );
  MUX2_X1 U94 ( .A(csr_rd_EX_wire[25]), .B(csr_rd_MW_reg[25]), .S(n2439), .Z(
        n925) );
  MUX2_X1 U95 ( .A(csr_rd_EX_wire[26]), .B(csr_rd_MW_reg[26]), .S(n2439), .Z(
        n924) );
  MUX2_X1 U96 ( .A(csr_rd_EX_wire[27]), .B(csr_rd_MW_reg[27]), .S(n2439), .Z(
        n923) );
  MUX2_X1 U97 ( .A(csr_rd_EX_wire[28]), .B(csr_rd_MW_reg[28]), .S(n2439), .Z(
        n922) );
  MUX2_X1 U98 ( .A(csr_rd_EX_wire[29]), .B(csr_rd_MW_reg[29]), .S(n2439), .Z(
        n921) );
  MUX2_X1 U99 ( .A(csr_rd_EX_wire[30]), .B(csr_rd_MW_reg[30]), .S(n2439), .Z(
        n920) );
  MUX2_X1 U100 ( .A(csr_rd_EX_wire[31]), .B(csr_rd_MW_reg[31]), .S(n2437), .Z(
        n919) );
  OAI22_X1 U107 ( .A1(n2440), .A2(address_EX_wire[3]), .B1(address_MW_reg[3]), 
        .B2(n2444), .ZN(n36) );
  INV_X1 U108 ( .A(n36), .ZN(n915) );
  OAI22_X1 U109 ( .A1(n2438), .A2(address_EX_wire[4]), .B1(address_MW_reg[4]), 
        .B2(n2444), .ZN(n37) );
  INV_X1 U110 ( .A(n37), .ZN(n914) );
  OAI22_X1 U111 ( .A1(n2442), .A2(address_EX_wire[5]), .B1(address_MW_reg[5]), 
        .B2(n2444), .ZN(n38) );
  INV_X1 U112 ( .A(n38), .ZN(n913) );
  OAI22_X1 U113 ( .A1(n2439), .A2(address_EX_wire[6]), .B1(address_MW_reg[6]), 
        .B2(n2444), .ZN(n39) );
  INV_X1 U114 ( .A(n39), .ZN(n912) );
  OAI22_X1 U115 ( .A1(n2437), .A2(address_EX_wire[7]), .B1(address_MW_reg[7]), 
        .B2(n2444), .ZN(n40) );
  INV_X1 U116 ( .A(n40), .ZN(n911) );
  AOI22_X1 U165 ( .A1(n2445), .A2(n244), .B1(n243), .B2(n2439), .ZN(n885) );
  AOI22_X1 U166 ( .A1(n2445), .A2(n246), .B1(n245), .B2(n2443), .ZN(n882) );
  AOI22_X1 U167 ( .A1(n2446), .A2(n248), .B1(n247), .B2(n2441), .ZN(n879) );
  AOI22_X1 U168 ( .A1(n2445), .A2(n250), .B1(n249), .B2(n2442), .ZN(n876) );
  AOI22_X1 U169 ( .A1(n2445), .A2(n252), .B1(n251), .B2(n2441), .ZN(n873) );
  AOI22_X1 U170 ( .A1(n2445), .A2(n254), .B1(n253), .B2(n2443), .ZN(n870) );
  AOI22_X1 U171 ( .A1(n2445), .A2(n256), .B1(n255), .B2(n2442), .ZN(n867) );
  AOI22_X1 U172 ( .A1(n2446), .A2(n258), .B1(n257), .B2(n2442), .ZN(n864) );
  AOI22_X1 U173 ( .A1(n2445), .A2(n260), .B1(n259), .B2(n2442), .ZN(n861) );
  AOI22_X1 U174 ( .A1(n2445), .A2(n262), .B1(n261), .B2(n2442), .ZN(n858) );
  AOI22_X1 U175 ( .A1(n2445), .A2(n264), .B1(n263), .B2(n2442), .ZN(n855) );
  AOI22_X1 U176 ( .A1(n2445), .A2(n266), .B1(n265), .B2(n2442), .ZN(n852) );
  AOI22_X1 U177 ( .A1(n2445), .A2(n268), .B1(n267), .B2(n2442), .ZN(n849) );
  AOI22_X1 U178 ( .A1(n2445), .A2(n270), .B1(n269), .B2(n2442), .ZN(n846) );
  AOI22_X1 U179 ( .A1(n2446), .A2(n272), .B1(n271), .B2(n2442), .ZN(n843) );
  AOI22_X1 U180 ( .A1(n2445), .A2(n274), .B1(n273), .B2(n2442), .ZN(n840) );
  AOI22_X1 U181 ( .A1(n2446), .A2(n276), .B1(n275), .B2(n2442), .ZN(n837) );
  AOI22_X1 U182 ( .A1(n2445), .A2(n278), .B1(n277), .B2(n2442), .ZN(n834) );
  AOI22_X1 U183 ( .A1(n2446), .A2(n280), .B1(n279), .B2(n2442), .ZN(n831) );
  AOI22_X1 U184 ( .A1(n2445), .A2(n282), .B1(n281), .B2(n2439), .ZN(n828) );
  AOI22_X1 U185 ( .A1(n2445), .A2(n284), .B1(n283), .B2(n2443), .ZN(n825) );
  AOI22_X1 U186 ( .A1(n2446), .A2(n286), .B1(n285), .B2(n2442), .ZN(n822) );
  AOI22_X1 U187 ( .A1(n2445), .A2(n288), .B1(n287), .B2(n2443), .ZN(n819) );
  AOI22_X1 U188 ( .A1(n2445), .A2(n290), .B1(n289), .B2(n2443), .ZN(n816) );
  AOI22_X1 U189 ( .A1(n2446), .A2(n292), .B1(n291), .B2(n2441), .ZN(n813) );
  AOI22_X1 U190 ( .A1(n2444), .A2(n294), .B1(n293), .B2(n2443), .ZN(n810) );
  AOI22_X1 U191 ( .A1(n2445), .A2(n296), .B1(n295), .B2(n2441), .ZN(n807) );
  AOI22_X1 U192 ( .A1(n2445), .A2(n298), .B1(n297), .B2(n2443), .ZN(n804) );
  AOI22_X1 U193 ( .A1(n2445), .A2(n300), .B1(n299), .B2(n2437), .ZN(n801) );
  AOI22_X1 U194 ( .A1(n2445), .A2(n302), .B1(n301), .B2(n2441), .ZN(n798) );
  AOI22_X1 U195 ( .A1(n2445), .A2(n304), .B1(n303), .B2(n2441), .ZN(n795) );
  AOI22_X1 U196 ( .A1(n2445), .A2(n306), .B1(n305), .B2(n2438), .ZN(n792) );
  NAND3_X1 U199 ( .A1(n1565), .A2(opcode_MW_reg[2]), .A3(opcode_MW_reg[4]), 
        .ZN(n66) );
  AOI22_X1 U203 ( .A1(n202), .A2(immediate_MW_reg[31]), .B1(n201), .B2(
        address_MW_reg[31]), .ZN(n71) );
  NAND3_X1 U205 ( .A1(n1210), .A2(n789), .A3(opcode_MW_reg[4]), .ZN(n67) );
  NOR3_X1 U207 ( .A1(n790), .A2(n1208), .A3(n67), .ZN(n203) );
  AOI22_X1 U208 ( .A1(n204), .A2(execution_result_MW_reg[31]), .B1(n2013), 
        .B2(csr_rd_MW_reg[31]), .ZN(n70) );
  AOI22_X1 U212 ( .A1(n2014), .A2(n2211), .B1(n2009), .B2(
        load_data_MW_wire[31]), .ZN(n69) );
  NAND3_X1 U213 ( .A1(n71), .A2(n70), .A3(n69), .ZN(n595) );
  NAND2_X1 U214 ( .A1(n1210), .A2(n1209), .ZN(n80) );
  OAI221_X1 U215 ( .B1(opcode_MW_reg[6]), .B2(n1209), .C1(n790), .C2(
        opcode_MW_reg[4]), .A(opcode_MW_reg[2]), .ZN(n79) );
  NOR2_X1 U216 ( .A1(n789), .A2(opcode_MW_reg[6]), .ZN(n77) );
  OAI22_X1 U217 ( .A1(n1209), .A2(n789), .B1(n790), .B2(opcode_MW_reg[5]), 
        .ZN(n76) );
  NOR4_X1 U218 ( .A1(n787), .A2(n77), .A3(n788), .A4(n76), .ZN(n78) );
  AOI22_X1 U220 ( .A1(n202), .A2(immediate_MW_reg[30]), .B1(n201), .B2(
        address_MW_reg[30]), .ZN(n84) );
  AOI22_X1 U221 ( .A1(n204), .A2(execution_result_MW_reg[30]), .B1(n2013), 
        .B2(csr_rd_MW_reg[30]), .ZN(n83) );
  AOI22_X1 U223 ( .A1(n2014), .A2(n2210), .B1(n2009), .B2(
        load_data_MW_wire[30]), .ZN(n82) );
  NAND3_X1 U224 ( .A1(n84), .A2(n83), .A3(n82), .ZN(n597) );
  AOI22_X1 U225 ( .A1(n202), .A2(immediate_MW_reg[29]), .B1(n201), .B2(
        address_MW_reg[29]), .ZN(n88) );
  AOI22_X1 U226 ( .A1(n204), .A2(execution_result_MW_reg[29]), .B1(n2013), 
        .B2(csr_rd_MW_reg[29]), .ZN(n87) );
  AOI22_X1 U228 ( .A1(n2014), .A2(n2209), .B1(n2009), .B2(
        load_data_MW_wire[29]), .ZN(n86) );
  NAND3_X1 U229 ( .A1(n88), .A2(n87), .A3(n86), .ZN(n599) );
  AOI22_X1 U230 ( .A1(n202), .A2(immediate_MW_reg[28]), .B1(n201), .B2(
        address_MW_reg[28]), .ZN(n92) );
  AOI22_X1 U231 ( .A1(n204), .A2(execution_result_MW_reg[28]), .B1(n2013), 
        .B2(csr_rd_MW_reg[28]), .ZN(n91) );
  AOI22_X1 U233 ( .A1(n2014), .A2(n2208), .B1(n2009), .B2(
        load_data_MW_wire[28]), .ZN(n90) );
  NAND3_X1 U234 ( .A1(n92), .A2(n91), .A3(n90), .ZN(n601) );
  AOI22_X1 U235 ( .A1(n202), .A2(immediate_MW_reg[27]), .B1(n201), .B2(
        address_MW_reg[27]), .ZN(n96) );
  AOI22_X1 U236 ( .A1(n204), .A2(execution_result_MW_reg[27]), .B1(n2013), 
        .B2(csr_rd_MW_reg[27]), .ZN(n95) );
  AOI22_X1 U238 ( .A1(n2014), .A2(n2207), .B1(n2009), .B2(
        load_data_MW_wire[27]), .ZN(n94) );
  NAND3_X1 U239 ( .A1(n96), .A2(n95), .A3(n94), .ZN(n603) );
  AOI22_X1 U240 ( .A1(n202), .A2(immediate_MW_reg[26]), .B1(n201), .B2(
        address_MW_reg[26]), .ZN(n100) );
  AOI22_X1 U241 ( .A1(n204), .A2(execution_result_MW_reg[26]), .B1(n2013), 
        .B2(csr_rd_MW_reg[26]), .ZN(n99) );
  AOI22_X1 U243 ( .A1(n2014), .A2(n2206), .B1(n2009), .B2(
        load_data_MW_wire[26]), .ZN(n98) );
  NAND3_X1 U244 ( .A1(n100), .A2(n99), .A3(n98), .ZN(n605) );
  AOI22_X1 U245 ( .A1(n202), .A2(immediate_MW_reg[25]), .B1(n201), .B2(
        address_MW_reg[25]), .ZN(n104) );
  AOI22_X1 U246 ( .A1(n204), .A2(execution_result_MW_reg[25]), .B1(n2013), 
        .B2(csr_rd_MW_reg[25]), .ZN(n103) );
  AOI22_X1 U248 ( .A1(n2014), .A2(n2205), .B1(n2009), .B2(
        load_data_MW_wire[25]), .ZN(n102) );
  NAND3_X1 U249 ( .A1(n104), .A2(n103), .A3(n102), .ZN(n607) );
  AOI22_X1 U250 ( .A1(n202), .A2(immediate_MW_reg[24]), .B1(n201), .B2(
        address_MW_reg[24]), .ZN(n108) );
  AOI22_X1 U251 ( .A1(n204), .A2(execution_result_MW_reg[24]), .B1(n2013), 
        .B2(csr_rd_MW_reg[24]), .ZN(n107) );
  AOI22_X1 U253 ( .A1(n2014), .A2(n2204), .B1(n2009), .B2(
        load_data_MW_wire[24]), .ZN(n106) );
  NAND3_X1 U254 ( .A1(n108), .A2(n107), .A3(n106), .ZN(n609) );
  AOI22_X1 U255 ( .A1(n202), .A2(immediate_MW_reg[23]), .B1(n201), .B2(
        address_MW_reg[23]), .ZN(n112) );
  AOI22_X1 U256 ( .A1(n204), .A2(execution_result_MW_reg[23]), .B1(n2013), 
        .B2(csr_rd_MW_reg[23]), .ZN(n111) );
  AOI22_X1 U258 ( .A1(n2014), .A2(n2203), .B1(n2009), .B2(
        load_data_MW_wire[23]), .ZN(n110) );
  NAND3_X1 U259 ( .A1(n112), .A2(n111), .A3(n110), .ZN(n611) );
  AOI22_X1 U260 ( .A1(n202), .A2(immediate_MW_reg[22]), .B1(n201), .B2(
        address_MW_reg[22]), .ZN(n116) );
  AOI22_X1 U261 ( .A1(n204), .A2(execution_result_MW_reg[22]), .B1(n2013), 
        .B2(csr_rd_MW_reg[22]), .ZN(n115) );
  AOI22_X1 U263 ( .A1(n2014), .A2(n2202), .B1(n2009), .B2(
        load_data_MW_wire[22]), .ZN(n114) );
  NAND3_X1 U264 ( .A1(n116), .A2(n115), .A3(n114), .ZN(n613) );
  AOI22_X1 U265 ( .A1(n202), .A2(immediate_MW_reg[21]), .B1(n201), .B2(
        address_MW_reg[21]), .ZN(n120) );
  AOI22_X1 U266 ( .A1(n204), .A2(execution_result_MW_reg[21]), .B1(n2013), 
        .B2(csr_rd_MW_reg[21]), .ZN(n119) );
  AOI22_X1 U268 ( .A1(n2014), .A2(n2201), .B1(n2009), .B2(
        load_data_MW_wire[21]), .ZN(n118) );
  NAND3_X1 U269 ( .A1(n120), .A2(n119), .A3(n118), .ZN(n615) );
  AOI22_X1 U270 ( .A1(n202), .A2(immediate_MW_reg[20]), .B1(n201), .B2(
        address_MW_reg[20]), .ZN(n124) );
  AOI22_X1 U271 ( .A1(n204), .A2(execution_result_MW_reg[20]), .B1(n2013), 
        .B2(csr_rd_MW_reg[20]), .ZN(n123) );
  AOI22_X1 U273 ( .A1(n2014), .A2(n2200), .B1(n2009), .B2(
        load_data_MW_wire[20]), .ZN(n122) );
  NAND3_X1 U274 ( .A1(n124), .A2(n123), .A3(n122), .ZN(n617) );
  AOI22_X1 U275 ( .A1(n202), .A2(immediate_MW_reg[19]), .B1(n201), .B2(
        address_MW_reg[19]), .ZN(n128) );
  AOI22_X1 U276 ( .A1(n204), .A2(execution_result_MW_reg[19]), .B1(n2013), 
        .B2(csr_rd_MW_reg[19]), .ZN(n127) );
  AOI22_X1 U278 ( .A1(n2014), .A2(n2199), .B1(n2009), .B2(
        load_data_MW_wire[19]), .ZN(n126) );
  NAND3_X1 U279 ( .A1(n128), .A2(n127), .A3(n126), .ZN(n619) );
  AOI22_X1 U280 ( .A1(n202), .A2(immediate_MW_reg[18]), .B1(n201), .B2(
        address_MW_reg[18]), .ZN(n132) );
  AOI22_X1 U281 ( .A1(n204), .A2(execution_result_MW_reg[18]), .B1(n2013), 
        .B2(csr_rd_MW_reg[18]), .ZN(n131) );
  AOI22_X1 U283 ( .A1(n2014), .A2(n2198), .B1(n2009), .B2(
        load_data_MW_wire[18]), .ZN(n130) );
  NAND3_X1 U284 ( .A1(n132), .A2(n131), .A3(n130), .ZN(n621) );
  AOI22_X1 U285 ( .A1(n202), .A2(immediate_MW_reg[17]), .B1(n201), .B2(
        address_MW_reg[17]), .ZN(n136) );
  AOI22_X1 U286 ( .A1(n204), .A2(execution_result_MW_reg[17]), .B1(n2013), 
        .B2(csr_rd_MW_reg[17]), .ZN(n135) );
  AOI22_X1 U288 ( .A1(n2014), .A2(n2197), .B1(n2009), .B2(
        load_data_MW_wire[17]), .ZN(n134) );
  NAND3_X1 U289 ( .A1(n136), .A2(n135), .A3(n134), .ZN(n623) );
  AOI22_X1 U290 ( .A1(n202), .A2(immediate_MW_reg[16]), .B1(n201), .B2(
        address_MW_reg[16]), .ZN(n140) );
  AOI22_X1 U291 ( .A1(n204), .A2(execution_result_MW_reg[16]), .B1(n2013), 
        .B2(csr_rd_MW_reg[16]), .ZN(n139) );
  AOI22_X1 U293 ( .A1(n2014), .A2(n2196), .B1(n2009), .B2(
        load_data_MW_wire[16]), .ZN(n138) );
  NAND3_X1 U294 ( .A1(n140), .A2(n139), .A3(n138), .ZN(n625) );
  AOI22_X1 U295 ( .A1(n202), .A2(immediate_MW_reg[15]), .B1(n201), .B2(
        address_MW_reg[15]), .ZN(n144) );
  AOI22_X1 U296 ( .A1(n204), .A2(execution_result_MW_reg[15]), .B1(n2013), 
        .B2(csr_rd_MW_reg[15]), .ZN(n143) );
  AOI22_X1 U298 ( .A1(n2014), .A2(n2195), .B1(n2009), .B2(
        load_data_MW_wire[15]), .ZN(n142) );
  NAND3_X1 U299 ( .A1(n144), .A2(n143), .A3(n142), .ZN(n627) );
  AOI22_X1 U300 ( .A1(n202), .A2(immediate_MW_reg[14]), .B1(n201), .B2(
        address_MW_reg[14]), .ZN(n148) );
  AOI22_X1 U301 ( .A1(n204), .A2(execution_result_MW_reg[14]), .B1(n2013), 
        .B2(csr_rd_MW_reg[14]), .ZN(n147) );
  AOI22_X1 U303 ( .A1(n2014), .A2(n2194), .B1(n2009), .B2(
        load_data_MW_wire[14]), .ZN(n146) );
  NAND3_X1 U304 ( .A1(n148), .A2(n147), .A3(n146), .ZN(n629) );
  AOI22_X1 U305 ( .A1(n202), .A2(immediate_MW_reg[13]), .B1(n201), .B2(
        address_MW_reg[13]), .ZN(n152) );
  AOI22_X1 U306 ( .A1(n204), .A2(execution_result_MW_reg[13]), .B1(n2013), 
        .B2(csr_rd_MW_reg[13]), .ZN(n151) );
  AOI22_X1 U308 ( .A1(n2014), .A2(n2193), .B1(n2009), .B2(
        load_data_MW_wire[13]), .ZN(n150) );
  NAND3_X1 U309 ( .A1(n152), .A2(n151), .A3(n150), .ZN(n631) );
  AOI22_X1 U310 ( .A1(n202), .A2(immediate_MW_reg[12]), .B1(n201), .B2(
        address_MW_reg[12]), .ZN(n156) );
  AOI22_X1 U311 ( .A1(n204), .A2(execution_result_MW_reg[12]), .B1(n2013), 
        .B2(csr_rd_MW_reg[12]), .ZN(n155) );
  AOI22_X1 U313 ( .A1(n2014), .A2(n2192), .B1(n2009), .B2(
        load_data_MW_wire[12]), .ZN(n154) );
  NAND3_X1 U314 ( .A1(n156), .A2(n155), .A3(n154), .ZN(n633) );
  AOI22_X1 U315 ( .A1(n202), .A2(immediate_MW_reg[11]), .B1(n201), .B2(
        address_MW_reg[11]), .ZN(n160) );
  AOI22_X1 U316 ( .A1(n204), .A2(execution_result_MW_reg[11]), .B1(n2013), 
        .B2(csr_rd_MW_reg[11]), .ZN(n159) );
  AOI22_X1 U318 ( .A1(n2014), .A2(n2191), .B1(n2009), .B2(
        load_data_MW_wire[11]), .ZN(n158) );
  NAND3_X1 U319 ( .A1(n160), .A2(n159), .A3(n158), .ZN(n635) );
  AOI22_X1 U320 ( .A1(n202), .A2(immediate_MW_reg[10]), .B1(n201), .B2(
        address_MW_reg[10]), .ZN(n164) );
  AOI22_X1 U321 ( .A1(n204), .A2(execution_result_MW_reg[10]), .B1(n2013), 
        .B2(csr_rd_MW_reg[10]), .ZN(n163) );
  AOI22_X1 U323 ( .A1(n2014), .A2(n2190), .B1(n2009), .B2(
        load_data_MW_wire[10]), .ZN(n162) );
  NAND3_X1 U324 ( .A1(n164), .A2(n163), .A3(n162), .ZN(n637) );
  AOI22_X1 U325 ( .A1(n202), .A2(immediate_MW_reg[9]), .B1(n201), .B2(
        address_MW_reg[9]), .ZN(n168) );
  AOI22_X1 U326 ( .A1(n204), .A2(execution_result_MW_reg[9]), .B1(n2013), .B2(
        csr_rd_MW_reg[9]), .ZN(n167) );
  AOI22_X1 U328 ( .A1(n2014), .A2(n2189), .B1(n2009), .B2(load_data_MW_wire[9]), .ZN(n166) );
  NAND3_X1 U329 ( .A1(n168), .A2(n167), .A3(n166), .ZN(n639) );
  AOI22_X1 U330 ( .A1(n202), .A2(immediate_MW_reg[8]), .B1(n201), .B2(
        address_MW_reg[8]), .ZN(n172) );
  AOI22_X1 U331 ( .A1(n204), .A2(execution_result_MW_reg[8]), .B1(n2013), .B2(
        csr_rd_MW_reg[8]), .ZN(n171) );
  AOI22_X1 U333 ( .A1(n2014), .A2(n2188), .B1(n2009), .B2(load_data_MW_wire[8]), .ZN(n170) );
  NAND3_X1 U334 ( .A1(n172), .A2(n171), .A3(n170), .ZN(n641) );
  AOI22_X1 U335 ( .A1(n202), .A2(immediate_MW_reg[7]), .B1(n201), .B2(
        address_MW_reg[7]), .ZN(n176) );
  AOI22_X1 U336 ( .A1(n204), .A2(execution_result_MW_reg[7]), .B1(n2013), .B2(
        csr_rd_MW_reg[7]), .ZN(n175) );
  AOI22_X1 U338 ( .A1(n2014), .A2(n2187), .B1(n2009), .B2(load_data_MW_wire[7]), .ZN(n174) );
  NAND3_X1 U339 ( .A1(n176), .A2(n175), .A3(n174), .ZN(n643) );
  AOI22_X1 U340 ( .A1(n202), .A2(immediate_MW_reg[6]), .B1(n201), .B2(
        address_MW_reg[6]), .ZN(n180) );
  AOI22_X1 U341 ( .A1(n204), .A2(execution_result_MW_reg[6]), .B1(n2013), .B2(
        csr_rd_MW_reg[6]), .ZN(n179) );
  AOI22_X1 U343 ( .A1(n2014), .A2(n2186), .B1(n2009), .B2(load_data_MW_wire[6]), .ZN(n178) );
  NAND3_X1 U344 ( .A1(n180), .A2(n179), .A3(n178), .ZN(n645) );
  AOI22_X1 U345 ( .A1(n202), .A2(immediate_MW_reg[5]), .B1(n201), .B2(
        address_MW_reg[5]), .ZN(n184) );
  AOI22_X1 U346 ( .A1(n204), .A2(execution_result_MW_reg[5]), .B1(n2013), .B2(
        csr_rd_MW_reg[5]), .ZN(n183) );
  AOI22_X1 U348 ( .A1(n2014), .A2(n2185), .B1(n2009), .B2(load_data_MW_wire[5]), .ZN(n182) );
  NAND3_X1 U349 ( .A1(n184), .A2(n183), .A3(n182), .ZN(n647) );
  AOI22_X1 U350 ( .A1(n202), .A2(immediate_MW_reg[4]), .B1(n201), .B2(
        address_MW_reg[4]), .ZN(n188) );
  AOI22_X1 U351 ( .A1(n204), .A2(execution_result_MW_reg[4]), .B1(n2013), .B2(
        csr_rd_MW_reg[4]), .ZN(n187) );
  AOI22_X1 U353 ( .A1(n2014), .A2(n2184), .B1(n205), .B2(load_data_MW_wire[4]), 
        .ZN(n186) );
  NAND3_X1 U354 ( .A1(n188), .A2(n187), .A3(n186), .ZN(n649) );
  AOI22_X1 U355 ( .A1(n202), .A2(immediate_MW_reg[3]), .B1(n201), .B2(
        address_MW_reg[3]), .ZN(n192) );
  AOI22_X1 U356 ( .A1(n204), .A2(execution_result_MW_reg[3]), .B1(n2013), .B2(
        csr_rd_MW_reg[3]), .ZN(n191) );
  AOI22_X1 U358 ( .A1(n2014), .A2(n2183), .B1(n205), .B2(load_data_MW_wire[3]), 
        .ZN(n190) );
  NAND3_X1 U359 ( .A1(n192), .A2(n191), .A3(n190), .ZN(n651) );
  AOI22_X1 U360 ( .A1(n202), .A2(immediate_MW_reg[2]), .B1(n201), .B2(
        address_MW_reg[2]), .ZN(n196) );
  AOI22_X1 U361 ( .A1(n204), .A2(execution_result_MW_reg[2]), .B1(n2013), .B2(
        csr_rd_MW_reg[2]), .ZN(n195) );
  AOI22_X1 U363 ( .A1(n2014), .A2(n2182), .B1(n2009), .B2(load_data_MW_wire[2]), .ZN(n194) );
  NAND3_X1 U364 ( .A1(n196), .A2(n195), .A3(n194), .ZN(n653) );
  AOI22_X1 U365 ( .A1(n202), .A2(immediate_MW_reg[1]), .B1(n201), .B2(
        address_MW_reg[1]), .ZN(n200) );
  AOI22_X1 U366 ( .A1(n204), .A2(execution_result_MW_reg[1]), .B1(n2013), .B2(
        csr_rd_MW_reg[1]), .ZN(n199) );
  AOI22_X1 U368 ( .A1(n2014), .A2(n2181), .B1(n205), .B2(load_data_MW_wire[1]), 
        .ZN(n198) );
  NAND3_X1 U369 ( .A1(n200), .A2(n199), .A3(n198), .ZN(n655) );
  AOI22_X1 U370 ( .A1(n202), .A2(immediate_MW_reg[0]), .B1(n201), .B2(
        address_MW_reg[0]), .ZN(n210) );
  AOI22_X1 U371 ( .A1(n204), .A2(execution_result_MW_reg[0]), .B1(n2013), .B2(
        csr_rd_MW_reg[0]), .ZN(n209) );
  AOI22_X1 U373 ( .A1(n2014), .A2(n2180), .B1(n205), .B2(load_data_MW_wire[0]), 
        .ZN(n208) );
  NAND3_X1 U374 ( .A1(n210), .A2(n209), .A3(n208), .ZN(n657) );
  AOI22_X1 U424 ( .A1(n1833), .A2(n2445), .B1(n1206), .B2(n2443), .ZN(n1581)
         );
  AOI22_X1 U425 ( .A1(n2445), .A2(n2061), .B1(n1205), .B2(n2437), .ZN(n1582)
         );
  AOI22_X1 U427 ( .A1(n2446), .A2(n1218), .B1(n1203), .B2(n2442), .ZN(n1584)
         );
  AOI22_X1 U428 ( .A1(n2444), .A2(n1219), .B1(n1202), .B2(n2438), .ZN(n1585)
         );
  AOI22_X1 U429 ( .A1(n2447), .A2(n1220), .B1(n1201), .B2(n2441), .ZN(n1586)
         );
  AOI22_X1 U430 ( .A1(n2446), .A2(n2068), .B1(n1200), .B2(n2438), .ZN(n1587)
         );
  AOI22_X1 U431 ( .A1(n2446), .A2(n1222), .B1(n1199), .B2(n2440), .ZN(n1588)
         );
  AOI22_X1 U432 ( .A1(n2444), .A2(n1223), .B1(n1198), .B2(n2438), .ZN(n1589)
         );
  AOI22_X1 U434 ( .A1(n2444), .A2(n1912), .B1(n1196), .B2(n2439), .ZN(n1591)
         );
  AOI22_X1 U435 ( .A1(n2446), .A2(n1911), .B1(n1195), .B2(n2440), .ZN(n1592)
         );
  AOI22_X1 U436 ( .A1(n2446), .A2(n2069), .B1(n1194), .B2(n2443), .ZN(n1593)
         );
  AOI22_X1 U437 ( .A1(n2444), .A2(n1913), .B1(n1193), .B2(n2443), .ZN(n1594)
         );
  AOI22_X1 U438 ( .A1(n2447), .A2(n2057), .B1(n1192), .B2(n2443), .ZN(n1595)
         );
  AOI22_X1 U439 ( .A1(n2446), .A2(n2060), .B1(n1191), .B2(n2443), .ZN(n1596)
         );
  AOI22_X1 U440 ( .A1(n2445), .A2(n1231), .B1(n1190), .B2(n2443), .ZN(n1597)
         );
  AOI22_X1 U441 ( .A1(n2444), .A2(n1232), .B1(n1189), .B2(n2443), .ZN(n1598)
         );
  AOI22_X1 U442 ( .A1(n2445), .A2(n2071), .B1(n1188), .B2(n2443), .ZN(n1599)
         );
  AOI22_X1 U443 ( .A1(n2446), .A2(n2075), .B1(n1187), .B2(n2443), .ZN(n1600)
         );
  AOI22_X1 U444 ( .A1(n2446), .A2(n1831), .B1(n1186), .B2(n2443), .ZN(n1601)
         );
  AOI22_X1 U449 ( .A1(n2447), .A2(n2070), .B1(n1181), .B2(n2441), .ZN(n1606)
         );
  AOI22_X1 U450 ( .A1(n2444), .A2(n2052), .B1(n1180), .B2(n2442), .ZN(n1607)
         );
  AOI22_X1 U451 ( .A1(n2446), .A2(n2074), .B1(n1179), .B2(n2437), .ZN(n1608)
         );
  AOI22_X1 U453 ( .A1(n2446), .A2(n1244), .B1(n1177), .B2(n2442), .ZN(n1610)
         );
  AOI22_X1 U454 ( .A1(n2446), .A2(n2073), .B1(n1176), .B2(n2438), .ZN(n1611)
         );
  MUX2_X1 U455 ( .A(pc_EX_reg[31]), .B(pc_FD_reg[31]), .S(n2151), .Z(n1612) );
  MUX2_X1 U458 ( .A(pc_EX_reg[30]), .B(pc_FD_reg[30]), .S(n2461), .Z(n1614) );
  MUX2_X1 U461 ( .A(pc_EX_reg[29]), .B(pc_FD_reg[29]), .S(n2465), .Z(n1616) );
  MUX2_X1 U464 ( .A(pc_EX_reg[28]), .B(pc_FD_reg[28]), .S(n2462), .Z(n1618) );
  MUX2_X1 U467 ( .A(pc_EX_reg[27]), .B(pc_FD_reg[27]), .S(n2466), .Z(n1620) );
  MUX2_X1 U470 ( .A(pc_EX_reg[26]), .B(pc_FD_reg[26]), .S(n2463), .Z(n1622) );
  MUX2_X1 U473 ( .A(pc_EX_reg[25]), .B(pc_FD_reg[25]), .S(n2151), .Z(n1624) );
  MUX2_X1 U476 ( .A(pc_EX_reg[24]), .B(pc_FD_reg[24]), .S(n2465), .Z(n1626) );
  MUX2_X1 U479 ( .A(pc_EX_reg[23]), .B(pc_FD_reg[23]), .S(n2462), .Z(n1628) );
  MUX2_X1 U482 ( .A(pc_EX_reg[22]), .B(pc_FD_reg[22]), .S(n2465), .Z(n1630) );
  MUX2_X1 U485 ( .A(pc_EX_reg[21]), .B(pc_FD_reg[21]), .S(n2467), .Z(n1632) );
  MUX2_X1 U488 ( .A(pc_EX_reg[20]), .B(pc_FD_reg[20]), .S(n2463), .Z(n1634) );
  MUX2_X1 U491 ( .A(pc_EX_reg[19]), .B(pc_FD_reg[19]), .S(n2462), .Z(n1636) );
  MUX2_X1 U494 ( .A(pc_EX_reg[18]), .B(pc_FD_reg[18]), .S(n2464), .Z(n1638) );
  MUX2_X1 U497 ( .A(pc_EX_reg[17]), .B(pc_FD_reg[17]), .S(n2463), .Z(n1640) );
  MUX2_X1 U500 ( .A(pc_EX_reg[16]), .B(pc_FD_reg[16]), .S(n2466), .Z(n1642) );
  MUX2_X1 U503 ( .A(pc_EX_reg[15]), .B(pc_FD_reg[15]), .S(n2462), .Z(n1644) );
  MUX2_X1 U506 ( .A(pc_EX_reg[14]), .B(pc_FD_reg[14]), .S(n2151), .Z(n1646) );
  MUX2_X1 U509 ( .A(pc_EX_reg[13]), .B(pc_FD_reg[13]), .S(n2462), .Z(n1648) );
  MUX2_X1 U512 ( .A(pc_EX_reg[12]), .B(pc_FD_reg[12]), .S(n2466), .Z(n1650) );
  MUX2_X1 U515 ( .A(pc_EX_reg[11]), .B(pc_FD_reg[11]), .S(n2464), .Z(n1652) );
  MUX2_X1 U518 ( .A(pc_EX_reg[10]), .B(pc_FD_reg[10]), .S(n2151), .Z(n1654) );
  MUX2_X1 U521 ( .A(pc_EX_reg[9]), .B(pc_FD_reg[9]), .S(n2464), .Z(n1656) );
  MUX2_X1 U524 ( .A(pc_EX_reg[8]), .B(pc_FD_reg[8]), .S(n2464), .Z(n1658) );
  MUX2_X1 U527 ( .A(pc_EX_reg[7]), .B(pc_FD_reg[7]), .S(n2467), .Z(n1660) );
  OAI21_X1 U528 ( .B1(n1247), .B2(n1131), .A(n1274), .ZN(n1661) );
  AOI22_X1 U529 ( .A1(n2006), .A2(address_EX_wire[7]), .B1(n2498), .B2(
        pc_FD_reg[7]), .ZN(n1274) );
  MUX2_X1 U530 ( .A(pc_EX_reg[6]), .B(pc_FD_reg[6]), .S(n2463), .Z(n1662) );
  OAI21_X1 U531 ( .B1(n1247), .B2(n1130), .A(n1275), .ZN(n1663) );
  AOI22_X1 U532 ( .A1(n2006), .A2(address_EX_wire[6]), .B1(n2498), .B2(
        pc_FD_reg[6]), .ZN(n1275) );
  MUX2_X1 U533 ( .A(pc_EX_reg[5]), .B(pc_FD_reg[5]), .S(n2152), .Z(n1664) );
  OAI21_X1 U534 ( .B1(n1247), .B2(n1129), .A(n1276), .ZN(n1665) );
  AOI22_X1 U535 ( .A1(n2006), .A2(address_EX_wire[5]), .B1(n2498), .B2(
        pc_FD_reg[5]), .ZN(n1276) );
  MUX2_X1 U536 ( .A(pc_EX_reg[4]), .B(pc_FD_reg[4]), .S(n2457), .Z(n1666) );
  OAI21_X1 U537 ( .B1(n1247), .B2(n1128), .A(n1277), .ZN(n1667) );
  AOI22_X1 U538 ( .A1(n2006), .A2(address_EX_wire[4]), .B1(n2498), .B2(
        pc_FD_reg[4]), .ZN(n1277) );
  MUX2_X1 U539 ( .A(pc_EX_reg[3]), .B(pc_FD_reg[3]), .S(n2458), .Z(n1668) );
  OAI21_X1 U540 ( .B1(n1247), .B2(n1127), .A(n1278), .ZN(n1669) );
  AOI22_X1 U541 ( .A1(n2006), .A2(address_EX_wire[3]), .B1(n2498), .B2(
        pc_FD_reg[3]), .ZN(n1278) );
  MUX2_X1 U542 ( .A(pc_EX_reg[2]), .B(pc_FD_reg[2]), .S(n2153), .Z(n1670) );
  OAI21_X1 U543 ( .B1(n1247), .B2(n1126), .A(n1279), .ZN(n1671) );
  AOI22_X1 U544 ( .A1(n2006), .A2(address_EX_wire[2]), .B1(n2498), .B2(
        pc_FD_reg[2]), .ZN(n1279) );
  MUX2_X1 U545 ( .A(pc_EX_reg[1]), .B(pc_FD_reg[1]), .S(n2153), .Z(n1672) );
  OAI21_X1 U546 ( .B1(n1247), .B2(n1125), .A(n1280), .ZN(n1673) );
  AOI22_X1 U547 ( .A1(n2006), .A2(address_EX_wire[1]), .B1(n2498), .B2(
        pc_FD_reg[1]), .ZN(n1280) );
  MUX2_X1 U548 ( .A(pc_EX_reg[0]), .B(pc_FD_reg[0]), .S(n2458), .Z(n1674) );
  OAI21_X1 U549 ( .B1(n1247), .B2(n1124), .A(n1281), .ZN(n1675) );
  AOI22_X1 U550 ( .A1(n2006), .A2(address_EX_wire[0]), .B1(n2498), .B2(
        pc_FD_reg[0]), .ZN(n1281) );
  MUX2_X1 U554 ( .A(next_pc_EX_reg[31]), .B(next_pc_FD_wire[31]), .S(n2458), 
        .Z(n1676) );
  MUX2_X1 U555 ( .A(next_pc_EX_reg[30]), .B(next_pc_FD_wire[30]), .S(n2457), 
        .Z(n1677) );
  MUX2_X1 U556 ( .A(next_pc_EX_reg[29]), .B(next_pc_FD_wire[29]), .S(n2457), 
        .Z(n1678) );
  MUX2_X1 U557 ( .A(next_pc_EX_reg[28]), .B(next_pc_FD_wire[28]), .S(n2460), 
        .Z(n1679) );
  MUX2_X1 U558 ( .A(next_pc_EX_reg[27]), .B(next_pc_FD_wire[27]), .S(n2460), 
        .Z(n1680) );
  MUX2_X1 U559 ( .A(next_pc_EX_reg[26]), .B(next_pc_FD_wire[26]), .S(n2152), 
        .Z(n1681) );
  MUX2_X1 U560 ( .A(next_pc_EX_reg[25]), .B(next_pc_FD_wire[25]), .S(n2457), 
        .Z(n1682) );
  MUX2_X1 U561 ( .A(next_pc_EX_reg[24]), .B(next_pc_FD_wire[24]), .S(n2461), 
        .Z(n1683) );
  MUX2_X1 U562 ( .A(next_pc_EX_reg[23]), .B(next_pc_FD_wire[23]), .S(n2457), 
        .Z(n1684) );
  MUX2_X1 U563 ( .A(next_pc_EX_reg[22]), .B(next_pc_FD_wire[22]), .S(n2458), 
        .Z(n1685) );
  MUX2_X1 U564 ( .A(next_pc_EX_reg[21]), .B(next_pc_FD_wire[21]), .S(n2458), 
        .Z(n1686) );
  MUX2_X1 U565 ( .A(next_pc_EX_reg[20]), .B(next_pc_FD_wire[20]), .S(n2459), 
        .Z(n1687) );
  MUX2_X1 U566 ( .A(next_pc_EX_reg[19]), .B(next_pc_FD_wire[19]), .S(n2461), 
        .Z(n1688) );
  MUX2_X1 U567 ( .A(next_pc_EX_reg[18]), .B(next_pc_FD_wire[18]), .S(n2152), 
        .Z(n1689) );
  MUX2_X1 U568 ( .A(next_pc_EX_reg[17]), .B(next_pc_FD_wire[17]), .S(n2153), 
        .Z(n1690) );
  MUX2_X1 U569 ( .A(next_pc_EX_reg[16]), .B(next_pc_FD_wire[16]), .S(n2457), 
        .Z(n1691) );
  MUX2_X1 U570 ( .A(next_pc_EX_reg[15]), .B(next_pc_FD_wire[15]), .S(n2458), 
        .Z(n1692) );
  MUX2_X1 U571 ( .A(next_pc_EX_reg[14]), .B(next_pc_FD_wire[14]), .S(n2460), 
        .Z(n1693) );
  MUX2_X1 U572 ( .A(next_pc_EX_reg[13]), .B(next_pc_FD_wire[13]), .S(n2459), 
        .Z(n1694) );
  MUX2_X1 U573 ( .A(next_pc_EX_reg[12]), .B(next_pc_FD_wire[12]), .S(n2461), 
        .Z(n1695) );
  MUX2_X1 U574 ( .A(next_pc_EX_reg[11]), .B(next_pc_FD_wire[11]), .S(n2152), 
        .Z(n1696) );
  MUX2_X1 U575 ( .A(next_pc_EX_reg[10]), .B(next_pc_FD_wire[10]), .S(n2457), 
        .Z(n1697) );
  MUX2_X1 U576 ( .A(next_pc_EX_reg[9]), .B(next_pc_FD_wire[9]), .S(n2458), .Z(
        n1698) );
  MUX2_X1 U577 ( .A(next_pc_EX_reg[8]), .B(next_pc_FD_wire[8]), .S(n2460), .Z(
        n1699) );
  MUX2_X1 U578 ( .A(next_pc_EX_reg[7]), .B(next_pc_FD_wire[7]), .S(n2459), .Z(
        n1700) );
  MUX2_X1 U579 ( .A(next_pc_EX_reg[6]), .B(next_pc_FD_wire[6]), .S(n2461), .Z(
        n1701) );
  MUX2_X1 U580 ( .A(next_pc_EX_reg[5]), .B(next_pc_FD_wire[5]), .S(n2152), .Z(
        n1702) );
  MUX2_X1 U581 ( .A(next_pc_EX_reg[4]), .B(next_pc_FD_wire[4]), .S(n2153), .Z(
        n1703) );
  MUX2_X1 U582 ( .A(next_pc_EX_reg[3]), .B(next_pc_FD_wire[3]), .S(n2457), .Z(
        n1704) );
  MUX2_X1 U583 ( .A(next_pc_EX_reg[2]), .B(next_pc_FD_wire[2]), .S(n2458), .Z(
        n1705) );
  MUX2_X1 U584 ( .A(next_pc_EX_reg[1]), .B(next_pc_FD_wire[1]), .S(n2460), .Z(
        n1706) );
  MUX2_X1 U585 ( .A(next_pc_EX_reg[0]), .B(next_pc_FD_wire[0]), .S(n2459), .Z(
        n1707) );
  AOI22_X1 U586 ( .A1(n2462), .A2(instruction_type_FD_wire[2]), .B1(n2007), 
        .B2(instruction_type_EX_reg[2]), .ZN(n1282) );
  AOI22_X1 U587 ( .A1(n2467), .A2(instruction_type_FD_wire[1]), .B1(n2007), 
        .B2(instruction_type_EX_reg[1]), .ZN(n1284) );
  AOI22_X1 U590 ( .A1(n2151), .A2(immediate_FD_wire[31]), .B1(n2007), .B2(
        immediate_EX_reg[31]), .ZN(n1287) );
  AOI22_X1 U591 ( .A1(n2465), .A2(immediate_FD_wire[30]), .B1(n2007), .B2(
        immediate_EX_reg[30]), .ZN(n1288) );
  AOI22_X1 U592 ( .A1(n2464), .A2(immediate_FD_wire[29]), .B1(n2007), .B2(
        immediate_EX_reg[29]), .ZN(n1289) );
  AOI22_X1 U593 ( .A1(n2465), .A2(immediate_FD_wire[28]), .B1(n2007), .B2(
        immediate_EX_reg[28]), .ZN(n1290) );
  AOI22_X1 U594 ( .A1(n2466), .A2(immediate_FD_wire[27]), .B1(n2007), .B2(
        immediate_EX_reg[27]), .ZN(n1291) );
  AOI22_X1 U595 ( .A1(n2151), .A2(immediate_FD_wire[26]), .B1(n2007), .B2(
        immediate_EX_reg[26]), .ZN(n1292) );
  AOI22_X1 U596 ( .A1(n2466), .A2(immediate_FD_wire[25]), .B1(n2007), .B2(
        immediate_EX_reg[25]), .ZN(n1293) );
  AOI22_X1 U597 ( .A1(n2463), .A2(immediate_FD_wire[24]), .B1(n2434), .B2(
        immediate_EX_reg[24]), .ZN(n1294) );
  AOI22_X1 U598 ( .A1(n2462), .A2(immediate_FD_wire[23]), .B1(n2434), .B2(
        immediate_EX_reg[23]), .ZN(n1295) );
  AOI22_X1 U599 ( .A1(n2466), .A2(immediate_FD_wire[22]), .B1(n2434), .B2(
        immediate_EX_reg[22]), .ZN(n1296) );
  AOI22_X1 U600 ( .A1(n2464), .A2(immediate_FD_wire[21]), .B1(n2434), .B2(
        immediate_EX_reg[21]), .ZN(n1297) );
  AOI22_X1 U601 ( .A1(n2465), .A2(immediate_FD_wire[20]), .B1(n2434), .B2(
        immediate_EX_reg[20]), .ZN(n1298) );
  AOI22_X1 U602 ( .A1(n2465), .A2(immediate_FD_wire[19]), .B1(n2434), .B2(
        immediate_EX_reg[19]), .ZN(n1299) );
  AOI22_X1 U603 ( .A1(n2151), .A2(immediate_FD_wire[18]), .B1(n2434), .B2(
        immediate_EX_reg[18]), .ZN(n1300) );
  AOI22_X1 U604 ( .A1(n2463), .A2(immediate_FD_wire[17]), .B1(n2434), .B2(
        immediate_EX_reg[17]), .ZN(n1301) );
  AOI22_X1 U605 ( .A1(n2467), .A2(immediate_FD_wire[16]), .B1(n2434), .B2(
        immediate_EX_reg[16]), .ZN(n1302) );
  AOI22_X1 U606 ( .A1(n2463), .A2(immediate_FD_wire[15]), .B1(n2434), .B2(
        immediate_EX_reg[15]), .ZN(n1303) );
  AOI22_X1 U607 ( .A1(n2463), .A2(immediate_FD_wire[14]), .B1(n2434), .B2(
        immediate_EX_reg[14]), .ZN(n1304) );
  AOI22_X1 U608 ( .A1(n2462), .A2(immediate_FD_wire[13]), .B1(n2434), .B2(
        immediate_EX_reg[13]), .ZN(n1305) );
  AOI22_X1 U609 ( .A1(n2462), .A2(immediate_FD_wire[12]), .B1(n2434), .B2(
        immediate_EX_reg[12]), .ZN(n1306) );
  AOI22_X1 U610 ( .A1(n2467), .A2(immediate_FD_wire[11]), .B1(n2434), .B2(
        immediate_EX_reg[11]), .ZN(n1307) );
  AOI22_X1 U611 ( .A1(n2463), .A2(immediate_FD_wire[10]), .B1(n2434), .B2(
        immediate_EX_reg[10]), .ZN(n1308) );
  AOI22_X1 U612 ( .A1(n2151), .A2(immediate_FD_wire[9]), .B1(n2434), .B2(
        immediate_EX_reg[9]), .ZN(n1309) );
  AOI22_X1 U613 ( .A1(n2464), .A2(immediate_FD_wire[8]), .B1(n2434), .B2(
        immediate_EX_reg[8]), .ZN(n1310) );
  AOI22_X1 U614 ( .A1(n2464), .A2(immediate_FD_wire[7]), .B1(n2434), .B2(
        immediate_EX_reg[7]), .ZN(n1311) );
  AOI22_X1 U615 ( .A1(n2464), .A2(immediate_FD_wire[6]), .B1(n2434), .B2(
        immediate_EX_reg[6]), .ZN(n1312) );
  AOI22_X1 U616 ( .A1(n2462), .A2(immediate_FD_wire[5]), .B1(n2434), .B2(
        immediate_EX_reg[5]), .ZN(n1313) );
  AOI22_X1 U617 ( .A1(n2467), .A2(immediate_FD_wire[4]), .B1(n2433), .B2(
        immediate_EX_reg[4]), .ZN(n1314) );
  AOI22_X1 U618 ( .A1(n2466), .A2(immediate_FD_wire[3]), .B1(n2433), .B2(
        immediate_EX_reg[3]), .ZN(n1315) );
  AOI22_X1 U619 ( .A1(n2468), .A2(immediate_FD_wire[2]), .B1(n2433), .B2(
        immediate_EX_reg[2]), .ZN(n1316) );
  AOI22_X1 U620 ( .A1(n2468), .A2(immediate_FD_wire[1]), .B1(n2433), .B2(
        immediate_EX_reg[1]), .ZN(n1317) );
  AOI22_X1 U621 ( .A1(n2468), .A2(immediate_FD_wire[0]), .B1(n2433), .B2(
        immediate_EX_reg[0]), .ZN(n1318) );
  MUX2_X1 U622 ( .A(csr_data_EX_reg[31]), .B(csr_data_FD_wire[31]), .S(n2461), 
        .Z(n1709) );
  MUX2_X1 U623 ( .A(csr_data_EX_reg[30]), .B(csr_data_FD_wire[30]), .S(n2459), 
        .Z(n1710) );
  MUX2_X1 U624 ( .A(csr_data_EX_reg[29]), .B(csr_data_FD_wire[29]), .S(n2460), 
        .Z(n1711) );
  MUX2_X1 U625 ( .A(csr_data_EX_reg[28]), .B(csr_data_FD_wire[28]), .S(n2458), 
        .Z(n1712) );
  MUX2_X1 U626 ( .A(csr_data_EX_reg[27]), .B(csr_data_FD_wire[27]), .S(n2457), 
        .Z(n1713) );
  MUX2_X1 U627 ( .A(csr_data_EX_reg[26]), .B(csr_data_FD_wire[26]), .S(n2152), 
        .Z(n1714) );
  MUX2_X1 U628 ( .A(csr_data_EX_reg[25]), .B(csr_data_FD_wire[25]), .S(n2461), 
        .Z(n1715) );
  MUX2_X1 U629 ( .A(csr_data_EX_reg[24]), .B(csr_data_FD_wire[24]), .S(n2459), 
        .Z(n1716) );
  MUX2_X1 U630 ( .A(csr_data_EX_reg[23]), .B(csr_data_FD_wire[23]), .S(n2457), 
        .Z(n1717) );
  MUX2_X1 U631 ( .A(csr_data_EX_reg[22]), .B(csr_data_FD_wire[22]), .S(n2152), 
        .Z(n1718) );
  MUX2_X1 U632 ( .A(csr_data_EX_reg[21]), .B(csr_data_FD_wire[21]), .S(n2152), 
        .Z(n1719) );
  MUX2_X1 U633 ( .A(csr_data_EX_reg[20]), .B(csr_data_FD_wire[20]), .S(n2152), 
        .Z(n1720) );
  MUX2_X1 U634 ( .A(csr_data_EX_reg[19]), .B(csr_data_FD_wire[19]), .S(n2461), 
        .Z(n1721) );
  MUX2_X1 U635 ( .A(csr_data_EX_reg[18]), .B(csr_data_FD_wire[18]), .S(n2461), 
        .Z(n1722) );
  MUX2_X1 U636 ( .A(csr_data_EX_reg[17]), .B(csr_data_FD_wire[17]), .S(n2461), 
        .Z(n1723) );
  MUX2_X1 U637 ( .A(csr_data_EX_reg[16]), .B(csr_data_FD_wire[16]), .S(n2459), 
        .Z(n1724) );
  MUX2_X1 U638 ( .A(csr_data_EX_reg[15]), .B(csr_data_FD_wire[15]), .S(n2459), 
        .Z(n1725) );
  MUX2_X1 U639 ( .A(csr_data_EX_reg[14]), .B(csr_data_FD_wire[14]), .S(n2459), 
        .Z(n1726) );
  MUX2_X1 U640 ( .A(csr_data_EX_reg[13]), .B(csr_data_FD_wire[13]), .S(n2460), 
        .Z(n1727) );
  MUX2_X1 U641 ( .A(csr_data_EX_reg[12]), .B(csr_data_FD_wire[12]), .S(n2460), 
        .Z(n1728) );
  MUX2_X1 U642 ( .A(csr_data_EX_reg[11]), .B(csr_data_FD_wire[11]), .S(n2153), 
        .Z(n1729) );
  MUX2_X1 U643 ( .A(csr_data_EX_reg[10]), .B(csr_data_FD_wire[10]), .S(n2152), 
        .Z(n1730) );
  MUX2_X1 U644 ( .A(csr_data_EX_reg[9]), .B(csr_data_FD_wire[9]), .S(n2461), 
        .Z(n1731) );
  MUX2_X1 U645 ( .A(csr_data_EX_reg[8]), .B(csr_data_FD_wire[8]), .S(n2459), 
        .Z(n1732) );
  MUX2_X1 U646 ( .A(csr_data_EX_reg[7]), .B(csr_data_FD_wire[7]), .S(n2460), 
        .Z(n1733) );
  MUX2_X1 U647 ( .A(csr_data_EX_reg[6]), .B(csr_data_FD_wire[6]), .S(n2458), 
        .Z(n1734) );
  MUX2_X1 U648 ( .A(csr_data_EX_reg[5]), .B(csr_data_FD_wire[5]), .S(n2457), 
        .Z(n1735) );
  MUX2_X1 U649 ( .A(csr_data_EX_reg[4]), .B(csr_data_FD_wire[4]), .S(n2153), 
        .Z(n1736) );
  MUX2_X1 U650 ( .A(csr_data_EX_reg[3]), .B(csr_data_FD_wire[3]), .S(n2152), 
        .Z(n1737) );
  MUX2_X1 U651 ( .A(csr_data_EX_reg[2]), .B(csr_data_FD_wire[2]), .S(n2459), 
        .Z(n1738) );
  MUX2_X1 U652 ( .A(csr_data_EX_reg[1]), .B(csr_data_FD_wire[1]), .S(n2460), 
        .Z(n1739) );
  MUX2_X1 U653 ( .A(csr_data_EX_reg[0]), .B(csr_data_FD_wire[0]), .S(n2458), 
        .Z(n1740) );
  AOI22_X1 U654 ( .A1(n2154), .A2(n2428), .B1(n2470), .B2(opcode_FD_wire[6]), 
        .ZN(n1319) );
  AOI22_X1 U655 ( .A1(n2414), .A2(n2428), .B1(n2470), .B2(opcode_FD_wire[5]), 
        .ZN(n1320) );
  OAI21_X1 U656 ( .B1(n2470), .B2(n1167), .A(n1321), .ZN(n1741) );
  AOI21_X1 U657 ( .B1(opcode_FD_wire[4]), .B2(n2469), .A(n2454), .ZN(n1321) );
  AOI22_X1 U659 ( .A1(n2072), .A2(n2428), .B1(n2470), .B2(opcode_FD_wire[2]), 
        .ZN(n1323) );
  NAND2_X1 U662 ( .A1(n2005), .A2(n1325), .ZN(n1743) );
  AOI22_X1 U663 ( .A1(opcode_EX_reg[0]), .A2(n2428), .B1(n2470), .B2(
        opcode_FD_wire[0]), .ZN(n1325) );
  AOI22_X1 U664 ( .A1(n2468), .A2(funct3_FD_wire[2]), .B1(n2433), .B2(
        funct3_EX_reg[2]), .ZN(n1326) );
  AOI22_X1 U665 ( .A1(n2468), .A2(funct3_FD_wire[1]), .B1(n2433), .B2(n2474), 
        .ZN(n1327) );
  AOI22_X1 U666 ( .A1(n2468), .A2(funct3_FD_wire[0]), .B1(n2433), .B2(
        funct3_EX_reg[0]), .ZN(n1328) );
  AOI22_X1 U667 ( .A1(n2468), .A2(funct7_FD_wire[6]), .B1(n2433), .B2(
        funct7_EX_reg[6]), .ZN(n1329) );
  AOI22_X1 U668 ( .A1(n2468), .A2(funct7_FD_wire[5]), .B1(n2433), .B2(
        funct7_EX_reg[5]), .ZN(n1330) );
  AOI22_X1 U669 ( .A1(n2468), .A2(funct7_FD_wire[4]), .B1(n2433), .B2(
        funct7_EX_reg[4]), .ZN(n1331) );
  AOI22_X1 U670 ( .A1(n2469), .A2(funct7_FD_wire[3]), .B1(n2433), .B2(
        funct7_EX_reg[3]), .ZN(n1332) );
  AOI22_X1 U671 ( .A1(n2468), .A2(funct7_FD_wire[2]), .B1(n2433), .B2(
        funct7_EX_reg[2]), .ZN(n1333) );
  AOI22_X1 U672 ( .A1(n2469), .A2(funct7_FD_wire[1]), .B1(n2433), .B2(
        funct7_EX_reg[1]), .ZN(n1334) );
  AOI22_X1 U673 ( .A1(n2468), .A2(funct7_FD_wire[0]), .B1(n2433), .B2(
        funct7_EX_reg[0]), .ZN(n1335) );
  AOI22_X1 U674 ( .A1(n2469), .A2(funct12_FD_wire[11]), .B1(n2433), .B2(
        funct12_EX_reg[11]), .ZN(n1336) );
  AOI22_X1 U675 ( .A1(n2469), .A2(funct12_FD_wire[10]), .B1(n2433), .B2(
        funct12_EX_reg[10]), .ZN(n1337) );
  AOI22_X1 U676 ( .A1(n2468), .A2(funct12_FD_wire[9]), .B1(n2433), .B2(
        funct12_EX_reg[9]), .ZN(n1338) );
  AOI22_X1 U677 ( .A1(n2469), .A2(funct12_FD_wire[8]), .B1(n2433), .B2(
        funct12_EX_reg[8]), .ZN(n1339) );
  AOI22_X1 U678 ( .A1(n2469), .A2(funct12_FD_wire[7]), .B1(n2433), .B2(
        funct12_EX_reg[7]), .ZN(n1340) );
  AOI22_X1 U679 ( .A1(n2469), .A2(funct12_FD_wire[6]), .B1(n2432), .B2(
        funct12_EX_reg[6]), .ZN(n1341) );
  AOI22_X1 U680 ( .A1(n2469), .A2(funct12_FD_wire[5]), .B1(n2432), .B2(
        funct12_EX_reg[5]), .ZN(n1342) );
  AOI22_X1 U681 ( .A1(n2468), .A2(funct12_FD_wire[4]), .B1(n2432), .B2(
        funct12_EX_reg[4]), .ZN(n1343) );
  AOI22_X1 U682 ( .A1(n2469), .A2(funct12_FD_wire[3]), .B1(n2432), .B2(
        funct12_EX_reg[3]), .ZN(n1344) );
  AOI22_X1 U683 ( .A1(n2469), .A2(funct12_FD_wire[2]), .B1(n2432), .B2(
        funct12_EX_reg[2]), .ZN(n1345) );
  AOI22_X1 U684 ( .A1(n2469), .A2(funct12_FD_wire[1]), .B1(n2432), .B2(
        funct12_EX_reg[1]), .ZN(n1346) );
  AOI22_X1 U685 ( .A1(n2469), .A2(funct12_FD_wire[0]), .B1(n2432), .B2(
        funct12_EX_reg[0]), .ZN(n1347) );
  MUX2_X1 U686 ( .A(read_index_1_EX_reg[4]), .B(read_index_1_FD_wire[4]), .S(
        n2465), .Z(n1744) );
  MUX2_X1 U687 ( .A(read_index_1_EX_reg[3]), .B(read_index_1_FD_wire[3]), .S(
        n2151), .Z(n1745) );
  MUX2_X1 U688 ( .A(read_index_1_EX_reg[2]), .B(read_index_1_FD_wire[2]), .S(
        n2151), .Z(n1746) );
  MUX2_X1 U689 ( .A(read_index_1_EX_reg[1]), .B(read_index_1_FD_wire[1]), .S(
        n2463), .Z(n1747) );
  MUX2_X1 U690 ( .A(read_index_1_EX_reg[0]), .B(read_index_1_FD_wire[0]), .S(
        n2467), .Z(n1748) );
  AOI22_X1 U691 ( .A1(write_index_EX_reg[4]), .A2(n2428), .B1(n2470), .B2(
        write_index_FD_wire[4]), .ZN(n1348) );
  AOI22_X1 U692 ( .A1(write_index_EX_reg[3]), .A2(n2428), .B1(n2470), .B2(
        write_index_FD_wire[3]), .ZN(n1349) );
  AOI22_X1 U693 ( .A1(write_index_EX_reg[2]), .A2(n2428), .B1(n2470), .B2(
        write_index_FD_wire[2]), .ZN(n1350) );
  AOI22_X1 U694 ( .A1(write_index_EX_reg[1]), .A2(n2428), .B1(n2470), .B2(
        write_index_FD_wire[1]), .ZN(n1351) );
  AOI22_X1 U695 ( .A1(write_index_EX_reg[0]), .A2(n2428), .B1(n2470), .B2(
        write_index_FD_wire[0]), .ZN(n1352) );
  MUX2_X1 U696 ( .A(csr_index_EX_reg[11]), .B(csr_index_FD_wire[11]), .S(n2466), .Z(n1749) );
  MUX2_X1 U697 ( .A(csr_index_EX_reg[10]), .B(csr_index_FD_wire[10]), .S(n2467), .Z(n1750) );
  MUX2_X1 U698 ( .A(csr_index_EX_reg[9]), .B(csr_index_FD_wire[9]), .S(n2465), 
        .Z(n1751) );
  MUX2_X1 U699 ( .A(csr_index_EX_reg[8]), .B(csr_index_FD_wire[8]), .S(n2464), 
        .Z(n1752) );
  MUX2_X1 U700 ( .A(csr_index_EX_reg[7]), .B(csr_index_FD_wire[7]), .S(n2466), 
        .Z(n1753) );
  MUX2_X1 U701 ( .A(csr_index_EX_reg[6]), .B(csr_index_FD_wire[6]), .S(n2467), 
        .Z(n1754) );
  MUX2_X1 U702 ( .A(csr_index_EX_reg[5]), .B(csr_index_FD_wire[5]), .S(n2467), 
        .Z(n1755) );
  MUX2_X1 U703 ( .A(csr_index_EX_reg[4]), .B(csr_index_FD_wire[4]), .S(n2464), 
        .Z(n1756) );
  MUX2_X1 U704 ( .A(csr_index_EX_reg[3]), .B(csr_index_FD_wire[3]), .S(n2462), 
        .Z(n1757) );
  MUX2_X1 U705 ( .A(csr_index_EX_reg[2]), .B(csr_index_FD_wire[2]), .S(n2463), 
        .Z(n1758) );
  MUX2_X1 U706 ( .A(csr_index_EX_reg[1]), .B(csr_index_FD_wire[1]), .S(n2151), 
        .Z(n1759) );
  MUX2_X1 U708 ( .A(write_enable_csr_EX_reg), .B(write_enable_csr_FD_wire), 
        .S(n2465), .Z(n1761) );
  AOI22_X1 U709 ( .A1(write_enable_EX_reg), .A2(n2428), .B1(n2470), .B2(
        write_enable_FD_wire), .ZN(n1353) );
  NAND2_X1 U717 ( .A1(n2005), .A2(n1361), .ZN(n1764) );
  NAND2_X1 U718 ( .A1(n2432), .A2(N458), .ZN(n1361) );
  NAND2_X1 U747 ( .A1(n2452), .A2(n1381), .ZN(n1774) );
  NAND2_X1 U748 ( .A1(n2429), .A2(N428), .ZN(n1381) );
  NAND2_X1 U750 ( .A1(n2452), .A2(n1383), .ZN(n1775) );
  NAND2_X1 U751 ( .A1(n2430), .A2(N425), .ZN(n1383) );
  NAND2_X1 U753 ( .A1(n2452), .A2(n1385), .ZN(n1776) );
  NAND2_X1 U754 ( .A1(n2430), .A2(N422), .ZN(n1385) );
  NAND2_X1 U756 ( .A1(n2452), .A2(n1387), .ZN(n1777) );
  NAND2_X1 U757 ( .A1(n2430), .A2(N419), .ZN(n1387) );
  NAND2_X1 U759 ( .A1(n2451), .A2(n1389), .ZN(n1778) );
  NAND2_X1 U760 ( .A1(n2429), .A2(N416), .ZN(n1389) );
  NAND2_X1 U762 ( .A1(n2451), .A2(n1391), .ZN(n1779) );
  NAND2_X1 U763 ( .A1(n2430), .A2(N413), .ZN(n1391) );
  NAND2_X1 U765 ( .A1(n2451), .A2(n1393), .ZN(n1780) );
  NAND2_X1 U766 ( .A1(n2429), .A2(N410), .ZN(n1393) );
  NAND2_X1 U768 ( .A1(n2451), .A2(n1395), .ZN(n1781) );
  NAND2_X1 U769 ( .A1(n2430), .A2(N407), .ZN(n1395) );
  NAND2_X1 U771 ( .A1(n2451), .A2(n1397), .ZN(n1782) );
  NAND2_X1 U772 ( .A1(n2429), .A2(N404), .ZN(n1397) );
  NAND2_X1 U774 ( .A1(n2451), .A2(n1399), .ZN(n1783) );
  NAND2_X1 U775 ( .A1(n2429), .A2(N401), .ZN(n1399) );
  NAND2_X1 U777 ( .A1(n2451), .A2(n1401), .ZN(n1784) );
  NAND2_X1 U778 ( .A1(n2430), .A2(N398), .ZN(n1401) );
  NAND2_X1 U780 ( .A1(n2451), .A2(n1403), .ZN(n1785) );
  NAND2_X1 U781 ( .A1(n2430), .A2(N395), .ZN(n1403) );
  NAND2_X1 U783 ( .A1(n2451), .A2(n1405), .ZN(n1786) );
  NAND2_X1 U784 ( .A1(n2430), .A2(N392), .ZN(n1405) );
  NAND2_X1 U786 ( .A1(n2451), .A2(n1407), .ZN(n1787) );
  NAND2_X1 U787 ( .A1(n2430), .A2(N389), .ZN(n1407) );
  NAND2_X1 U789 ( .A1(n2451), .A2(n1409), .ZN(n1788) );
  NAND2_X1 U790 ( .A1(n2430), .A2(N386), .ZN(n1409) );
  NAND2_X1 U792 ( .A1(n2451), .A2(n1411), .ZN(n1789) );
  NAND2_X1 U793 ( .A1(n2430), .A2(N383), .ZN(n1411) );
  NAND2_X1 U795 ( .A1(n2450), .A2(n1413), .ZN(n1790) );
  NAND2_X1 U796 ( .A1(n2429), .A2(N380), .ZN(n1413) );
  NAND2_X1 U798 ( .A1(n2450), .A2(n1415), .ZN(n1791) );
  NAND2_X1 U799 ( .A1(n2430), .A2(N377), .ZN(n1415) );
  NAND2_X1 U801 ( .A1(n2450), .A2(n1417), .ZN(n1792) );
  NAND2_X1 U802 ( .A1(n2430), .A2(N374), .ZN(n1417) );
  NAND2_X1 U804 ( .A1(n2450), .A2(n1419), .ZN(n1793) );
  NAND2_X1 U805 ( .A1(n2430), .A2(N371), .ZN(n1419) );
  NAND2_X1 U806 ( .A1(n2450), .A2(n1420), .ZN(n1794) );
  NAND2_X1 U807 ( .A1(n2430), .A2(N560), .ZN(n1420) );
  NAND2_X1 U809 ( .A1(n2450), .A2(n1424), .ZN(n1795) );
  NAND2_X1 U810 ( .A1(n2430), .A2(N557), .ZN(n1424) );
  NAND2_X1 U812 ( .A1(n2450), .A2(n1426), .ZN(n1796) );
  NAND2_X1 U813 ( .A1(n2430), .A2(N554), .ZN(n1426) );
  NAND2_X1 U815 ( .A1(n2450), .A2(n1428), .ZN(n1797) );
  NAND2_X1 U816 ( .A1(n2430), .A2(N551), .ZN(n1428) );
  NAND2_X1 U818 ( .A1(n2450), .A2(n1430), .ZN(n1798) );
  NAND2_X1 U819 ( .A1(n2431), .A2(N548), .ZN(n1430) );
  NAND2_X1 U821 ( .A1(n2450), .A2(n1432), .ZN(n1799) );
  NAND2_X1 U822 ( .A1(n2431), .A2(N545), .ZN(n1432) );
  NAND2_X1 U824 ( .A1(n2450), .A2(n1434), .ZN(n1800) );
  NAND2_X1 U825 ( .A1(n2431), .A2(N542), .ZN(n1434) );
  NAND2_X1 U827 ( .A1(n2450), .A2(n1436), .ZN(n1801) );
  NAND2_X1 U828 ( .A1(n2431), .A2(N539), .ZN(n1436) );
  NAND2_X1 U830 ( .A1(n2005), .A2(n1438), .ZN(n1802) );
  NAND2_X1 U831 ( .A1(n2431), .A2(N536), .ZN(n1438) );
  NAND2_X1 U833 ( .A1(n2005), .A2(n1440), .ZN(n1803) );
  NAND2_X1 U834 ( .A1(n2431), .A2(N533), .ZN(n1440) );
  NAND2_X1 U842 ( .A1(n2005), .A2(n1446), .ZN(n1806) );
  NAND2_X1 U843 ( .A1(n2431), .A2(N524), .ZN(n1446) );
  NAND2_X1 U845 ( .A1(n2005), .A2(n1448), .ZN(n1807) );
  NAND2_X1 U846 ( .A1(n2431), .A2(N521), .ZN(n1448) );
  NAND2_X1 U848 ( .A1(n2005), .A2(n1450), .ZN(n1808) );
  NAND2_X1 U849 ( .A1(n2431), .A2(N518), .ZN(n1450) );
  NAND2_X1 U851 ( .A1(n2005), .A2(n1452), .ZN(n1809) );
  NAND2_X1 U852 ( .A1(n2431), .A2(N515), .ZN(n1452) );
  NAND2_X1 U854 ( .A1(n2005), .A2(n1454), .ZN(n1810) );
  NAND2_X1 U855 ( .A1(n2431), .A2(N512), .ZN(n1454) );
  NAND2_X1 U857 ( .A1(n2005), .A2(n1456), .ZN(n1811) );
  NAND2_X1 U858 ( .A1(n2431), .A2(N509), .ZN(n1456) );
  NAND2_X1 U860 ( .A1(n2005), .A2(n1458), .ZN(n1812) );
  NAND2_X1 U861 ( .A1(n2431), .A2(N506), .ZN(n1458) );
  NAND2_X1 U863 ( .A1(n2005), .A2(n1460), .ZN(n1813) );
  NAND2_X1 U864 ( .A1(n2431), .A2(N503), .ZN(n1460) );
  NAND2_X1 U866 ( .A1(n2449), .A2(n1462), .ZN(n1814) );
  NAND2_X1 U867 ( .A1(n2431), .A2(N500), .ZN(n1462) );
  NAND2_X1 U869 ( .A1(n2449), .A2(n1464), .ZN(n1815) );
  NAND2_X1 U870 ( .A1(n2431), .A2(N497), .ZN(n1464) );
  NAND2_X1 U872 ( .A1(n2449), .A2(n1466), .ZN(n1816) );
  NAND2_X1 U873 ( .A1(n2431), .A2(N494), .ZN(n1466) );
  NAND2_X1 U875 ( .A1(n2449), .A2(n1468), .ZN(n1817) );
  NAND2_X1 U876 ( .A1(n2431), .A2(N491), .ZN(n1468) );
  NAND2_X1 U878 ( .A1(n2449), .A2(n1470), .ZN(n1818) );
  NAND2_X1 U879 ( .A1(n2432), .A2(N488), .ZN(n1470) );
  NAND2_X1 U881 ( .A1(n2449), .A2(n1472), .ZN(n1819) );
  NAND2_X1 U882 ( .A1(n2432), .A2(N485), .ZN(n1472) );
  NAND2_X1 U884 ( .A1(n2449), .A2(n1474), .ZN(n1820) );
  NAND2_X1 U885 ( .A1(n2432), .A2(N482), .ZN(n1474) );
  NAND2_X1 U887 ( .A1(n2449), .A2(n1476), .ZN(n1821) );
  NAND2_X1 U888 ( .A1(n2432), .A2(N479), .ZN(n1476) );
  NAND2_X1 U890 ( .A1(n2449), .A2(n1478), .ZN(n1822) );
  NAND2_X1 U891 ( .A1(n2432), .A2(N476), .ZN(n1478) );
  NAND2_X1 U893 ( .A1(n2449), .A2(n1480), .ZN(n1823) );
  NAND2_X1 U894 ( .A1(n2432), .A2(N473), .ZN(n1480) );
  NAND2_X1 U896 ( .A1(n2449), .A2(n1482), .ZN(n1824) );
  NAND2_X1 U897 ( .A1(n2429), .A2(N470), .ZN(n1482) );
  NAND2_X1 U899 ( .A1(n2449), .A2(n1484), .ZN(n1825) );
  NAND2_X1 U900 ( .A1(n2432), .A2(N467), .ZN(n1484) );
  AOI222_X1 U948 ( .A1(n2448), .A2(alu_output_EX_wire[2]), .B1(n2008), .B2(
        div_output_EX_wire[2]), .C1(mul_output_EX_wire[2]), .C2(n2011), .ZN(
        n1216) );
  AOI222_X1 U992 ( .A1(n2448), .A2(alu_output_EX_wire[1]), .B1(n2008), .B2(
        div_output_EX_wire[1]), .C1(mul_output_EX_wire[1]), .C2(n2011), .ZN(
        n1215) );
  AOI222_X1 U1041 ( .A1(n2448), .A2(alu_output_EX_wire[0]), .B1(n2011), .B2(
        mul_output_EX_wire[0]), .C1(n2008), .C2(div_output_EX_wire[0]), .ZN(
        n1214) );
  NOR3_X1 U1045 ( .A1(funct7_EX_reg[1]), .A2(funct7_EX_reg[2]), .A3(n1559), 
        .ZN(n1563) );
  NOR3_X1 U1047 ( .A1(funct7_EX_reg[4]), .A2(funct7_EX_reg[5]), .A3(n1166), 
        .ZN(n1562) );
  NOR4_X1 U1048 ( .A1(n2154), .A2(n2072), .A3(funct7_EX_reg[3]), .A4(
        funct7_EX_reg[6]), .ZN(n1561) );
  NOR2_X1 U1050 ( .A1(opcode_MW_reg[6]), .A2(opcode_MW_reg[3]), .ZN(n1565) );
  NOR2_X1 U1051 ( .A1(n2440), .A2(n1170), .ZN(N717) );
  NOR2_X1 U1052 ( .A1(n2438), .A2(n1171), .ZN(N716) );
  NOR2_X1 U1053 ( .A1(n2437), .A2(n1172), .ZN(N715) );
  AND2_X1 U1054 ( .A1(n2446), .A2(write_index_EX_reg[1]), .ZN(N714) );
  NOR2_X1 U1055 ( .A1(n2443), .A2(n1173), .ZN(N713) );
  AND2_X1 U1056 ( .A1(n2447), .A2(immediate_EX_reg[31]), .ZN(N712) );
  AND2_X1 U1057 ( .A1(n2447), .A2(immediate_EX_reg[30]), .ZN(N711) );
  AND2_X1 U1058 ( .A1(n2447), .A2(immediate_EX_reg[29]), .ZN(N710) );
  AND2_X1 U1059 ( .A1(n2447), .A2(immediate_EX_reg[28]), .ZN(N709) );
  AND2_X1 U1060 ( .A1(n2446), .A2(immediate_EX_reg[27]), .ZN(N708) );
  AND2_X1 U1061 ( .A1(n2446), .A2(immediate_EX_reg[26]), .ZN(N707) );
  AND2_X1 U1062 ( .A1(n2446), .A2(immediate_EX_reg[25]), .ZN(N706) );
  AND2_X1 U1063 ( .A1(n2446), .A2(immediate_EX_reg[24]), .ZN(N705) );
  AND2_X1 U1064 ( .A1(n2447), .A2(immediate_EX_reg[23]), .ZN(N704) );
  AND2_X1 U1065 ( .A1(n2446), .A2(immediate_EX_reg[22]), .ZN(N703) );
  AND2_X1 U1066 ( .A1(n2446), .A2(immediate_EX_reg[21]), .ZN(N702) );
  AND2_X1 U1067 ( .A1(n2446), .A2(immediate_EX_reg[20]), .ZN(N701) );
  AND2_X1 U1068 ( .A1(n2446), .A2(immediate_EX_reg[19]), .ZN(N700) );
  AND2_X1 U1069 ( .A1(n2445), .A2(immediate_EX_reg[18]), .ZN(N699) );
  AND2_X1 U1070 ( .A1(n2446), .A2(immediate_EX_reg[17]), .ZN(N698) );
  AND2_X1 U1071 ( .A1(n2446), .A2(immediate_EX_reg[16]), .ZN(N697) );
  AND2_X1 U1072 ( .A1(n2446), .A2(immediate_EX_reg[15]), .ZN(N696) );
  AND2_X1 U1073 ( .A1(n2445), .A2(immediate_EX_reg[14]), .ZN(N695) );
  AND2_X1 U1074 ( .A1(n2446), .A2(immediate_EX_reg[13]), .ZN(N694) );
  AND2_X1 U1075 ( .A1(n2446), .A2(immediate_EX_reg[12]), .ZN(N693) );
  AND2_X1 U1076 ( .A1(n2446), .A2(immediate_EX_reg[11]), .ZN(N692) );
  AND2_X1 U1077 ( .A1(n2446), .A2(immediate_EX_reg[10]), .ZN(N691) );
  AND2_X1 U1078 ( .A1(n2447), .A2(immediate_EX_reg[9]), .ZN(N690) );
  AND2_X1 U1079 ( .A1(n2446), .A2(immediate_EX_reg[8]), .ZN(N689) );
  AND2_X1 U1080 ( .A1(n2447), .A2(immediate_EX_reg[7]), .ZN(N688) );
  AND2_X1 U1081 ( .A1(n2446), .A2(immediate_EX_reg[6]), .ZN(N687) );
  AND2_X1 U1082 ( .A1(n2447), .A2(immediate_EX_reg[5]), .ZN(N686) );
  AND2_X1 U1083 ( .A1(n2447), .A2(immediate_EX_reg[4]), .ZN(N685) );
  AND2_X1 U1084 ( .A1(n2447), .A2(immediate_EX_reg[3]), .ZN(N684) );
  AND2_X1 U1085 ( .A1(n2447), .A2(immediate_EX_reg[2]), .ZN(N683) );
  AND2_X1 U1086 ( .A1(n2446), .A2(immediate_EX_reg[1]), .ZN(N682) );
  AND2_X1 U1087 ( .A1(n2446), .A2(immediate_EX_reg[0]), .ZN(N681) );
  AND2_X1 U1088 ( .A1(n2446), .A2(funct12_EX_reg[11]), .ZN(N680) );
  AND2_X1 U1089 ( .A1(n2447), .A2(funct12_EX_reg[10]), .ZN(N679) );
  AND2_X1 U1090 ( .A1(n2444), .A2(funct12_EX_reg[9]), .ZN(N678) );
  AND2_X1 U1091 ( .A1(n2444), .A2(funct12_EX_reg[8]), .ZN(N677) );
  AND2_X1 U1092 ( .A1(n2444), .A2(funct12_EX_reg[7]), .ZN(N676) );
  AND2_X1 U1093 ( .A1(n2444), .A2(funct12_EX_reg[6]), .ZN(N675) );
  AND2_X1 U1094 ( .A1(n2444), .A2(funct12_EX_reg[5]), .ZN(N674) );
  AND2_X1 U1095 ( .A1(n2444), .A2(funct12_EX_reg[4]), .ZN(N673) );
  AND2_X1 U1096 ( .A1(n2447), .A2(funct12_EX_reg[3]), .ZN(N672) );
  AND2_X1 U1097 ( .A1(n2446), .A2(funct12_EX_reg[2]), .ZN(N671) );
  AND2_X1 U1098 ( .A1(n2446), .A2(funct12_EX_reg[1]), .ZN(N670) );
  AND2_X1 U1099 ( .A1(n2445), .A2(funct12_EX_reg[0]), .ZN(N669) );
  AND2_X1 U1100 ( .A1(n2445), .A2(funct7_EX_reg[6]), .ZN(N668) );
  AND2_X1 U1101 ( .A1(n2446), .A2(funct7_EX_reg[5]), .ZN(N667) );
  AND2_X1 U1102 ( .A1(n2446), .A2(funct7_EX_reg[4]), .ZN(N666) );
  AND2_X1 U1103 ( .A1(n2446), .A2(funct7_EX_reg[3]), .ZN(N665) );
  AND2_X1 U1104 ( .A1(n2445), .A2(funct7_EX_reg[2]), .ZN(N664) );
  AND2_X1 U1105 ( .A1(n2445), .A2(funct7_EX_reg[1]), .ZN(N663) );
  AND2_X1 U1106 ( .A1(n2447), .A2(funct7_EX_reg[0]), .ZN(N662) );
  NOR2_X1 U1107 ( .A1(n2439), .A2(n1169), .ZN(N661) );
  AND2_X1 U1108 ( .A1(n2444), .A2(n2474), .ZN(N660) );
  AND2_X1 U1109 ( .A1(n2444), .A2(funct3_EX_reg[0]), .ZN(N659) );
  NOR2_X1 U1110 ( .A1(n2442), .A2(n1165), .ZN(N658) );
  NOR2_X1 U1111 ( .A1(n2441), .A2(n1166), .ZN(N657) );
  NAND2_X1 U1112 ( .A1(n2444), .A2(n1167), .ZN(N656) );
  NOR2_X1 U1114 ( .A1(n2443), .A2(n1168), .ZN(N654) );
  AND2_X1 U1115 ( .A1(n2446), .A2(write_enable_EX_reg), .ZN(N651) );
  NAND3_X1 U1119 ( .A1(write_enable_EX_reg), .A2(n1569), .A3(n1167), .ZN(n1568) );
  NAND4_X1 U1122 ( .A1(read_enable_1_FD_wire), .A2(n1570), .A3(n1571), .A4(
        n1572), .ZN(n1567) );
  XNOR2_X1 U1123 ( .A(write_index_EX_reg[1]), .B(read_index_1_FD_wire[1]), 
        .ZN(n1572) );
  AOI221_X1 U1124 ( .B1(n1170), .B2(read_index_1_FD_wire[4]), .C1(
        read_index_1_FD_wire[3]), .C2(n1171), .A(n1573), .ZN(n1571) );
  OAI22_X1 U1125 ( .A1(n1170), .A2(read_index_1_FD_wire[4]), .B1(n1171), .B2(
        read_index_1_FD_wire[3]), .ZN(n1573) );
  AOI221_X1 U1126 ( .B1(n1172), .B2(read_index_1_FD_wire[2]), .C1(
        read_index_1_FD_wire[0]), .C2(n1173), .A(n1574), .ZN(n1570) );
  OAI22_X1 U1127 ( .A1(n1172), .A2(read_index_1_FD_wire[2]), .B1(n1173), .B2(
        read_index_1_FD_wire[0]), .ZN(n1574) );
  NAND4_X1 U1128 ( .A1(read_enable_2_FD_wire), .A2(n1575), .A3(n1576), .A4(
        n1577), .ZN(n1566) );
  XNOR2_X1 U1129 ( .A(write_index_EX_reg[1]), .B(read_index_2_FD_wire[1]), 
        .ZN(n1577) );
  AOI221_X1 U1130 ( .B1(n1170), .B2(read_index_2_FD_wire[4]), .C1(
        read_index_2_FD_wire[3]), .C2(n1171), .A(n1578), .ZN(n1576) );
  OAI22_X1 U1131 ( .A1(n1170), .A2(read_index_2_FD_wire[4]), .B1(n1171), .B2(
        read_index_2_FD_wire[3]), .ZN(n1578) );
  AOI221_X1 U1132 ( .B1(n1172), .B2(read_index_2_FD_wire[2]), .C1(
        read_index_2_FD_wire[0]), .C2(n1173), .A(n1579), .ZN(n1575) );
  OAI22_X1 U1133 ( .A1(n1172), .A2(read_index_2_FD_wire[2]), .B1(n1173), .B2(
        read_index_2_FD_wire[0]), .ZN(n1579) );
  DFF_X2 \opcode_EX_reg_reg[0]  ( .D(n1743), .CK(clk), .Q(opcode_EX_reg[0]), 
        .QN(n1959) );
  DFF_X1 \opcode_EX_reg_reg[4]  ( .D(n1741), .CK(clk), .Q(opcode_EX_reg[4]), 
        .QN(n1167) );
  DFF_X1 \opcode_EX_reg_reg[2]  ( .D(n1161), .CK(clk), .Q(opcode_EX_reg[2]), 
        .QN(n1168) );
  DFF_X1 \opcode_EX_reg_reg[1]  ( .D(n1742), .CK(clk), .Q(opcode_EX_reg[1]), 
        .QN(n1960) );
  AOI22_X1 U447 ( .A1(n2444), .A2(n2091), .B1(n1183), .B2(n2443), .ZN(n1604)
         );
  AOI22_X1 U446 ( .A1(n2447), .A2(n2087), .B1(n1184), .B2(n2443), .ZN(n1603)
         );
  TBUF_X1 \instruction_FD_reg_tri[0]  ( .A(N290), .EN(N291), .Z(
        instruction_FD_reg[0]) );
  TBUF_X1 \instruction_FD_reg_tri[1]  ( .A(N287), .EN(N288), .Z(
        instruction_FD_reg[1]) );
  TBUF_X1 \instruction_FD_reg_tri[14]  ( .A(N248), .EN(N249), .Z(
        instruction_FD_reg[14]) );
  TBUF_X1 \instruction_FD_reg_tri[3]  ( .A(N281), .EN(N282), .Z(
        instruction_FD_reg[3]) );
  TBUF_X1 \instruction_FD_reg_tri[11]  ( .A(N257), .EN(N258), .Z(
        instruction_FD_reg[11]) );
  TBUF_X1 \instruction_FD_reg_tri[8]  ( .A(N266), .EN(N267), .Z(
        instruction_FD_reg[8]) );
  TBUF_X1 \instruction_FD_reg_tri[9]  ( .A(N263), .EN(N264), .Z(
        instruction_FD_reg[9]) );
  TBUF_X1 \instruction_FD_reg_tri[13]  ( .A(N251), .EN(N252), .Z(
        instruction_FD_reg[13]) );
  TBUF_X1 \instruction_FD_reg_tri[10]  ( .A(N260), .EN(N261), .Z(
        instruction_FD_reg[10]) );
  TBUF_X1 \instruction_FD_reg_tri[12]  ( .A(N254), .EN(N255), .Z(
        instruction_FD_reg[12]) );
  TBUF_X1 \instruction_FD_reg_tri[7]  ( .A(N269), .EN(N270), .Z(
        instruction_FD_reg[7]) );
  TBUF_X1 \instruction_FD_reg_tri[29]  ( .A(N203), .EN(N204), .Z(
        instruction_FD_reg[29]) );
  TBUF_X1 \instruction_FD_reg_tri[28]  ( .A(N206), .EN(N207), .Z(
        instruction_FD_reg[28]) );
  TBUF_X1 \instruction_FD_reg_tri[25]  ( .A(N215), .EN(N216), .Z(
        instruction_FD_reg[25]) );
  TBUF_X1 \instruction_FD_reg_tri[26]  ( .A(N212), .EN(N213), .Z(
        instruction_FD_reg[26]) );
  TBUF_X1 \instruction_FD_reg_tri[2]  ( .A(N284), .EN(N285), .Z(
        instruction_FD_reg[2]) );
  TBUF_X1 \instruction_FD_reg_tri[5]  ( .A(N275), .EN(N276), .Z(
        instruction_FD_reg[5]) );
  TBUF_X1 \instruction_FD_reg_tri[4]  ( .A(N278), .EN(N279), .Z(
        instruction_FD_reg[4]) );
  TBUF_X1 \instruction_FD_reg_tri[6]  ( .A(N272), .EN(N273), .Z(
        instruction_FD_reg[6]) );
  TBUF_X1 \instruction_FD_reg_tri[19]  ( .A(N233), .EN(N234), .Z(
        instruction_FD_reg[19]) );
  TBUF_X1 \instruction_FD_reg_tri[18]  ( .A(N236), .EN(N237), .Z(
        instruction_FD_reg[18]) );
  TBUF_X1 \instruction_FD_reg_tri[31]  ( .A(N197), .EN(N198), .Z(
        instruction_FD_reg[31]) );
  TBUF_X1 \instruction_FD_reg_tri[17]  ( .A(N239), .EN(N240), .Z(
        instruction_FD_reg[17]) );
  TBUF_X1 \instruction_FD_reg_tri[24]  ( .A(N218), .EN(N219), .Z(
        instruction_FD_reg[24]) );
  TBUF_X1 \instruction_FD_reg_tri[23]  ( .A(N221), .EN(N222), .Z(
        instruction_FD_reg[23]) );
  TBUF_X1 \instruction_FD_reg_tri[30]  ( .A(N200), .EN(N201), .Z(
        instruction_FD_reg[30]) );
  TBUF_X1 \instruction_FD_reg_tri[15]  ( .A(N245), .EN(N246), .Z(
        instruction_FD_reg[15]) );
  TBUF_X1 \instruction_FD_reg_tri[27]  ( .A(N209), .EN(N210), .Z(
        instruction_FD_reg[27]) );
  TBUF_X1 \instruction_FD_reg_tri[16]  ( .A(N242), .EN(N243), .Z(
        instruction_FD_reg[16]) );
  TBUF_X1 \instruction_FD_reg_tri[22]  ( .A(N224), .EN(N225), .Z(
        instruction_FD_reg[22]) );
  TBUF_X1 \instruction_FD_reg_tri[20]  ( .A(N230), .EN(N231), .Z(
        instruction_FD_reg[20]) );
  TBUF_X1 \instruction_FD_reg_tri[21]  ( .A(N227), .EN(N228), .Z(
        instruction_FD_reg[21]) );
  INV_X1 U414 ( .A(n1323), .ZN(n1161) );
  INV_X1 U411 ( .A(n1349), .ZN(n1158) );
  INV_X1 U412 ( .A(n1348), .ZN(n1159) );
  INV_X1 U409 ( .A(n1352), .ZN(n1156) );
  INV_X1 U410 ( .A(n1350), .ZN(n1157) );
  INV_X1 U413 ( .A(n1326), .ZN(n1160) );
  INV_X1 U383 ( .A(next_pc_FD_wire[6]), .ZN(n1130) );
  INV_X1 U384 ( .A(next_pc_FD_wire[7]), .ZN(n1131) );
  INV_X1 U382 ( .A(next_pc_FD_wire[5]), .ZN(n1129) );
  INV_X1 U377 ( .A(next_pc_FD_wire[0]), .ZN(n1124) );
  INV_X1 U379 ( .A(next_pc_FD_wire[2]), .ZN(n1126) );
  INV_X1 U380 ( .A(next_pc_FD_wire[3]), .ZN(n1127) );
  INV_X1 U378 ( .A(next_pc_FD_wire[1]), .ZN(n1125) );
  INV_X1 U381 ( .A(next_pc_FD_wire[4]), .ZN(n1128) );
  INV_X1 U49 ( .A(rs2_EX_reg[21]), .ZN(n23) );
  INV_X1 U15 ( .A(rs2_EX_reg[4]), .ZN(n6) );
  INV_X1 U53 ( .A(rs2_EX_reg[23]), .ZN(n25) );
  INV_X1 U41 ( .A(rs2_EX_reg[17]), .ZN(n19) );
  INV_X1 U55 ( .A(rs2_EX_reg[24]), .ZN(n26) );
  INV_X1 U61 ( .A(rs2_EX_reg[27]), .ZN(n29) );
  INV_X1 U63 ( .A(rs2_EX_reg[28]), .ZN(n30) );
  INV_X1 U67 ( .A(rs2_EX_reg[30]), .ZN(n32) );
  INV_X1 U57 ( .A(rs2_EX_reg[25]), .ZN(n27) );
  INV_X1 U65 ( .A(rs2_EX_reg[29]), .ZN(n31) );
  INV_X1 U59 ( .A(rs2_EX_reg[26]), .ZN(n28) );
  INV_X1 U47 ( .A(rs2_EX_reg[20]), .ZN(n22) );
  INV_X1 U37 ( .A(rs2_EX_reg[15]), .ZN(n17) );
  INV_X1 U17 ( .A(rs2_EX_reg[5]), .ZN(n7) );
  INV_X1 U45 ( .A(rs2_EX_reg[19]), .ZN(n21) );
  INV_X1 U23 ( .A(rs2_EX_reg[8]), .ZN(n10) );
  INV_X1 U25 ( .A(rs2_EX_reg[9]), .ZN(n11) );
  INV_X1 U31 ( .A(rs2_EX_reg[12]), .ZN(n14) );
  INV_X1 U19 ( .A(rs2_EX_reg[6]), .ZN(n8) );
  INV_X1 U27 ( .A(rs2_EX_reg[10]), .ZN(n12) );
  INV_X1 U11 ( .A(rs2_EX_reg[2]), .ZN(n4) );
  INV_X1 U9 ( .A(rs2_EX_reg[1]), .ZN(n3) );
  INV_X1 U4 ( .A(rs2_EX_reg[0]), .ZN(n1) );
  INV_X1 U29 ( .A(rs2_EX_reg[11]), .ZN(n13) );
  INV_X1 U13 ( .A(rs2_EX_reg[3]), .ZN(n5) );
  INV_X1 U39 ( .A(rs2_EX_reg[16]), .ZN(n18) );
  INV_X1 U33 ( .A(rs2_EX_reg[13]), .ZN(n15) );
  INV_X1 U43 ( .A(rs2_EX_reg[18]), .ZN(n20) );
  NAND2_X1 U1121 ( .A1(opcode_EX_reg[0]), .A2(opcode_EX_reg[1]), .ZN(n1564) );
  DFF_X2 \rs2_EX_reg_reg[28]  ( .D(n2505), .CK(clk), .Q(), .QN(N475) );
  MUX2_X1 U707 ( .A(csr_index_EX_reg[0]), .B(csr_index_FD_wire[0]), .S(n2466), 
        .Z(n1760) );
  DFF_X1 \opcode_EX_reg_reg[6]  ( .D(n1163), .CK(clk), .Q(opcode_EX_reg[6]), 
        .QN(n1165) );
  DFF_X2 \rs2_EX_reg_reg[19]  ( .D(n1461), .CK(clk), .Q(), .QN(N502) );
  DFF_X2 \rs2_EX_reg_reg[16]  ( .D(n1455), .CK(clk), .Q(), .QN(N511) );
  DFF_X2 \rs1_EX_reg_reg[19]  ( .D(n1396), .CK(clk), .Q(), .QN(N406) );
  DFF_X2 \rs1_EX_reg_reg[16]  ( .D(n1390), .CK(clk), .Q(), .QN(N415) );
  DFF_X2 \rs1_EX_reg_reg[28]  ( .D(n2506), .CK(clk), .Q(), .QN(N379) );
  DFF_X2 \rs2_EX_reg_reg[23]  ( .D(n1469), .CK(clk), .Q(), .QN(N490) );
  DFF_X2 \rs1_EX_reg_reg[23]  ( .D(n1404), .CK(clk), .Q(), .QN(N394) );
  DFF_X1 \opcode_EX_reg_reg[3]  ( .D(n1322), .CK(clk), .Q(), .QN(
        opcode_EX_reg[3]) );
  DFF_X2 \rs2_EX_reg_reg[10]  ( .D(n1443), .CK(clk), .Q(), .QN(N529) );
  DFF_X1 \rs2_EX_reg_reg[31]  ( .D(n2508), .CK(clk), .Q(), .QN(N466) );
  DFF_X1 \rs1_EX_reg_reg[31]  ( .D(n2507), .CK(clk), .Q(), .QN(N370) );
  DFF_X2 \rs1_EX_reg_reg[5]  ( .D(n1368), .CK(clk), .Q(), .QN(N448) );
  DFF_X2 \rs2_EX_reg_reg[5]  ( .D(n1433), .CK(clk), .Q(), .QN(N544) );
  AOI211_X1 U1118 ( .C1(n1566), .C2(n1567), .A(n1564), .B(n1568), .ZN(n1485)
         );
  NAND2_X2 U1116 ( .A1(n1354), .A2(n2475), .ZN(N193) );
  DFF_X2 \rs1_EX_reg_reg[3]  ( .D(n1364), .CK(clk), .Q(), .QN(N454) );
  DFF_X1 \opcode_MW_reg_reg[1]  ( .D(n1962), .CK(clk), .Q(opcode_MW_reg[1]), 
        .QN(n788) );
  DFF_X1 \opcode_MW_reg_reg[0]  ( .D(n1961), .CK(clk), .Q(opcode_MW_reg[0]), 
        .QN(n787) );
  DFF_X1 \opcode_EX_reg_reg[5]  ( .D(n1320), .CK(clk), .Q(n1166), .QN(
        opcode_EX_reg[5]) );
  TBUF_X2 \rs1_EX_reg_tri[10]  ( .A(N433), .EN(N434), .Z(rs1_EX_reg[10]) );
  TBUF_X2 \rs1_EX_reg_tri[0]  ( .A(N463), .EN(N464), .Z(rs1_EX_reg[0]) );
  TBUF_X2 \rs1_EX_reg_tri[1]  ( .A(N460), .EN(N461), .Z(rs1_EX_reg[1]) );
  DFF_X2 \rs2_EX_reg_reg[24]  ( .D(n1471), .CK(clk), .Q(), .QN(N487) );
  DFF_X2 \rs1_EX_reg_reg[24]  ( .D(n1406), .CK(clk), .Q(), .QN(N391) );
  AOI21_X1 U1134 ( .B1(mul_output_EX_wire[12]), .B2(n2011), .A(n2241), .ZN(
        n1827) );
  CLKBUF_X1 U1135 ( .A(address_EX_wire[28]), .Z(n2093) );
  AOI222_X2 U1136 ( .A1(n2448), .A2(alu_output_EX_wire[30]), .B1(n2008), .B2(
        div_output_EX_wire[30]), .C1(mul_output_EX_wire[30]), .C2(n2011), .ZN(
        n1244) );
  AND2_X2 U1137 ( .A1(n2136), .A2(n2137), .ZN(n1830) );
  INV_X4 U1138 ( .A(n1830), .ZN(n2135) );
  CLKBUF_X1 U1139 ( .A(address_EX_wire[23]), .Z(n2098) );
  CLKBUF_X2 U1140 ( .A(n1235), .Z(n1831) );
  CLKBUF_X1 U1141 ( .A(n2103), .Z(n1909) );
  CLKBUF_X1 U1142 ( .A(address_EX_wire[24]), .Z(n2097) );
  OAI21_X1 U1143 ( .B1(n1235), .B2(n1488), .A(n2308), .ZN(n1832) );
  AOI21_X2 U1144 ( .B1(mul_output_EX_wire[21]), .B2(n2011), .A(n2232), .ZN(
        n1235) );
  AOI222_X1 U1145 ( .A1(n2448), .A2(alu_output_EX_wire[1]), .B1(n2008), .B2(
        div_output_EX_wire[1]), .C1(mul_output_EX_wire[1]), .C2(n2011), .ZN(
        n1833) );
  AND2_X2 U1146 ( .A1(n2477), .A2(n1166), .ZN(n2504) );
  NAND2_X1 U1147 ( .A1(address_EX_wire[31]), .A2(n2504), .ZN(n1834) );
  NAND2_X1 U1148 ( .A1(n1834), .A2(n1969), .ZN(n1910) );
  NAND2_X1 U1149 ( .A1(n1898), .A2(n1897), .ZN(\_2_net_[23] ) );
  AOI21_X1 U1150 ( .B1(FW_source_1[23]), .B2(n2422), .A(n1903), .ZN(n1404) );
  AOI21_X1 U1151 ( .B1(FW_source_2[31]), .B2(n2501), .A(n1838), .ZN(n2508) );
  NAND2_X1 U1152 ( .A1(n2429), .A2(N370), .ZN(n1837) );
  NAND2_X1 U1153 ( .A1(n2268), .A2(RF_source_1[31]), .ZN(n1836) );
  NAND2_X1 U1154 ( .A1(n1836), .A2(n1837), .ZN(n1835) );
  AOI21_X1 U1155 ( .B1(FW_source_1[31]), .B2(n2500), .A(n1835), .ZN(n2507) );
  NAND2_X1 U1156 ( .A1(n2007), .A2(N466), .ZN(n1840) );
  NAND2_X1 U1157 ( .A1(n2004), .A2(RF_source_2[31]), .ZN(n1839) );
  NAND2_X1 U1158 ( .A1(n1839), .A2(n1840), .ZN(n1838) );
  INV_X2 U1159 ( .A(n1844), .ZN(n1843) );
  NAND2_X2 U1160 ( .A1(n2448), .A2(alu_output_EX_wire[4]), .ZN(n1844) );
  AOI21_X1 U1161 ( .B1(mul_output_EX_wire[4]), .B2(n2011), .A(n1843), .ZN(
        n1841) );
  AND2_X1 U1162 ( .A1(n1841), .A2(n1842), .ZN(n1218) );
  NAND2_X1 U1163 ( .A1(div_output_EX_wire[4]), .A2(n2008), .ZN(n1842) );
  NAND2_X1 U1164 ( .A1(n2293), .A2(immediate_EX_reg[4]), .ZN(n1848) );
  NAND2_X1 U1165 ( .A1(csr_rd_EX_wire[4]), .A2(n2436), .ZN(n1847) );
  NAND2_X1 U1166 ( .A1(n1847), .A2(n1848), .ZN(n1846) );
  AOI21_X1 U1167 ( .B1(address_EX_wire[4]), .B2(n2504), .A(n1846), .ZN(n1845)
         );
  OAI21_X1 U1168 ( .B1(n1218), .B2(n1488), .A(n1845), .ZN(\_2_net_[4] ) );
  NAND2_X1 U1169 ( .A1(n2429), .A2(N451), .ZN(n1851) );
  NAND2_X1 U1170 ( .A1(n2268), .A2(RF_source_1[4]), .ZN(n1850) );
  NAND2_X1 U1171 ( .A1(n1850), .A2(n1851), .ZN(n1849) );
  AOI21_X1 U1172 ( .B1(FW_source_1[4]), .B2(n2500), .A(n1849), .ZN(n1366) );
  NAND2_X1 U1173 ( .A1(n2429), .A2(N547), .ZN(n1854) );
  NAND2_X1 U1174 ( .A1(n2004), .A2(RF_source_2[4]), .ZN(n1853) );
  NAND2_X1 U1175 ( .A1(n1853), .A2(n1854), .ZN(n1852) );
  AOI21_X1 U1176 ( .B1(FW_source_2[4]), .B2(n2501), .A(n1852), .ZN(n1431) );
  AND2_X2 U1177 ( .A1(n2443), .A2(n1185), .ZN(n1856) );
  AOI21_X1 U1178 ( .B1(n2011), .B2(mul_output_EX_wire[22]), .A(n1859), .ZN(
        n1855) );
  AOI21_X1 U1179 ( .B1(n1857), .B2(n2445), .A(n1856), .ZN(n1602) );
  OR2_X1 U1180 ( .A1(n1855), .A2(n1488), .ZN(n1858) );
  BUF_X1 U1181 ( .A(n1855), .Z(n1857) );
  OAI211_X1 U1182 ( .C1(n2080), .C2(n2081), .A(n1858), .B(n2104), .ZN(n2055)
         );
  OAI211_X1 U1183 ( .C1(n2080), .C2(n2081), .A(n1858), .B(n2104), .ZN(
        \_2_net_[22] ) );
  NAND2_X1 U1184 ( .A1(n2448), .A2(alu_output_EX_wire[22]), .ZN(n1861) );
  NAND2_X1 U1185 ( .A1(div_output_EX_wire[22]), .A2(n2502), .ZN(n1860) );
  NAND2_X1 U1186 ( .A1(n1860), .A2(n1861), .ZN(n1859) );
  INV_X2 U1187 ( .A(n1488), .ZN(n1862) );
  AND2_X2 U1188 ( .A1(n2437), .A2(n1197), .ZN(n1864) );
  OR2_X1 U1189 ( .A1(n1865), .A2(n1894), .ZN(n1866) );
  NAND2_X1 U1190 ( .A1(n1866), .A2(n1862), .ZN(n2027) );
  AND2_X1 U1191 ( .A1(mul_output_EX_wire[10]), .A2(n2011), .ZN(n1865) );
  BUF_X1 U1192 ( .A(n1865), .Z(n1867) );
  NOR2_X1 U1193 ( .A1(n1867), .A2(n1894), .ZN(n1863) );
  AOI21_X1 U1194 ( .B1(n1863), .B2(n2446), .A(n1864), .ZN(n1590) );
  NAND2_X1 U1195 ( .A1(n2027), .A2(n2023), .ZN(\_2_net_[10] ) );
  AOI21_X1 U1196 ( .B1(FW_source_2[10]), .B2(n2501), .A(n2028), .ZN(n1443) );
  NAND2_X1 U1197 ( .A1(n1494), .A2(alu_output_EX_wire[9]), .ZN(n1870) );
  NAND2_X1 U1198 ( .A1(div_output_EX_wire[9]), .A2(n2435), .ZN(n1869) );
  NAND2_X1 U1199 ( .A1(n1869), .A2(n1870), .ZN(n1868) );
  AOI21_X1 U1200 ( .B1(mul_output_EX_wire[9]), .B2(n2011), .A(n1868), .ZN(
        n1223) );
  OR2_X1 U1201 ( .A1(n2418), .A2(n2175), .ZN(n1874) );
  NAND2_X1 U1202 ( .A1(csr_rd_EX_wire[9]), .A2(n2436), .ZN(n1873) );
  NAND2_X1 U1203 ( .A1(n1873), .A2(n1874), .ZN(n1872) );
  AOI21_X1 U1204 ( .B1(address_EX_wire[9]), .B2(n2479), .A(n1872), .ZN(n1871)
         );
  OAI21_X1 U1205 ( .B1(n1223), .B2(n1488), .A(n1871), .ZN(\_2_net_[9] ) );
  NAND2_X1 U1206 ( .A1(n2428), .A2(N436), .ZN(n1877) );
  NAND2_X1 U1207 ( .A1(n2424), .A2(RF_source_1[9]), .ZN(n1876) );
  NAND2_X1 U1208 ( .A1(n1876), .A2(n1877), .ZN(n1875) );
  AOI21_X1 U1209 ( .B1(FW_source_1[9]), .B2(n2422), .A(n1875), .ZN(n1376) );
  NAND2_X1 U1210 ( .A1(n2427), .A2(N532), .ZN(n1880) );
  NAND2_X1 U1211 ( .A1(n2004), .A2(RF_source_2[9]), .ZN(n1879) );
  NAND2_X1 U1212 ( .A1(n1879), .A2(n1880), .ZN(n1878) );
  AOI21_X1 U1213 ( .B1(FW_source_2[9]), .B2(n2425), .A(n1878), .ZN(n1441) );
  AOI21_X2 U1214 ( .B1(n1883), .B2(n1884), .A(n1885), .ZN(n1882) );
  NAND2_X2 U1215 ( .A1(n1886), .A2(n1887), .ZN(n1885) );
  INV_X2 U1216 ( .A(n1888), .ZN(n1887) );
  NOR2_X2 U1217 ( .A1(n2418), .A2(n2158), .ZN(n1888) );
  NAND2_X2 U1218 ( .A1(csr_rd_EX_wire[24]), .A2(n2436), .ZN(n1886) );
  INV_X2 U1219 ( .A(n1488), .ZN(n1884) );
  NAND2_X1 U1220 ( .A1(address_EX_wire[24]), .A2(n2479), .ZN(n1881) );
  NAND2_X1 U1221 ( .A1(n1881), .A2(n1882), .ZN(\_2_net_[24] ) );
  INV_X1 U1222 ( .A(n2100), .ZN(n1889) );
  NAND2_X1 U1223 ( .A1(n1889), .A2(n1890), .ZN(n1883) );
  NAND2_X1 U1224 ( .A1(mul_output_EX_wire[24]), .A2(n2011), .ZN(n1890) );
  NAND2_X1 U1225 ( .A1(n2426), .A2(N391), .ZN(n1893) );
  NAND2_X1 U1226 ( .A1(n2268), .A2(RF_source_1[24]), .ZN(n1892) );
  NAND2_X1 U1227 ( .A1(n1892), .A2(n1893), .ZN(n1891) );
  AOI21_X1 U1228 ( .B1(FW_source_1[24]), .B2(n2422), .A(n1891), .ZN(n1406) );
  NAND2_X2 U1229 ( .A1(n1494), .A2(alu_output_EX_wire[10]), .ZN(n1896) );
  NAND2_X1 U1230 ( .A1(div_output_EX_wire[10]), .A2(n2435), .ZN(n1895) );
  NAND2_X1 U1231 ( .A1(n1895), .A2(n1896), .ZN(n1894) );
  AOI22_X1 U1232 ( .A1(csr_rd_EX_wire[23]), .A2(n2436), .B1(
        immediate_EX_reg[23]), .B2(n2293), .ZN(n1902) );
  NAND2_X1 U1233 ( .A1(mul_output_EX_wire[23]), .A2(n2011), .ZN(n1899) );
  INV_X1 U1234 ( .A(n1902), .ZN(n1901) );
  NAND2_X1 U1235 ( .A1(n1899), .A2(n1830), .ZN(n1900) );
  AOI21_X1 U1236 ( .B1(n1900), .B2(n2144), .A(n1901), .ZN(n1897) );
  NAND2_X1 U1237 ( .A1(address_EX_wire[23]), .A2(n2479), .ZN(n1898) );
  NAND2_X1 U1238 ( .A1(n2426), .A2(N394), .ZN(n1905) );
  NAND2_X1 U1239 ( .A1(n2424), .A2(RF_source_1[23]), .ZN(n1904) );
  NAND2_X1 U1240 ( .A1(n1904), .A2(n1905), .ZN(n1903) );
  NAND2_X1 U1241 ( .A1(n2007), .A2(N490), .ZN(n1908) );
  NAND2_X1 U1242 ( .A1(n2269), .A2(RF_source_2[23]), .ZN(n1907) );
  NAND2_X1 U1243 ( .A1(n1907), .A2(n1908), .ZN(n1906) );
  AOI21_X1 U1244 ( .B1(FW_source_2[23]), .B2(n2425), .A(n1906), .ZN(n1469) );
  BUF_X1 U1245 ( .A(n1827), .Z(n1911) );
  AOI21_X1 U1246 ( .B1(mul_output_EX_wire[11]), .B2(n2011), .A(n2238), .ZN(
        n1912) );
  AOI21_X1 U1247 ( .B1(mul_output_EX_wire[14]), .B2(n2011), .A(n2244), .ZN(
        n1913) );
  NAND2_X1 U1248 ( .A1(n2448), .A2(alu_output_EX_wire[19]), .ZN(n1990) );
  NAND2_X1 U1249 ( .A1(n2448), .A2(alu_output_EX_wire[29]), .ZN(n2002) );
  NAND2_X1 U1250 ( .A1(csr_rd_EX_wire[29]), .A2(n2436), .ZN(n1999) );
  NAND2_X1 U1251 ( .A1(csr_rd_EX_wire[3]), .A2(n2436), .ZN(n1979) );
  NAND2_X1 U1252 ( .A1(n2293), .A2(immediate_EX_reg[3]), .ZN(n1980) );
  NAND2_X1 U1253 ( .A1(n1986), .A2(n1990), .ZN(n1989) );
  NAND2_X1 U1254 ( .A1(n1999), .A2(n1957), .ZN(n1998) );
  NAND2_X1 U1255 ( .A1(n1979), .A2(n1980), .ZN(n1978) );
  NAND2_X1 U1256 ( .A1(n2448), .A2(alu_output_EX_wire[28]), .ZN(n2124) );
  NAND2_X1 U1257 ( .A1(n2448), .A2(alu_output_EX_wire[24]), .ZN(n2102) );
  NAND2_X1 U1258 ( .A1(n2448), .A2(alu_output_EX_wire[23]), .ZN(n2137) );
  NAND2_X1 U1259 ( .A1(n2448), .A2(alu_output_EX_wire[31]), .ZN(n2064) );
  NAND2_X1 U1260 ( .A1(csr_rd_EX_wire[6]), .A2(n2436), .ZN(n1914) );
  OAI21_X1 U1261 ( .B1(n2168), .B2(n2418), .A(n1914), .ZN(n1915) );
  AOI21_X1 U1262 ( .B1(address_EX_wire[6]), .B2(n2479), .A(n1915), .ZN(n1916)
         );
  OAI21_X1 U1263 ( .B1(n1220), .B2(n1488), .A(n1916), .ZN(\_2_net_[6] ) );
  AOI222_X1 U1264 ( .A1(address_EX_wire[17]), .A2(n2421), .B1(
        next_pc_FD_wire[17]), .B2(n2496), .C1(pc_FD_reg[17]), .C2(n2420), .ZN(
        n1917) );
  INV_X1 U1265 ( .A(n1917), .ZN(n1641) );
  NAND2_X1 U1266 ( .A1(N431), .A2(n2430), .ZN(n1918) );
  NAND2_X1 U1267 ( .A1(n2452), .A2(n1918), .ZN(n1773) );
  AOI222_X1 U1268 ( .A1(n2010), .A2(n2421), .B1(next_pc_FD_wire[16]), .B2(
        n2496), .C1(pc_FD_reg[16]), .C2(n2420), .ZN(n1919) );
  INV_X1 U1269 ( .A(n1919), .ZN(n1643) );
  NAND2_X1 U1270 ( .A1(N527), .A2(n2431), .ZN(n1920) );
  NAND2_X1 U1271 ( .A1(n2005), .A2(n1920), .ZN(n1805) );
  INV_X1 U1272 ( .A(n2430), .ZN(n1921) );
  OAI21_X1 U1273 ( .B1(n2085), .B2(n1921), .A(n2452), .ZN(n1772) );
  AOI222_X1 U1274 ( .A1(address_EX_wire[15]), .A2(n2421), .B1(
        next_pc_FD_wire[15]), .B2(n2496), .C1(pc_FD_reg[15]), .C2(n2420), .ZN(
        n1922) );
  INV_X1 U1275 ( .A(n1922), .ZN(n1645) );
  NAND2_X1 U1276 ( .A1(N530), .A2(n2431), .ZN(n1923) );
  NAND2_X1 U1277 ( .A1(n2005), .A2(n1923), .ZN(n1804) );
  NAND2_X1 U1278 ( .A1(N437), .A2(n2429), .ZN(n1924) );
  NAND2_X1 U1279 ( .A1(n2452), .A2(n1924), .ZN(n1771) );
  NOR2_X1 U1280 ( .A1(n2418), .A2(n2157), .ZN(n1925) );
  AOI21_X1 U1281 ( .B1(csr_rd_EX_wire[19]), .B2(n2436), .A(n1925), .ZN(n1986)
         );
  AOI22_X1 U1282 ( .A1(opcode_FD_wire[1]), .A2(n2470), .B1(n2428), .B2(
        opcode_EX_reg[1]), .ZN(n1926) );
  NAND2_X1 U1283 ( .A1(n2005), .A2(n1926), .ZN(n1742) );
  AOI222_X1 U1284 ( .A1(address_EX_wire[14]), .A2(n2421), .B1(
        next_pc_FD_wire[14]), .B2(n2496), .C1(pc_FD_reg[14]), .C2(n2420), .ZN(
        n1927) );
  INV_X1 U1285 ( .A(n1927), .ZN(n1647) );
  NAND2_X1 U1286 ( .A1(N449), .A2(n2432), .ZN(n1928) );
  NAND2_X1 U1287 ( .A1(n2452), .A2(n1928), .ZN(n1767) );
  AOI22_X1 U1288 ( .A1(csr_rd_EX_wire[28]), .A2(n2436), .B1(n2293), .B2(
        immediate_EX_reg[28]), .ZN(n1929) );
  INV_X1 U1289 ( .A(n1929), .ZN(n1966) );
  AOI222_X1 U1290 ( .A1(address_EX_wire[11]), .A2(n2421), .B1(
        next_pc_FD_wire[11]), .B2(n2496), .C1(pc_FD_reg[11]), .C2(n2420), .ZN(
        n1930) );
  INV_X1 U1291 ( .A(n1930), .ZN(n1653) );
  AOI22_X1 U1292 ( .A1(instruction_type_EX_reg[0]), .A2(n2007), .B1(
        instruction_type_FD_wire[0]), .B2(n2465), .ZN(n1931) );
  NAND2_X1 U1293 ( .A1(n2005), .A2(n1931), .ZN(n1708) );
  NAND2_X1 U1294 ( .A1(N452), .A2(n2432), .ZN(n1932) );
  NAND2_X1 U1295 ( .A1(n2452), .A2(n1932), .ZN(n1766) );
  AOI222_X1 U1296 ( .A1(address_EX_wire[10]), .A2(n2421), .B1(
        next_pc_FD_wire[10]), .B2(n2496), .C1(pc_FD_reg[10]), .C2(n2420), .ZN(
        n1933) );
  INV_X1 U1297 ( .A(n1933), .ZN(n1655) );
  NAND2_X1 U1298 ( .A1(N440), .A2(n2429), .ZN(n1934) );
  NAND2_X1 U1299 ( .A1(n2452), .A2(n1934), .ZN(n1770) );
  NAND2_X1 U1300 ( .A1(N455), .A2(n2432), .ZN(n1935) );
  NAND2_X1 U1301 ( .A1(n2005), .A2(n1935), .ZN(n1765) );
  AOI222_X1 U1302 ( .A1(n2006), .A2(n2090), .B1(next_pc_FD_wire[19]), .B2(
        n2496), .C1(pc_FD_reg[19]), .C2(n2419), .ZN(n1936) );
  INV_X1 U1303 ( .A(n1936), .ZN(n1637) );
  OAI22_X1 U1304 ( .A1(address_MW_reg[2]), .A2(n2444), .B1(n2438), .B2(
        address_EX_wire[2]), .ZN(n1937) );
  INV_X1 U1305 ( .A(n1937), .ZN(n916) );
  OAI22_X1 U1306 ( .A1(address_MW_reg[0]), .A2(n2444), .B1(n2440), .B2(
        address_EX_wire[0]), .ZN(n1938) );
  INV_X1 U1307 ( .A(n1938), .ZN(n918) );
  NAND2_X1 U1308 ( .A1(N443), .A2(n2429), .ZN(n1939) );
  NAND2_X1 U1309 ( .A1(n2452), .A2(n1939), .ZN(n1769) );
  NAND2_X1 U1310 ( .A1(N461), .A2(n2432), .ZN(n1940) );
  NAND2_X1 U1311 ( .A1(n2005), .A2(n1940), .ZN(n1763) );
  NAND2_X1 U1312 ( .A1(n2436), .A2(csr_rd_EX_wire[20]), .ZN(n1941) );
  OAI21_X1 U1313 ( .B1(n2167), .B2(n2418), .A(n1941), .ZN(n2307) );
  NAND2_X1 U1314 ( .A1(n2436), .A2(csr_rd_EX_wire[13]), .ZN(n1942) );
  OAI21_X1 U1315 ( .B1(n2176), .B2(n2418), .A(n1942), .ZN(n2325) );
  NAND2_X1 U1316 ( .A1(n2436), .A2(csr_rd_EX_wire[16]), .ZN(n1943) );
  OAI21_X1 U1317 ( .B1(n2174), .B2(n2418), .A(n1943), .ZN(n2126) );
  AND2_X1 U1318 ( .A1(alu_output_EX_wire[18]), .A2(n2448), .ZN(n1944) );
  AOI211_X1 U1319 ( .C1(mul_output_EX_wire[18]), .C2(n2011), .A(n1944), .B(
        n2323), .ZN(n1232) );
  AOI22_X1 U1320 ( .A1(n2470), .A2(opcode_FD_wire[3]), .B1(n2428), .B2(n2077), 
        .ZN(n1322) );
  AOI222_X1 U1321 ( .A1(alu_output_EX_wire[29]), .A2(n2448), .B1(n2011), .B2(
        mul_output_EX_wire[29]), .C1(div_output_EX_wire[29]), .C2(n2008), .ZN(
        n1945) );
  AOI22_X1 U1322 ( .A1(n2442), .A2(n1178), .B1(n1945), .B2(n2444), .ZN(n1609)
         );
  AOI211_X1 U1323 ( .C1(mul_output_EX_wire[25]), .C2(n2011), .A(n2291), .B(
        n2292), .ZN(n1946) );
  AOI22_X1 U1324 ( .A1(n2443), .A2(n1182), .B1(n1946), .B2(n2446), .ZN(n1605)
         );
  AOI222_X1 U1325 ( .A1(alu_output_EX_wire[3]), .A2(n2448), .B1(n2011), .B2(
        mul_output_EX_wire[3]), .C1(div_output_EX_wire[3]), .C2(n2008), .ZN(
        n1947) );
  AOI22_X1 U1326 ( .A1(n2439), .A2(n1204), .B1(n1947), .B2(n2444), .ZN(n1583)
         );
  AOI222_X1 U1327 ( .A1(address_EX_wire[13]), .A2(n2421), .B1(
        next_pc_FD_wire[13]), .B2(n2496), .C1(pc_FD_reg[13]), .C2(n2420), .ZN(
        n1948) );
  INV_X1 U1328 ( .A(n1948), .ZN(n1649) );
  OAI22_X1 U1329 ( .A1(address_MW_reg[1]), .A2(n2444), .B1(n2437), .B2(
        address_EX_wire[1]), .ZN(n1949) );
  INV_X1 U1330 ( .A(n1949), .ZN(n917) );
  INV_X1 U1331 ( .A(rs2_EX_reg[22]), .ZN(n1950) );
  AOI22_X1 U1332 ( .A1(n2439), .A2(n234), .B1(n2444), .B2(n1950), .ZN(n1100)
         );
  INV_X1 U1333 ( .A(rs2_EX_reg[14]), .ZN(n1951) );
  AOI22_X1 U1334 ( .A1(n2439), .A2(n226), .B1(n2444), .B2(n1951), .ZN(n1108)
         );
  INV_X1 U1335 ( .A(rs2_EX_reg[7]), .ZN(n1952) );
  AOI22_X1 U1336 ( .A1(n2443), .A2(n219), .B1(n2444), .B2(n1952), .ZN(n1115)
         );
  NAND2_X1 U1337 ( .A1(N446), .A2(n2429), .ZN(n1953) );
  NAND2_X1 U1338 ( .A1(n2452), .A2(n1953), .ZN(n1768) );
  NAND2_X1 U1339 ( .A1(N464), .A2(n2432), .ZN(n1954) );
  NAND2_X1 U1340 ( .A1(n2005), .A2(n1954), .ZN(n1762) );
  AOI222_X1 U1341 ( .A1(alu_output_EX_wire[0]), .A2(n2448), .B1(
        div_output_EX_wire[0]), .B2(n2008), .C1(mul_output_EX_wire[0]), .C2(
        n2011), .ZN(n1955) );
  AOI22_X1 U1342 ( .A1(n2440), .A2(n1207), .B1(n1955), .B2(n2445), .ZN(n1580)
         );
  INV_X1 U1343 ( .A(rs2_EX_reg[31]), .ZN(n1956) );
  AOI22_X1 U1344 ( .A1(n2441), .A2(n212), .B1(n2444), .B2(n1956), .ZN(n1122)
         );
  INV_X2 U1345 ( .A(reset), .ZN(n2475) );
  AND2_X4 U1346 ( .A1(n2480), .A2(FW_enable_2), .ZN(n2501) );
  AND2_X4 U1347 ( .A1(n2480), .A2(FW_enable_1), .ZN(n2500) );
  INV_X2 U1348 ( .A(n2480), .ZN(n2262) );
  BUF_X4 U1349 ( .A(n2262), .Z(n2429) );
  CLKBUF_X3 U1350 ( .A(n2262), .Z(n2427) );
  INV_X2 U1351 ( .A(n1247), .ZN(n2496) );
  INV_X4 U1352 ( .A(n2144), .ZN(n1488) );
  OR2_X1 U1353 ( .A1(n2418), .A2(n2165), .ZN(n1957) );
  AND2_X1 U1354 ( .A1(n1494), .A2(alu_output_EX_wire[6]), .ZN(n1958) );
  BUF_X4 U1355 ( .A(funct3_EX_reg[1]), .Z(n2474) );
  NAND2_X1 U1356 ( .A1(n2447), .A2(n1959), .ZN(n1961) );
  NAND2_X1 U1357 ( .A1(n2447), .A2(n1960), .ZN(n1962) );
  INV_X1 U1358 ( .A(n2122), .ZN(n1968) );
  NAND2_X1 U1359 ( .A1(mul_output_EX_wire[28]), .A2(n2011), .ZN(n1967) );
  NAND2_X1 U1360 ( .A1(n1967), .A2(n1968), .ZN(n1965) );
  AOI21_X1 U1361 ( .B1(n1965), .B2(n2144), .A(n1966), .ZN(n1964) );
  NAND2_X1 U1362 ( .A1(address_EX_wire[28]), .A2(n2504), .ZN(n1963) );
  NAND2_X1 U1363 ( .A1(n1963), .A2(n1964), .ZN(\_2_net_[28] ) );
  AND2_X1 U1364 ( .A1(n2293), .A2(immediate_EX_reg[31]), .ZN(n1972) );
  AOI21_X1 U1365 ( .B1(csr_rd_EX_wire[31]), .B2(n2436), .A(n1972), .ZN(n1971)
         );
  AOI21_X1 U1366 ( .B1(mul_output_EX_wire[31]), .B2(n2011), .A(n2103), .ZN(
        n1245) );
  OAI21_X1 U1367 ( .B1(n1245), .B2(n1488), .A(n1971), .ZN(n1970) );
  INV_X1 U1368 ( .A(n1970), .ZN(n1969) );
  NAND2_X1 U1369 ( .A1(n2007), .A2(N487), .ZN(n1975) );
  NAND2_X1 U1370 ( .A1(n2269), .A2(RF_source_2[24]), .ZN(n1974) );
  NAND2_X1 U1371 ( .A1(n1974), .A2(n1975), .ZN(n1973) );
  AOI21_X1 U1372 ( .B1(FW_source_2[24]), .B2(n2425), .A(n1973), .ZN(n1471) );
  AOI222_X1 U1373 ( .A1(mul_output_EX_wire[3]), .A2(n2011), .B1(
        div_output_EX_wire[3]), .B2(n2008), .C1(n2448), .C2(
        alu_output_EX_wire[3]), .ZN(n1976) );
  OAI21_X1 U1374 ( .B1(n1976), .B2(n1488), .A(n1977), .ZN(\_2_net_[3] ) );
  AOI21_X1 U1375 ( .B1(address_EX_wire[3]), .B2(n2504), .A(n1978), .ZN(n1977)
         );
  NAND2_X1 U1376 ( .A1(n2428), .A2(N454), .ZN(n1983) );
  NAND2_X1 U1377 ( .A1(n2424), .A2(RF_source_1[3]), .ZN(n1982) );
  NAND2_X1 U1378 ( .A1(n1982), .A2(n1983), .ZN(n1981) );
  AOI21_X1 U1379 ( .B1(FW_source_1[3]), .B2(n2500), .A(n1981), .ZN(n1364) );
  NAND2_X1 U1380 ( .A1(address_EX_wire[19]), .A2(n2479), .ZN(n1984) );
  NAND2_X1 U1381 ( .A1(n1984), .A2(n1985), .ZN(\_2_net_[19] ) );
  AOI21_X1 U1382 ( .B1(div_output_EX_wire[19]), .B2(n2008), .A(n1989), .ZN(
        n1987) );
  NAND2_X1 U1383 ( .A1(mul_output_EX_wire[19]), .A2(n2011), .ZN(n1988) );
  AND2_X1 U1384 ( .A1(n1986), .A2(n1488), .ZN(n1991) );
  AND2_X1 U1385 ( .A1(n1987), .A2(n1988), .ZN(n1992) );
  OR2_X1 U1386 ( .A1(n1992), .A2(n1991), .ZN(n1985) );
  NAND2_X1 U1387 ( .A1(n2007), .A2(N502), .ZN(n1995) );
  NAND2_X1 U1388 ( .A1(n2269), .A2(RF_source_2[19]), .ZN(n1994) );
  NAND2_X1 U1389 ( .A1(n1994), .A2(n1995), .ZN(n1993) );
  AOI21_X1 U1390 ( .B1(FW_source_2[19]), .B2(n2501), .A(n1993), .ZN(n1461) );
  NAND2_X1 U1391 ( .A1(div_output_EX_wire[29]), .A2(n2008), .ZN(n2001) );
  NAND2_X1 U1392 ( .A1(n2001), .A2(n2002), .ZN(n2000) );
  AOI21_X1 U1393 ( .B1(mul_output_EX_wire[29]), .B2(n2011), .A(n2000), .ZN(
        n1996) );
  OAI21_X1 U1394 ( .B1(n1996), .B2(n1488), .A(n1997), .ZN(\_2_net_[29] ) );
  AOI21_X1 U1395 ( .B1(address_EX_wire[29]), .B2(n2479), .A(n1998), .ZN(n1997)
         );
  NOR2_X1 U1396 ( .A1(n2453), .A2(n1354), .ZN(n1246) );
  BUF_X1 U1397 ( .A(n2266), .Z(n2268) );
  BUF_X2 U1398 ( .A(n2266), .Z(n2423) );
  BUF_X2 U1399 ( .A(n2267), .Z(n2004) );
  BUF_X1 U1400 ( .A(n2426), .Z(n2433) );
  BUF_X1 U1401 ( .A(n2426), .Z(n2430) );
  INV_X2 U1402 ( .A(n2453), .ZN(n2005) );
  BUF_X1 U1403 ( .A(n2262), .Z(n2432) );
  BUF_X2 U1404 ( .A(n2499), .Z(n2006) );
  BUF_X1 U1405 ( .A(n2501), .Z(n2425) );
  BUF_X1 U1406 ( .A(n2426), .Z(n2434) );
  BUF_X1 U1407 ( .A(n2262), .Z(n2431) );
  BUF_X1 U1408 ( .A(n2500), .Z(n2422) );
  BUF_X1 U1409 ( .A(n2426), .Z(n2428) );
  BUF_X2 U1410 ( .A(n2426), .Z(n2007) );
  BUF_X1 U1411 ( .A(n2444), .Z(n2447) );
  BUF_X1 U1412 ( .A(n2502), .Z(n2435) );
  CLKBUF_X3 U1413 ( .A(n2503), .Z(n2011) );
  BUF_X4 U1414 ( .A(n2504), .Z(n2479) );
  BUF_X2 U1415 ( .A(n2502), .Z(n2008) );
  BUF_X2 U1416 ( .A(n203), .Z(n2013) );
  BUF_X2 U1417 ( .A(n207), .Z(n2014) );
  BUF_X2 U1418 ( .A(n205), .Z(n2009) );
  INV_X1 U1419 ( .A(n1165), .ZN(n2154) );
  BUF_X2 U1420 ( .A(n2456), .Z(n2468) );
  BUF_X2 U1421 ( .A(n2456), .Z(n2470) );
  BUF_X2 U1422 ( .A(n2455), .Z(n2469) );
  BUF_X1 U1423 ( .A(n2498), .Z(n2419) );
  BUF_X1 U1424 ( .A(n2498), .Z(n2420) );
  BUF_X1 U1425 ( .A(n2499), .Z(n2421) );
  BUF_X1 U1426 ( .A(n2267), .Z(n2269) );
  INV_X1 U1427 ( .A(n2454), .ZN(n2451) );
  INV_X1 U1428 ( .A(n2454), .ZN(n2449) );
  INV_X1 U1429 ( .A(n2454), .ZN(n2452) );
  INV_X1 U1430 ( .A(n2454), .ZN(n2450) );
  INV_X1 U1431 ( .A(n2483), .ZN(n2498) );
  INV_X1 U1432 ( .A(n2480), .ZN(n2426) );
  OR2_X1 U1433 ( .A1(n2509), .A2(n1485), .ZN(n1354) );
  INV_X1 U1434 ( .A(n2444), .ZN(n2441) );
  INV_X1 U1435 ( .A(n2444), .ZN(n2442) );
  INV_X1 U1436 ( .A(n2444), .ZN(n2440) );
  INV_X1 U1437 ( .A(n2444), .ZN(n2439) );
  INV_X1 U1438 ( .A(n2444), .ZN(n2437) );
  INV_X1 U1439 ( .A(n2444), .ZN(n2438) );
  BUF_X2 U1440 ( .A(n2444), .Z(n2446) );
  INV_X1 U1441 ( .A(n2444), .ZN(n2443) );
  BUF_X2 U1442 ( .A(n2444), .Z(n2445) );
  NAND2_X1 U1443 ( .A1(n2035), .A2(n2036), .ZN(n2034) );
  NAND2_X1 U1444 ( .A1(n2130), .A2(n2131), .ZN(n2129) );
  NAND2_X1 U1445 ( .A1(csr_rd_EX_wire[18]), .A2(n2436), .ZN(n2130) );
  NAND2_X1 U1446 ( .A1(n2472), .A2(n2473), .ZN(n2509) );
  NAND2_X1 U1447 ( .A1(csr_rd_EX_wire[25]), .A2(n2436), .ZN(n2035) );
  AOI21_X1 U1448 ( .B1(csr_rd_EX_wire[22]), .B2(n2436), .A(n2105), .ZN(n2104)
         );
  OR2_X1 U1449 ( .A1(n2418), .A2(n2159), .ZN(n2036) );
  INV_X1 U1450 ( .A(mul_busy_EX_wire), .ZN(n2473) );
  NOR2_X1 U1451 ( .A1(n1494), .A2(n1169), .ZN(n2502) );
  NOR2_X1 U1452 ( .A1(n2418), .A2(n2166), .ZN(n2105) );
  OR2_X1 U1453 ( .A1(n2418), .A2(n2160), .ZN(n2131) );
  INV_X1 U1454 ( .A(n2293), .ZN(n2418) );
  AND2_X1 U1455 ( .A1(n2477), .A2(n2414), .ZN(n2293) );
  INV_X2 U1456 ( .A(n2156), .ZN(n2436) );
  BUF_X1 U1457 ( .A(n596), .Z(n2471) );
  OR4_X1 U1458 ( .A1(n1559), .A2(n1166), .A3(n2072), .A4(n1165), .ZN(n2156) );
  CLKBUF_X1 U1459 ( .A(rs1_EX_reg[0]), .Z(n2062) );
  AND4_X1 U1460 ( .A1(n1210), .A2(n1209), .A3(n1208), .A4(n1565), .ZN(n205) );
  BUF_X1 U1461 ( .A(opcode_EX_reg[3]), .Z(n2077) );
  CLKBUF_X1 U1462 ( .A(reset), .Z(n2476) );
  NAND2_X1 U1463 ( .A1(mul_output_EX_wire[6]), .A2(n2011), .ZN(n2015) );
  AND2_X1 U1464 ( .A1(n2015), .A2(n2016), .ZN(n1220) );
  AOI21_X1 U1465 ( .B1(div_output_EX_wire[6]), .B2(n2435), .A(n1958), .ZN(
        n2016) );
  NAND2_X1 U1466 ( .A1(n2427), .A2(N541), .ZN(n2019) );
  NAND2_X1 U1467 ( .A1(n2004), .A2(RF_source_2[6]), .ZN(n2018) );
  NAND2_X1 U1468 ( .A1(n2018), .A2(n2019), .ZN(n2017) );
  AOI21_X1 U1469 ( .B1(FW_source_2[6]), .B2(n2501), .A(n2017), .ZN(n1435) );
  NAND2_X1 U1470 ( .A1(n2427), .A2(N445), .ZN(n2022) );
  NAND2_X1 U1471 ( .A1(n2423), .A2(RF_source_1[6]), .ZN(n2021) );
  NAND2_X1 U1472 ( .A1(n2021), .A2(n2022), .ZN(n2020) );
  AOI21_X1 U1473 ( .B1(FW_source_1[6]), .B2(n2500), .A(n2020), .ZN(n1370) );
  OR2_X1 U1474 ( .A1(n2418), .A2(n2171), .ZN(n2026) );
  NAND2_X1 U1475 ( .A1(csr_rd_EX_wire[10]), .A2(n2436), .ZN(n2025) );
  NAND2_X1 U1476 ( .A1(n2025), .A2(n2026), .ZN(n2024) );
  AOI21_X1 U1477 ( .B1(address_EX_wire[10]), .B2(n2479), .A(n2024), .ZN(n2023)
         );
  NAND2_X1 U1478 ( .A1(n2427), .A2(N529), .ZN(n2030) );
  NAND2_X1 U1479 ( .A1(n2004), .A2(RF_source_2[10]), .ZN(n2029) );
  NAND2_X1 U1480 ( .A1(n2029), .A2(n2030), .ZN(n2028) );
  AND2_X1 U1481 ( .A1(div_output_EX_wire[25]), .A2(n2008), .ZN(n2292) );
  NOR2_X1 U1482 ( .A1(n2292), .A2(n2291), .ZN(n2037) );
  NAND2_X1 U1483 ( .A1(n2037), .A2(n2038), .ZN(n2033) );
  NAND2_X1 U1484 ( .A1(mul_output_EX_wire[25]), .A2(n2011), .ZN(n2038) );
  AOI21_X1 U1485 ( .B1(n2033), .B2(n2144), .A(n2034), .ZN(n2031) );
  NAND2_X1 U1486 ( .A1(n2031), .A2(n2032), .ZN(\_2_net_[25] ) );
  NAND2_X1 U1487 ( .A1(address_EX_wire[25]), .A2(n2479), .ZN(n2032) );
  NAND2_X1 U1488 ( .A1(n2007), .A2(N475), .ZN(n2041) );
  NAND2_X1 U1489 ( .A1(n2004), .A2(RF_source_2[28]), .ZN(n2040) );
  NAND2_X1 U1490 ( .A1(n2040), .A2(n2041), .ZN(n2039) );
  AOI21_X1 U1491 ( .B1(FW_source_2[28]), .B2(n2425), .A(n2039), .ZN(n2505) );
  AOI222_X2 U1492 ( .A1(mul_output_EX_wire[5]), .A2(n2011), .B1(
        div_output_EX_wire[5]), .B2(n2435), .C1(n1494), .C2(
        alu_output_EX_wire[5]), .ZN(n1219) );
  NAND2_X1 U1493 ( .A1(n2293), .A2(immediate_EX_reg[5]), .ZN(n2045) );
  NAND2_X1 U1494 ( .A1(csr_rd_EX_wire[5]), .A2(n2436), .ZN(n2044) );
  NAND2_X1 U1495 ( .A1(n2044), .A2(n2045), .ZN(n2043) );
  AOI21_X1 U1496 ( .B1(address_EX_wire[5]), .B2(n2479), .A(n2043), .ZN(n2042)
         );
  OAI21_X1 U1497 ( .B1(n1219), .B2(n1488), .A(n2042), .ZN(\_2_net_[5] ) );
  NAND2_X1 U1498 ( .A1(n2427), .A2(N544), .ZN(n2048) );
  NAND2_X1 U1499 ( .A1(n2004), .A2(RF_source_2[5]), .ZN(n2047) );
  NAND2_X1 U1500 ( .A1(n2047), .A2(n2048), .ZN(n2046) );
  AOI21_X1 U1501 ( .B1(FW_source_2[5]), .B2(n2501), .A(n2046), .ZN(n1433) );
  NAND2_X1 U1502 ( .A1(n2427), .A2(N448), .ZN(n2051) );
  NAND2_X1 U1503 ( .A1(n2424), .A2(RF_source_1[5]), .ZN(n2050) );
  NAND2_X1 U1504 ( .A1(n2050), .A2(n2051), .ZN(n2049) );
  AOI21_X1 U1505 ( .B1(FW_source_1[5]), .B2(n2500), .A(n2049), .ZN(n1368) );
  AOI222_X1 U1506 ( .A1(n2448), .A2(alu_output_EX_wire[27]), .B1(n2008), .B2(
        div_output_EX_wire[27]), .C1(mul_output_EX_wire[27]), .C2(n2011), .ZN(
        n2052) );
  INV_X1 U1507 ( .A(n2012), .ZN(n2472) );
  AOI21_X1 U1508 ( .B1(n2444), .B2(n1485), .A(n2413), .ZN(n2056) );
  AOI222_X1 U1509 ( .A1(n2448), .A2(alu_output_EX_wire[15]), .B1(n2435), .B2(
        div_output_EX_wire[15]), .C1(mul_output_EX_wire[15]), .C2(n2011), .ZN(
        n2057) );
  AOI222_X1 U1510 ( .A1(n2448), .A2(alu_output_EX_wire[16]), .B1(n2435), .B2(
        div_output_EX_wire[16]), .C1(mul_output_EX_wire[16]), .C2(n2011), .ZN(
        n2060) );
  AOI222_X1 U1511 ( .A1(n2448), .A2(alu_output_EX_wire[2]), .B1(n2008), .B2(
        div_output_EX_wire[2]), .C1(mul_output_EX_wire[2]), .C2(n2011), .ZN(
        n2061) );
  NAND2_X1 U1512 ( .A1(div_output_EX_wire[31]), .A2(n2008), .ZN(n2063) );
  NAND2_X1 U1513 ( .A1(n2063), .A2(n2064), .ZN(n2103) );
  NAND2_X1 U1514 ( .A1(n2007), .A2(N511), .ZN(n2067) );
  NAND2_X1 U1515 ( .A1(n2269), .A2(RF_source_2[16]), .ZN(n2066) );
  NAND2_X1 U1516 ( .A1(n2066), .A2(n2067), .ZN(n2065) );
  AOI21_X1 U1517 ( .B1(FW_source_2[16]), .B2(n2501), .A(n2065), .ZN(n1455) );
  AOI222_X1 U1518 ( .A1(n1494), .A2(alu_output_EX_wire[7]), .B1(n2435), .B2(
        div_output_EX_wire[7]), .C1(mul_output_EX_wire[7]), .C2(n2011), .ZN(
        n2068) );
  AOI222_X1 U1519 ( .A1(n1494), .A2(alu_output_EX_wire[13]), .B1(n2435), .B2(
        div_output_EX_wire[13]), .C1(mul_output_EX_wire[13]), .C2(n2011), .ZN(
        n2069) );
  AOI222_X1 U1520 ( .A1(n2448), .A2(alu_output_EX_wire[26]), .B1(n2008), .B2(
        div_output_EX_wire[26]), .C1(mul_output_EX_wire[26]), .C2(n2011), .ZN(
        n2070) );
  AOI222_X1 U1521 ( .A1(n2448), .A2(alu_output_EX_wire[19]), .B1(
        div_output_EX_wire[19]), .B2(n2008), .C1(mul_output_EX_wire[19]), .C2(
        n2011), .ZN(n2071) );
  INV_X1 U1522 ( .A(n1168), .ZN(n2072) );
  AOI21_X1 U1523 ( .B1(mul_output_EX_wire[31]), .B2(n2011), .A(n1909), .ZN(
        n2073) );
  AOI21_X1 U1524 ( .B1(mul_output_EX_wire[28]), .B2(n2011), .A(n2122), .ZN(
        n2074) );
  AOI21_X1 U1525 ( .B1(mul_output_EX_wire[20]), .B2(n2011), .A(n2229), .ZN(
        n2075) );
  NAND2_X1 U1526 ( .A1(n2418), .A2(n2156), .ZN(n2079) );
  NOR2_X1 U1527 ( .A1(n2079), .A2(n2479), .ZN(n2144) );
  INV_X1 U1528 ( .A(address_EX_wire[22]), .ZN(n2080) );
  INV_X1 U1529 ( .A(n2479), .ZN(n2081) );
  AOI21_X1 U1530 ( .B1(n2444), .B2(n1485), .A(n2413), .ZN(n1285) );
  BUF_X1 U1531 ( .A(address_EX_wire[25]), .Z(n2086) );
  CLKBUF_X3 U1532 ( .A(n1246), .Z(n2456) );
  CLKBUF_X3 U1533 ( .A(n1246), .Z(n2455) );
  CLKBUF_X3 U1534 ( .A(n2455), .Z(n2457) );
  CLKBUF_X3 U1535 ( .A(n2456), .Z(n2467) );
  CLKBUF_X3 U1536 ( .A(n2456), .Z(n2466) );
  CLKBUF_X3 U1537 ( .A(n2456), .Z(n2151) );
  CLKBUF_X3 U1538 ( .A(n2456), .Z(n2462) );
  CLKBUF_X3 U1539 ( .A(n2456), .Z(n2465) );
  AOI21_X1 U1540 ( .B1(mul_output_EX_wire[23]), .B2(n2011), .A(n2135), .ZN(
        n2087) );
  BUF_X1 U1541 ( .A(address_EX_wire[19]), .Z(n2090) );
  AOI21_X1 U1542 ( .B1(mul_output_EX_wire[24]), .B2(n2011), .A(n2100), .ZN(
        n2091) );
  BUF_X1 U1543 ( .A(address_EX_wire[21]), .Z(n2092) );
  OR2_X1 U1544 ( .A1(n1234), .A2(n1488), .ZN(n2094) );
  NAND2_X1 U1545 ( .A1(n2094), .A2(n2306), .ZN(\_2_net_[20] ) );
  BUF_X1 U1546 ( .A(address_EX_wire[22]), .Z(n2099) );
  NAND2_X1 U1547 ( .A1(div_output_EX_wire[24]), .A2(n2008), .ZN(n2101) );
  NAND2_X1 U1548 ( .A1(n2101), .A2(n2102), .ZN(n2100) );
  OR2_X1 U1549 ( .A1(n2418), .A2(n2163), .ZN(n2109) );
  NAND2_X1 U1550 ( .A1(csr_rd_EX_wire[26]), .A2(n2436), .ZN(n2108) );
  NAND2_X1 U1551 ( .A1(n2108), .A2(n2109), .ZN(n2107) );
  AOI21_X1 U1552 ( .B1(address_EX_wire[26]), .B2(n2479), .A(n2107), .ZN(n2106)
         );
  OAI21_X1 U1553 ( .B1(n1240), .B2(n1488), .A(n2106), .ZN(\_2_net_[26] ) );
  NAND2_X1 U1554 ( .A1(n2007), .A2(N481), .ZN(n2112) );
  NAND2_X1 U1555 ( .A1(n2269), .A2(RF_source_2[26]), .ZN(n2111) );
  NAND2_X1 U1556 ( .A1(n2111), .A2(n2112), .ZN(n2110) );
  AOI21_X1 U1557 ( .B1(FW_source_2[26]), .B2(n2425), .A(n2110), .ZN(n1475) );
  NAND2_X1 U1558 ( .A1(n2262), .A2(N385), .ZN(n2115) );
  NAND2_X1 U1559 ( .A1(n2424), .A2(RF_source_1[26]), .ZN(n2114) );
  NAND2_X1 U1560 ( .A1(n2114), .A2(n2115), .ZN(n2113) );
  AOI21_X1 U1561 ( .B1(FW_source_1[26]), .B2(n2422), .A(n2113), .ZN(n1410) );
  INV_X4 U1562 ( .A(n2509), .ZN(n2444) );
  NAND2_X1 U1563 ( .A1(n2125), .A2(n2127), .ZN(\_2_net_[16] ) );
  OR2_X2 U1564 ( .A1(jump_branch_enable_EX_wire), .A2(n2444), .ZN(n2480) );
  NOR2_X1 U1565 ( .A1(n2262), .A2(FW_enable_1), .ZN(n2266) );
  NAND2_X1 U1566 ( .A1(n2427), .A2(N472), .ZN(n2118) );
  NAND2_X1 U1567 ( .A1(n2004), .A2(RF_source_2[29]), .ZN(n2117) );
  NAND2_X1 U1568 ( .A1(n2117), .A2(n2118), .ZN(n2116) );
  AOI21_X1 U1569 ( .B1(FW_source_2[29]), .B2(n2425), .A(n2116), .ZN(n1481) );
  AND2_X1 U1570 ( .A1(n2262), .A2(N376), .ZN(n2121) );
  AND2_X1 U1571 ( .A1(n2268), .A2(RF_source_1[29]), .ZN(n2120) );
  OR2_X1 U1572 ( .A1(n2120), .A2(n2121), .ZN(n2119) );
  AOI21_X1 U1573 ( .B1(FW_source_1[29]), .B2(n2500), .A(n2119), .ZN(n1416) );
  NAND2_X1 U1574 ( .A1(div_output_EX_wire[28]), .A2(n2008), .ZN(n2123) );
  NAND2_X1 U1575 ( .A1(n2123), .A2(n2124), .ZN(n2122) );
  OR2_X1 U1576 ( .A1(n1230), .A2(n1488), .ZN(n2127) );
  AOI21_X1 U1577 ( .B1(n2010), .B2(n2479), .A(n2126), .ZN(n2125) );
  AOI21_X1 U1578 ( .B1(address_EX_wire[18]), .B2(n2479), .A(n2129), .ZN(n2128)
         );
  OAI21_X1 U1579 ( .B1(n1232), .B2(n1488), .A(n2128), .ZN(\_2_net_[18] ) );
  NAND2_X1 U1580 ( .A1(n2007), .A2(N505), .ZN(n2134) );
  NAND2_X1 U1581 ( .A1(n2269), .A2(RF_source_2[18]), .ZN(n2133) );
  NAND2_X1 U1582 ( .A1(n2133), .A2(n2134), .ZN(n2132) );
  AOI21_X1 U1583 ( .B1(FW_source_2[18]), .B2(n2425), .A(n2132), .ZN(n1459) );
  NAND2_X1 U1584 ( .A1(div_output_EX_wire[23]), .A2(n2008), .ZN(n2136) );
  AOI21_X1 U1585 ( .B1(FW_source_2[22]), .B2(n2425), .A(n2138), .ZN(n1467) );
  AOI21_X1 U1586 ( .B1(FW_source_1[22]), .B2(n2422), .A(n2141), .ZN(n1402) );
  NAND2_X1 U1587 ( .A1(n2429), .A2(N493), .ZN(n2140) );
  NAND2_X1 U1588 ( .A1(n2269), .A2(RF_source_2[22]), .ZN(n2139) );
  NAND2_X1 U1589 ( .A1(n2139), .A2(n2140), .ZN(n2138) );
  NAND2_X1 U1590 ( .A1(n2426), .A2(N397), .ZN(n2143) );
  NAND2_X1 U1591 ( .A1(n2423), .A2(RF_source_1[22]), .ZN(n2142) );
  NAND2_X1 U1592 ( .A1(n2142), .A2(n2143), .ZN(n2141) );
  NAND2_X1 U1593 ( .A1(n2007), .A2(N484), .ZN(n2147) );
  NAND2_X1 U1594 ( .A1(n2269), .A2(RF_source_2[25]), .ZN(n2146) );
  NAND2_X1 U1595 ( .A1(n2146), .A2(n2147), .ZN(n2145) );
  AOI21_X1 U1596 ( .B1(FW_source_2[25]), .B2(n2425), .A(n2145), .ZN(n1473) );
  NAND2_X1 U1597 ( .A1(n2262), .A2(N379), .ZN(n2150) );
  NAND2_X1 U1598 ( .A1(n2424), .A2(RF_source_1[28]), .ZN(n2149) );
  NAND2_X1 U1599 ( .A1(n2149), .A2(n2150), .ZN(n2148) );
  AOI21_X1 U1600 ( .B1(FW_source_1[28]), .B2(n2422), .A(n2148), .ZN(n2506) );
  AND2_X1 U1601 ( .A1(n2446), .A2(n2077), .ZN(N655) );
  NOR4_X1 U1602 ( .A1(n2072), .A2(n2154), .A3(n2077), .A4(n2414), .ZN(n1569)
         );
  OR3_X1 U1603 ( .A1(n1564), .A2(n2077), .A3(n1167), .ZN(n1559) );
  CLKBUF_X3 U1604 ( .A(n2456), .Z(n2463) );
  CLKBUF_X3 U1605 ( .A(n2456), .Z(n2464) );
  CLKBUF_X3 U1606 ( .A(n2455), .Z(n2152) );
  CLKBUF_X3 U1607 ( .A(n2455), .Z(n2153) );
  BUF_X2 U1608 ( .A(opcode_EX_reg[5]), .Z(n2414) );
  CLKBUF_X3 U1609 ( .A(n2455), .Z(n2461) );
  CLKBUF_X3 U1610 ( .A(n2455), .Z(n2458) );
  CLKBUF_X3 U1611 ( .A(n2455), .Z(n2459) );
  CLKBUF_X3 U1612 ( .A(n2455), .Z(n2460) );
  INV_X1 U1613 ( .A(n1285), .ZN(n2453) );
  NOR2_X4 U1614 ( .A1(opcode_MW_reg[6]), .A2(n67), .ZN(n204) );
  OR2_X2 U1615 ( .A1(n2413), .A2(n2417), .ZN(n1247) );
  BUF_X1 U1616 ( .A(n2266), .Z(n2424) );
  NOR2_X1 U1617 ( .A1(n2426), .A2(FW_enable_2), .ZN(n2267) );
  BUF_X2 U1618 ( .A(jump_branch_enable_EX_wire), .Z(n2413) );
  BUF_X2 U1619 ( .A(n1494), .Z(n2448) );
  NOR2_X4 U1620 ( .A1(opcode_MW_reg[5]), .A2(n66), .ZN(n201) );
  NOR2_X4 U1621 ( .A1(n1208), .A2(n66), .ZN(n202) );
  OAI211_X2 U1622 ( .C1(n1208), .C2(n80), .A(n79), .B(n78), .ZN(n596) );
  NOR4_X1 U1623 ( .A1(n790), .A2(n1210), .A3(n1208), .A4(opcode_MW_reg[4]), 
        .ZN(n207) );
  AOI22_X1 U1624 ( .A1(address_EX_wire[29]), .A2(n2006), .B1(n2419), .B2(
        pc_FD_reg[29]), .ZN(n2226) );
  AOI22_X1 U1625 ( .A1(n2006), .A2(address_EX_wire[30]), .B1(n2419), .B2(
        pc_FD_reg[30]), .ZN(n2224) );
  AOI222_X1 U1626 ( .A1(n2006), .A2(n2097), .B1(n2419), .B2(pc_FD_reg[24]), 
        .C1(n2496), .C2(next_pc_FD_wire[24]), .ZN(n2487) );
  NAND2_X1 U1627 ( .A1(n2316), .A2(n2213), .ZN(n2315) );
  NAND2_X1 U1628 ( .A1(csr_rd_EX_wire[8]), .A2(n2436), .ZN(n2316) );
  AOI21_X1 U1629 ( .B1(mul_output_EX_wire[8]), .B2(n2011), .A(n2235), .ZN(
        n1222) );
  NAND2_X1 U1630 ( .A1(n1494), .A2(alu_output_EX_wire[8]), .ZN(n2237) );
  NAND2_X1 U1631 ( .A1(n2319), .A2(n2214), .ZN(n2318) );
  NAND2_X1 U1632 ( .A1(csr_rd_EX_wire[11]), .A2(n2436), .ZN(n2319) );
  AOI21_X1 U1633 ( .B1(mul_output_EX_wire[11]), .B2(n2011), .A(n2238), .ZN(
        n1225) );
  NAND2_X1 U1634 ( .A1(n1494), .A2(alu_output_EX_wire[11]), .ZN(n2240) );
  OR2_X1 U1635 ( .A1(n2413), .A2(n2482), .ZN(n2483) );
  NAND2_X1 U1636 ( .A1(n1354), .A2(n2475), .ZN(n2482) );
  NOR2_X1 U1637 ( .A1(n2481), .A2(reset), .ZN(n2499) );
  INV_X1 U1638 ( .A(n2413), .ZN(n2481) );
  AOI21_X1 U1639 ( .B1(address_EX_wire[0]), .B2(n2504), .A(n2251), .ZN(n2250)
         );
  NAND2_X1 U1640 ( .A1(n2252), .A2(n2253), .ZN(n2251) );
  NAND2_X1 U1641 ( .A1(n2293), .A2(immediate_EX_reg[0]), .ZN(n2253) );
  NAND2_X1 U1642 ( .A1(csr_rd_EX_wire[0]), .A2(n2436), .ZN(n2252) );
  AOI21_X1 U1643 ( .B1(address_EX_wire[1]), .B2(n2504), .A(n2255), .ZN(n2254)
         );
  NAND2_X1 U1644 ( .A1(n2256), .A2(n2257), .ZN(n2255) );
  NAND2_X1 U1645 ( .A1(n2293), .A2(immediate_EX_reg[1]), .ZN(n2257) );
  NAND2_X1 U1646 ( .A1(csr_rd_EX_wire[1]), .A2(n2436), .ZN(n2256) );
  AOI21_X1 U1647 ( .B1(address_EX_wire[2]), .B2(n2504), .A(n2259), .ZN(n2258)
         );
  NAND2_X1 U1648 ( .A1(n2260), .A2(n2261), .ZN(n2259) );
  NAND2_X1 U1649 ( .A1(n2293), .A2(immediate_EX_reg[2]), .ZN(n2261) );
  NAND2_X1 U1650 ( .A1(csr_rd_EX_wire[2]), .A2(n2436), .ZN(n2260) );
  NAND2_X1 U1651 ( .A1(n2334), .A2(n2218), .ZN(n2333) );
  NAND2_X1 U1652 ( .A1(csr_rd_EX_wire[17]), .A2(n2436), .ZN(n2334) );
  AOI21_X1 U1653 ( .B1(mul_output_EX_wire[17]), .B2(n2011), .A(n2247), .ZN(
        n1231) );
  NAND2_X1 U1654 ( .A1(n2448), .A2(alu_output_EX_wire[17]), .ZN(n2249) );
  NAND2_X1 U1655 ( .A1(n2296), .A2(n2212), .ZN(n2295) );
  NAND2_X1 U1656 ( .A1(csr_rd_EX_wire[7]), .A2(n2436), .ZN(n2296) );
  AOI222_X1 U1657 ( .A1(n1494), .A2(alu_output_EX_wire[7]), .B1(n2435), .B2(
        div_output_EX_wire[7]), .C1(mul_output_EX_wire[7]), .C2(n2011), .ZN(
        n1221) );
  NAND2_X1 U1658 ( .A1(n2322), .A2(n2215), .ZN(n2321) );
  NAND2_X1 U1659 ( .A1(csr_rd_EX_wire[12]), .A2(n2436), .ZN(n2322) );
  AOI21_X1 U1660 ( .B1(mul_output_EX_wire[12]), .B2(n2011), .A(n2241), .ZN(
        n1226) );
  NAND2_X1 U1661 ( .A1(n1494), .A2(alu_output_EX_wire[12]), .ZN(n2243) );
  NAND2_X1 U1662 ( .A1(n2429), .A2(N553), .ZN(n2284) );
  NAND2_X1 U1663 ( .A1(n2429), .A2(N460), .ZN(n2281) );
  NAND2_X1 U1664 ( .A1(n2429), .A2(N463), .ZN(n2275) );
  NAND2_X1 U1665 ( .A1(n2429), .A2(N559), .ZN(n2272) );
  NAND2_X1 U1666 ( .A1(n2429), .A2(N556), .ZN(n2278) );
  NAND2_X1 U1667 ( .A1(n2429), .A2(N457), .ZN(n2287) );
  NAND2_X1 U1668 ( .A1(n2429), .A2(N550), .ZN(n2290) );
  NAND2_X1 U1669 ( .A1(n2426), .A2(N382), .ZN(n2355) );
  NAND2_X1 U1670 ( .A1(n2423), .A2(RF_source_1[27]), .ZN(n2354) );
  NAND2_X1 U1671 ( .A1(n2313), .A2(n2221), .ZN(n2312) );
  NAND2_X1 U1672 ( .A1(csr_rd_EX_wire[27]), .A2(n2436), .ZN(n2313) );
  AOI222_X1 U1673 ( .A1(n2448), .A2(alu_output_EX_wire[27]), .B1(n2008), .B2(
        div_output_EX_wire[27]), .C1(mul_output_EX_wire[27]), .C2(n2011), .ZN(
        n1241) );
  NAND2_X1 U1674 ( .A1(n2427), .A2(N535), .ZN(n2391) );
  NAND2_X1 U1675 ( .A1(n2004), .A2(RF_source_2[8]), .ZN(n2390) );
  NAND2_X1 U1676 ( .A1(n2427), .A2(N523), .ZN(n2397) );
  NAND2_X1 U1677 ( .A1(n2004), .A2(RF_source_2[12]), .ZN(n2396) );
  NAND2_X1 U1678 ( .A1(n2428), .A2(N439), .ZN(n2394) );
  NAND2_X1 U1679 ( .A1(n2424), .A2(RF_source_1[8]), .ZN(n2393) );
  NAND2_X1 U1680 ( .A1(n2007), .A2(N412), .ZN(n2388) );
  NAND2_X1 U1681 ( .A1(n2423), .A2(RF_source_1[17]), .ZN(n2387) );
  NAND2_X1 U1682 ( .A1(n2427), .A2(N508), .ZN(n2385) );
  NAND2_X1 U1683 ( .A1(n2004), .A2(RF_source_2[17]), .ZN(n2384) );
  NAND2_X1 U1684 ( .A1(n2427), .A2(N427), .ZN(n2400) );
  NAND2_X1 U1685 ( .A1(n2268), .A2(RF_source_1[12]), .ZN(n2399) );
  NAND2_X1 U1686 ( .A1(n2428), .A2(N430), .ZN(n2412) );
  NAND2_X1 U1687 ( .A1(n2268), .A2(RF_source_1[11]), .ZN(n2411) );
  NAND2_X1 U1688 ( .A1(n2427), .A2(N442), .ZN(n2406) );
  NAND2_X1 U1689 ( .A1(n2268), .A2(RF_source_1[7]), .ZN(n2405) );
  NAND2_X1 U1690 ( .A1(n2427), .A2(N538), .ZN(n2403) );
  NAND2_X1 U1691 ( .A1(n2004), .A2(RF_source_2[7]), .ZN(n2402) );
  NAND2_X1 U1692 ( .A1(n2427), .A2(N526), .ZN(n2409) );
  NAND2_X1 U1693 ( .A1(n2004), .A2(RF_source_2[11]), .ZN(n2408) );
  NAND2_X1 U1694 ( .A1(n2007), .A2(N373), .ZN(n2340) );
  NAND2_X1 U1695 ( .A1(n2424), .A2(RF_source_1[30]), .ZN(n2339) );
  NAND2_X1 U1696 ( .A1(n2429), .A2(N469), .ZN(n2265) );
  NAND2_X1 U1697 ( .A1(n2302), .A2(n2219), .ZN(n2301) );
  NAND2_X1 U1698 ( .A1(csr_rd_EX_wire[30]), .A2(n2436), .ZN(n2302) );
  NAND2_X1 U1699 ( .A1(n2262), .A2(N406), .ZN(n2337) );
  NAND2_X1 U1700 ( .A1(n2423), .A2(RF_source_1[19]), .ZN(n2336) );
  NAND2_X1 U1701 ( .A1(n2429), .A2(N418), .ZN(n2382) );
  NAND2_X1 U1702 ( .A1(n2268), .A2(RF_source_1[15]), .ZN(n2381) );
  NAND2_X1 U1703 ( .A1(n2007), .A2(N478), .ZN(n2358) );
  NAND2_X1 U1704 ( .A1(n2269), .A2(RF_source_2[27]), .ZN(n2357) );
  NAND2_X1 U1705 ( .A1(n2426), .A2(N400), .ZN(n2349) );
  NAND2_X1 U1706 ( .A1(n2424), .A2(RF_source_1[21]), .ZN(n2348) );
  NAND2_X1 U1707 ( .A1(n2007), .A2(N496), .ZN(n2352) );
  NAND2_X1 U1708 ( .A1(n2269), .A2(RF_source_2[21]), .ZN(n2351) );
  NAND2_X1 U1709 ( .A1(n2310), .A2(n2220), .ZN(n2309) );
  NAND2_X1 U1710 ( .A1(csr_rd_EX_wire[21]), .A2(n2436), .ZN(n2310) );
  NAND2_X1 U1711 ( .A1(n2448), .A2(alu_output_EX_wire[21]), .ZN(n2234) );
  NAND2_X1 U1712 ( .A1(n2428), .A2(N433), .ZN(n2364) );
  NAND2_X1 U1713 ( .A1(n2423), .A2(RF_source_1[10]), .ZN(n2363) );
  NAND2_X1 U1714 ( .A1(n2007), .A2(N517), .ZN(n2373) );
  NAND2_X1 U1715 ( .A1(n2004), .A2(RF_source_2[14]), .ZN(n2372) );
  NAND2_X1 U1716 ( .A1(n2427), .A2(N421), .ZN(n2376) );
  NAND2_X1 U1717 ( .A1(n2423), .A2(RF_source_1[14]), .ZN(n2375) );
  NAND2_X1 U1718 ( .A1(n2328), .A2(n2216), .ZN(n2327) );
  NAND2_X1 U1719 ( .A1(csr_rd_EX_wire[14]), .A2(n2436), .ZN(n2328) );
  AOI21_X1 U1720 ( .B1(mul_output_EX_wire[14]), .B2(n2011), .A(n2244), .ZN(
        n1228) );
  NAND2_X1 U1721 ( .A1(n1494), .A2(alu_output_EX_wire[14]), .ZN(n2246) );
  NAND2_X1 U1722 ( .A1(n2427), .A2(N424), .ZN(n2370) );
  NAND2_X1 U1723 ( .A1(n2423), .A2(RF_source_1[13]), .ZN(n2369) );
  NAND2_X1 U1724 ( .A1(n2429), .A2(N520), .ZN(n2367) );
  NAND2_X1 U1725 ( .A1(n2004), .A2(RF_source_2[13]), .ZN(n2366) );
  AOI222_X1 U1726 ( .A1(n1494), .A2(alu_output_EX_wire[13]), .B1(n2435), .B2(
        div_output_EX_wire[13]), .C1(mul_output_EX_wire[13]), .C2(n2011), .ZN(
        n1227) );
  NAND2_X1 U1727 ( .A1(n2429), .A2(N409), .ZN(n2361) );
  NAND2_X1 U1728 ( .A1(n2268), .A2(RF_source_1[18]), .ZN(n2360) );
  NAND2_X1 U1729 ( .A1(n2007), .A2(N514), .ZN(n2379) );
  NAND2_X1 U1730 ( .A1(n2269), .A2(RF_source_2[15]), .ZN(n2378) );
  NAND2_X1 U1731 ( .A1(n2331), .A2(n2217), .ZN(n2330) );
  NAND2_X1 U1732 ( .A1(csr_rd_EX_wire[15]), .A2(n2436), .ZN(n2331) );
  AOI222_X1 U1733 ( .A1(n2448), .A2(alu_output_EX_wire[15]), .B1(n2435), .B2(
        div_output_EX_wire[15]), .C1(mul_output_EX_wire[15]), .C2(n2011), .ZN(
        n1229) );
  NAND2_X1 U1734 ( .A1(n2007), .A2(N415), .ZN(n2305) );
  NAND2_X1 U1735 ( .A1(n2268), .A2(RF_source_1[16]), .ZN(n2304) );
  AOI222_X1 U1736 ( .A1(n2448), .A2(alu_output_EX_wire[16]), .B1(n2435), .B2(
        div_output_EX_wire[16]), .C1(mul_output_EX_wire[16]), .C2(n2011), .ZN(
        n1230) );
  AOI222_X1 U1737 ( .A1(n2448), .A2(alu_output_EX_wire[26]), .B1(n2008), .B2(
        div_output_EX_wire[26]), .C1(mul_output_EX_wire[26]), .C2(n2011), .ZN(
        n1240) );
  NAND2_X1 U1738 ( .A1(n2007), .A2(N499), .ZN(n2346) );
  NAND2_X1 U1739 ( .A1(n2269), .A2(RF_source_2[20]), .ZN(n2345) );
  NAND2_X1 U1740 ( .A1(n2262), .A2(N403), .ZN(n2343) );
  NAND2_X1 U1741 ( .A1(n2424), .A2(RF_source_1[20]), .ZN(n2342) );
  AOI21_X1 U1742 ( .B1(mul_output_EX_wire[20]), .B2(n2011), .A(n2229), .ZN(
        n1234) );
  NAND2_X1 U1743 ( .A1(n2448), .A2(alu_output_EX_wire[20]), .ZN(n2231) );
  NAND2_X1 U1744 ( .A1(n2262), .A2(N388), .ZN(n2299) );
  NAND2_X1 U1745 ( .A1(n2423), .A2(RF_source_1[25]), .ZN(n2298) );
  NOR2_X1 U1746 ( .A1(n1494), .A2(funct3_EX_reg[2]), .ZN(n2503) );
  AND2_X1 U1747 ( .A1(n1562), .A2(funct7_EX_reg[0]), .ZN(n2478) );
  OR2_X1 U1748 ( .A1(n2418), .A2(n2169), .ZN(n2212) );
  OR2_X1 U1749 ( .A1(n2418), .A2(n2170), .ZN(n2213) );
  OR2_X1 U1750 ( .A1(n2418), .A2(n2172), .ZN(n2214) );
  OR2_X1 U1751 ( .A1(n2418), .A2(n2173), .ZN(n2215) );
  OR2_X1 U1752 ( .A1(n2418), .A2(n2177), .ZN(n2216) );
  OR2_X1 U1753 ( .A1(n2418), .A2(n2178), .ZN(n2217) );
  OR2_X1 U1754 ( .A1(n2418), .A2(n2179), .ZN(n2218) );
  OR2_X1 U1755 ( .A1(n2418), .A2(n2161), .ZN(n2219) );
  OR2_X1 U1756 ( .A1(n2418), .A2(n2162), .ZN(n2220) );
  OR2_X1 U1757 ( .A1(n2418), .A2(n2164), .ZN(n2221) );
  AND2_X1 U1758 ( .A1(n2419), .A2(pc_FD_reg[28]), .ZN(n2222) );
  NAND2_X1 U1759 ( .A1(next_pc_FD_wire[30]), .A2(n2496), .ZN(n2223) );
  NAND2_X1 U1760 ( .A1(n2223), .A2(n2224), .ZN(n1615) );
  NAND2_X1 U1761 ( .A1(next_pc_FD_wire[29]), .A2(n2496), .ZN(n2225) );
  NAND2_X1 U1762 ( .A1(n2225), .A2(n2226), .ZN(n1617) );
  NAND2_X1 U1763 ( .A1(next_pc_FD_wire[28]), .A2(n2496), .ZN(n2227) );
  NAND2_X1 U1764 ( .A1(n2227), .A2(n2228), .ZN(n1619) );
  AOI21_X1 U1765 ( .B1(n2093), .B2(n2421), .A(n2222), .ZN(n2228) );
  NAND2_X1 U1766 ( .A1(div_output_EX_wire[20]), .A2(n2008), .ZN(n2230) );
  NAND2_X1 U1767 ( .A1(n2230), .A2(n2231), .ZN(n2229) );
  NAND2_X1 U1768 ( .A1(div_output_EX_wire[21]), .A2(n2008), .ZN(n2233) );
  NAND2_X1 U1769 ( .A1(n2233), .A2(n2234), .ZN(n2232) );
  NAND2_X1 U1770 ( .A1(div_output_EX_wire[8]), .A2(n2435), .ZN(n2236) );
  NAND2_X1 U1771 ( .A1(n2236), .A2(n2237), .ZN(n2235) );
  NAND2_X1 U1772 ( .A1(div_output_EX_wire[11]), .A2(n2435), .ZN(n2239) );
  NAND2_X1 U1773 ( .A1(n2239), .A2(n2240), .ZN(n2238) );
  NAND2_X1 U1774 ( .A1(div_output_EX_wire[12]), .A2(n2435), .ZN(n2242) );
  NAND2_X1 U1775 ( .A1(n2242), .A2(n2243), .ZN(n2241) );
  NAND2_X1 U1776 ( .A1(div_output_EX_wire[14]), .A2(n2435), .ZN(n2245) );
  NAND2_X1 U1777 ( .A1(n2245), .A2(n2246), .ZN(n2244) );
  NAND2_X1 U1778 ( .A1(div_output_EX_wire[17]), .A2(n2008), .ZN(n2248) );
  NAND2_X1 U1779 ( .A1(n2248), .A2(n2249), .ZN(n2247) );
  OAI21_X1 U1780 ( .B1(n1214), .B2(n1488), .A(n2250), .ZN(\_2_net_[0] ) );
  OAI21_X1 U1781 ( .B1(n1215), .B2(n1488), .A(n2254), .ZN(\_2_net_[1] ) );
  OAI21_X1 U1782 ( .B1(n1216), .B2(n1488), .A(n2258), .ZN(\_2_net_[2] ) );
  AOI21_X1 U1783 ( .B1(FW_source_1[25]), .B2(n2422), .A(n2297), .ZN(n1408) );
  NAND2_X1 U1784 ( .A1(n2269), .A2(RF_source_2[30]), .ZN(n2264) );
  NAND2_X1 U1785 ( .A1(n2264), .A2(n2265), .ZN(n2263) );
  AOI21_X1 U1786 ( .B1(FW_source_2[30]), .B2(n2501), .A(n2263), .ZN(n1483) );
  AOI21_X1 U1787 ( .B1(FW_source_1[14]), .B2(n2500), .A(n2374), .ZN(n1386) );
  AOI21_X1 U1788 ( .B1(FW_source_1[15]), .B2(n2500), .A(n2380), .ZN(n1388) );
  AOI21_X1 U1789 ( .B1(FW_source_2[15]), .B2(n2501), .A(n2377), .ZN(n1453) );
  AOI21_X1 U1790 ( .B1(FW_source_1[16]), .B2(n2422), .A(n2303), .ZN(n1390) );
  AOI21_X1 U1791 ( .B1(FW_source_2[20]), .B2(n2501), .A(n2344), .ZN(n1463) );
  AOI21_X1 U1792 ( .B1(FW_source_1[18]), .B2(n2500), .A(n2359), .ZN(n1394) );
  AOI21_X1 U1793 ( .B1(FW_source_1[19]), .B2(n2500), .A(n2335), .ZN(n1396) );
  NAND2_X1 U1794 ( .A1(n2004), .A2(RF_source_2[0]), .ZN(n2271) );
  NAND2_X1 U1795 ( .A1(n2271), .A2(n2272), .ZN(n2270) );
  AOI21_X1 U1796 ( .B1(FW_source_2[0]), .B2(n2501), .A(n2270), .ZN(n1421) );
  NAND2_X1 U1797 ( .A1(n2268), .A2(RF_source_1[0]), .ZN(n2274) );
  NAND2_X1 U1798 ( .A1(n2274), .A2(n2275), .ZN(n2273) );
  AOI21_X1 U1799 ( .B1(FW_source_1[0]), .B2(n2500), .A(n2273), .ZN(n1356) );
  NAND2_X1 U1800 ( .A1(n2004), .A2(RF_source_2[1]), .ZN(n2277) );
  NAND2_X1 U1801 ( .A1(n2277), .A2(n2278), .ZN(n2276) );
  AOI21_X1 U1802 ( .B1(FW_source_2[1]), .B2(n2501), .A(n2276), .ZN(n1425) );
  NAND2_X1 U1803 ( .A1(n2424), .A2(RF_source_1[1]), .ZN(n2280) );
  NAND2_X1 U1804 ( .A1(n2280), .A2(n2281), .ZN(n2279) );
  AOI21_X1 U1805 ( .B1(FW_source_1[1]), .B2(n2500), .A(n2279), .ZN(n1360) );
  NAND2_X1 U1806 ( .A1(n2004), .A2(RF_source_2[2]), .ZN(n2283) );
  NAND2_X1 U1807 ( .A1(n2283), .A2(n2284), .ZN(n2282) );
  AOI21_X1 U1808 ( .B1(FW_source_2[2]), .B2(n2501), .A(n2282), .ZN(n1427) );
  NAND2_X1 U1809 ( .A1(n2423), .A2(RF_source_1[2]), .ZN(n2286) );
  NAND2_X1 U1810 ( .A1(n2286), .A2(n2287), .ZN(n2285) );
  AOI21_X1 U1811 ( .B1(FW_source_1[2]), .B2(n2500), .A(n2285), .ZN(n1362) );
  NAND2_X1 U1812 ( .A1(n2004), .A2(RF_source_2[3]), .ZN(n2289) );
  NAND2_X1 U1813 ( .A1(n2289), .A2(n2290), .ZN(n2288) );
  AOI21_X1 U1814 ( .B1(FW_source_2[3]), .B2(n2501), .A(n2288), .ZN(n1429) );
  AND2_X1 U1815 ( .A1(n2448), .A2(alu_output_EX_wire[25]), .ZN(n2291) );
  AOI21_X1 U1816 ( .B1(address_EX_wire[7]), .B2(n2479), .A(n2295), .ZN(n2294)
         );
  OAI21_X1 U1817 ( .B1(n1221), .B2(n1488), .A(n2294), .ZN(\_2_net_[7] ) );
  NAND2_X1 U1818 ( .A1(n2298), .A2(n2299), .ZN(n2297) );
  AOI21_X1 U1819 ( .B1(address_EX_wire[30]), .B2(n2479), .A(n2301), .ZN(n2300)
         );
  OAI21_X1 U1820 ( .B1(n1244), .B2(n1488), .A(n2300), .ZN(\_2_net_[30] ) );
  NAND2_X1 U1821 ( .A1(n2304), .A2(n2305), .ZN(n2303) );
  AOI21_X1 U1822 ( .B1(address_EX_wire[20]), .B2(n2479), .A(n2307), .ZN(n2306)
         );
  AOI21_X1 U1823 ( .B1(address_EX_wire[21]), .B2(n2479), .A(n2309), .ZN(n2308)
         );
  OAI21_X1 U1824 ( .B1(n1235), .B2(n1488), .A(n2308), .ZN(\_2_net_[21] ) );
  AOI21_X1 U1825 ( .B1(address_EX_wire[27]), .B2(n2479), .A(n2312), .ZN(n2311)
         );
  OAI21_X1 U1826 ( .B1(n1241), .B2(n1488), .A(n2311), .ZN(\_2_net_[27] ) );
  AOI21_X1 U1827 ( .B1(address_EX_wire[8]), .B2(n2479), .A(n2315), .ZN(n2314)
         );
  OAI21_X1 U1828 ( .B1(n1222), .B2(n1488), .A(n2314), .ZN(\_2_net_[8] ) );
  AOI21_X1 U1829 ( .B1(address_EX_wire[11]), .B2(n2479), .A(n2318), .ZN(n2317)
         );
  OAI21_X1 U1830 ( .B1(n1225), .B2(n1488), .A(n2317), .ZN(\_2_net_[11] ) );
  AOI21_X1 U1831 ( .B1(address_EX_wire[12]), .B2(n2479), .A(n2321), .ZN(n2320)
         );
  OAI21_X1 U1832 ( .B1(n1226), .B2(n1488), .A(n2320), .ZN(\_2_net_[12] ) );
  AND2_X1 U1833 ( .A1(div_output_EX_wire[18]), .A2(n2008), .ZN(n2323) );
  AOI21_X1 U1834 ( .B1(address_EX_wire[13]), .B2(n2479), .A(n2325), .ZN(n2324)
         );
  OAI21_X1 U1835 ( .B1(n1227), .B2(n1488), .A(n2324), .ZN(\_2_net_[13] ) );
  AOI21_X1 U1836 ( .B1(address_EX_wire[14]), .B2(n2479), .A(n2327), .ZN(n2326)
         );
  OAI21_X1 U1837 ( .B1(n1228), .B2(n1488), .A(n2326), .ZN(\_2_net_[14] ) );
  AOI21_X1 U1838 ( .B1(address_EX_wire[15]), .B2(n2479), .A(n2330), .ZN(n2329)
         );
  OAI21_X1 U1839 ( .B1(n1229), .B2(n1488), .A(n2329), .ZN(\_2_net_[15] ) );
  AOI21_X1 U1840 ( .B1(address_EX_wire[17]), .B2(n2479), .A(n2333), .ZN(n2332)
         );
  OAI21_X1 U1841 ( .B1(n1231), .B2(n1488), .A(n2332), .ZN(\_2_net_[17] ) );
  NAND2_X1 U1842 ( .A1(n2336), .A2(n2337), .ZN(n2335) );
  NAND2_X1 U1843 ( .A1(n2339), .A2(n2340), .ZN(n2338) );
  AOI21_X1 U1844 ( .B1(FW_source_1[30]), .B2(n2500), .A(n2338), .ZN(n1418) );
  NAND2_X1 U1845 ( .A1(n2342), .A2(n2343), .ZN(n2341) );
  AOI21_X1 U1846 ( .B1(FW_source_1[20]), .B2(n2422), .A(n2341), .ZN(n1398) );
  NAND2_X1 U1847 ( .A1(n2345), .A2(n2346), .ZN(n2344) );
  NAND2_X1 U1848 ( .A1(n2348), .A2(n2349), .ZN(n2347) );
  AOI21_X1 U1849 ( .B1(FW_source_1[21]), .B2(n2422), .A(n2347), .ZN(n1400) );
  NAND2_X1 U1850 ( .A1(n2351), .A2(n2352), .ZN(n2350) );
  AOI21_X1 U1851 ( .B1(FW_source_2[21]), .B2(n2425), .A(n2350), .ZN(n1465) );
  NAND2_X1 U1852 ( .A1(n2354), .A2(n2355), .ZN(n2353) );
  AOI21_X1 U1853 ( .B1(FW_source_1[27]), .B2(n2422), .A(n2353), .ZN(n1412) );
  NAND2_X1 U1854 ( .A1(n2357), .A2(n2358), .ZN(n2356) );
  AOI21_X1 U1855 ( .B1(FW_source_2[27]), .B2(n2425), .A(n2356), .ZN(n1477) );
  NAND2_X1 U1856 ( .A1(n2360), .A2(n2361), .ZN(n2359) );
  NAND2_X1 U1857 ( .A1(n2363), .A2(n2364), .ZN(n2362) );
  AOI21_X1 U1858 ( .B1(FW_source_1[10]), .B2(n2500), .A(n2362), .ZN(n1378) );
  NAND2_X1 U1859 ( .A1(n2366), .A2(n2367), .ZN(n2365) );
  AOI21_X1 U1860 ( .B1(FW_source_2[13]), .B2(n2501), .A(n2365), .ZN(n1449) );
  NAND2_X1 U1861 ( .A1(n2369), .A2(n2370), .ZN(n2368) );
  AOI21_X1 U1862 ( .B1(FW_source_1[13]), .B2(n2500), .A(n2368), .ZN(n1384) );
  NAND2_X1 U1863 ( .A1(n2372), .A2(n2373), .ZN(n2371) );
  AOI21_X1 U1864 ( .B1(FW_source_2[14]), .B2(n2501), .A(n2371), .ZN(n1451) );
  NAND2_X1 U1865 ( .A1(n2375), .A2(n2376), .ZN(n2374) );
  NAND2_X1 U1866 ( .A1(n2378), .A2(n2379), .ZN(n2377) );
  NAND2_X1 U1867 ( .A1(n2381), .A2(n2382), .ZN(n2380) );
  NAND2_X1 U1868 ( .A1(n2384), .A2(n2385), .ZN(n2383) );
  AOI21_X1 U1869 ( .B1(FW_source_2[17]), .B2(n2501), .A(n2383), .ZN(n1457) );
  NAND2_X1 U1870 ( .A1(n2387), .A2(n2388), .ZN(n2386) );
  AOI21_X1 U1871 ( .B1(FW_source_1[17]), .B2(n2500), .A(n2386), .ZN(n1392) );
  NAND2_X1 U1872 ( .A1(n2390), .A2(n2391), .ZN(n2389) );
  AOI21_X1 U1873 ( .B1(FW_source_2[8]), .B2(n2501), .A(n2389), .ZN(n1439) );
  NAND2_X1 U1874 ( .A1(n2393), .A2(n2394), .ZN(n2392) );
  AOI21_X1 U1875 ( .B1(FW_source_1[8]), .B2(n2500), .A(n2392), .ZN(n1374) );
  NAND2_X1 U1876 ( .A1(n2396), .A2(n2397), .ZN(n2395) );
  AOI21_X1 U1877 ( .B1(FW_source_2[12]), .B2(n2501), .A(n2395), .ZN(n1447) );
  NAND2_X1 U1878 ( .A1(n2399), .A2(n2400), .ZN(n2398) );
  AOI21_X1 U1879 ( .B1(FW_source_1[12]), .B2(n2500), .A(n2398), .ZN(n1382) );
  NAND2_X1 U1880 ( .A1(n2402), .A2(n2403), .ZN(n2401) );
  AOI21_X1 U1881 ( .B1(FW_source_2[7]), .B2(n2425), .A(n2401), .ZN(n1437) );
  NAND2_X1 U1882 ( .A1(n2405), .A2(n2406), .ZN(n2404) );
  AOI21_X1 U1883 ( .B1(FW_source_1[7]), .B2(n2422), .A(n2404), .ZN(n1372) );
  NAND2_X1 U1884 ( .A1(n2408), .A2(n2409), .ZN(n2407) );
  AOI21_X1 U1885 ( .B1(FW_source_2[11]), .B2(n2425), .A(n2407), .ZN(n1445) );
  NAND2_X1 U1886 ( .A1(n2411), .A2(n2412), .ZN(n2410) );
  AOI21_X1 U1887 ( .B1(FW_source_1[11]), .B2(n2422), .A(n2410), .ZN(n1380) );
  INV_X1 U1888 ( .A(n1319), .ZN(n1163) );
  NOR3_X1 U1889 ( .A1(n1559), .A2(n1168), .A3(n2154), .ZN(n2477) );
  INV_X1 U1890 ( .A(n1167), .ZN(n2415) );
  BUF_X1 U1891 ( .A(address_EX_wire[31]), .Z(n2416) );
  AOI222_X1 U1892 ( .A1(n2416), .A2(n2421), .B1(n2420), .B2(pc_FD_reg[31]), 
        .C1(n2496), .C2(next_pc_FD_wire[31]), .ZN(n2497) );
  INV_X1 U1893 ( .A(n2492), .ZN(n1639) );
  INV_X1 U1894 ( .A(n2485), .ZN(n1623) );
  INV_X1 U1895 ( .A(n2491), .ZN(n1635) );
  INV_X1 U1896 ( .A(n2488), .ZN(n1629) );
  INV_X1 U1897 ( .A(n2484), .ZN(n1621) );
  AOI222_X1 U1898 ( .A1(n2006), .A2(address_EX_wire[18]), .B1(n2420), .B2(
        pc_FD_reg[18]), .C1(n2496), .C2(next_pc_FD_wire[18]), .ZN(n2492) );
  INV_X1 U1899 ( .A(n2489), .ZN(n1631) );
  AOI222_X1 U1900 ( .A1(n2006), .A2(n2099), .B1(n2419), .B2(pc_FD_reg[22]), 
        .C1(n2496), .C2(next_pc_FD_wire[22]), .ZN(n2489) );
  AOI222_X1 U1901 ( .A1(n2006), .A2(address_EX_wire[26]), .B1(n2419), .B2(
        pc_FD_reg[26]), .C1(n2496), .C2(next_pc_FD_wire[26]), .ZN(n2485) );
  INV_X1 U1902 ( .A(n2490), .ZN(n1633) );
  AOI222_X1 U1903 ( .A1(n2006), .A2(n2092), .B1(n2419), .B2(pc_FD_reg[21]), 
        .C1(n2496), .C2(next_pc_FD_wire[21]), .ZN(n2490) );
  AOI222_X1 U1904 ( .A1(n2006), .A2(n2098), .B1(n2419), .B2(pc_FD_reg[23]), 
        .C1(n2496), .C2(next_pc_FD_wire[23]), .ZN(n2488) );
  INV_X1 U1905 ( .A(n2486), .ZN(n1625) );
  AOI222_X1 U1906 ( .A1(n2006), .A2(n2086), .B1(n2419), .B2(pc_FD_reg[25]), 
        .C1(n2496), .C2(next_pc_FD_wire[25]), .ZN(n2486) );
  AOI222_X1 U1907 ( .A1(n2006), .A2(address_EX_wire[27]), .B1(n2419), .B2(
        pc_FD_reg[27]), .C1(n2496), .C2(next_pc_FD_wire[27]), .ZN(n2484) );
  AOI222_X1 U1908 ( .A1(n2006), .A2(address_EX_wire[20]), .B1(n2419), .B2(
        pc_FD_reg[20]), .C1(n2496), .C2(next_pc_FD_wire[20]), .ZN(n2491) );
  INV_X1 U1909 ( .A(n2495), .ZN(n1659) );
  INV_X1 U1910 ( .A(n2494), .ZN(n1657) );
  AOI222_X1 U1911 ( .A1(n2421), .A2(address_EX_wire[9]), .B1(n2420), .B2(
        pc_FD_reg[9]), .C1(n2496), .C2(next_pc_FD_wire[9]), .ZN(n2494) );
  AOI222_X1 U1912 ( .A1(n2421), .A2(address_EX_wire[8]), .B1(n2420), .B2(
        pc_FD_reg[8]), .C1(n2496), .C2(next_pc_FD_wire[8]), .ZN(n2495) );
  INV_X1 U1913 ( .A(n2497), .ZN(n1613) );
  INV_X1 U1914 ( .A(n2493), .ZN(n1651) );
  AOI222_X1 U1915 ( .A1(n2421), .A2(address_EX_wire[12]), .B1(n2420), .B2(
        pc_FD_reg[12]), .C1(n2496), .C2(next_pc_FD_wire[12]), .ZN(n2493) );
  INV_X1 U1916 ( .A(n2487), .ZN(n1627) );
  OR2_X1 U1917 ( .A1(n1354), .A2(reset), .ZN(n2417) );
  NOR2_X1 U1918 ( .A1(n1354), .A2(reset), .ZN(_0_net_) );
  INV_X1 U1919 ( .A(n2056), .ZN(n2454) );
  NAND3_X1 U1920 ( .A1(n1563), .A2(n1561), .A3(n2478), .ZN(n1494) );
  MUX2_X1 U1921 ( .A(n2416), .B(address_MW_reg[31]), .S(n2437), .Z(n887) );
  MUX2_X1 U1922 ( .A(address_EX_wire[30]), .B(address_MW_reg[30]), .S(n2437), 
        .Z(n888) );
  MUX2_X1 U1923 ( .A(address_EX_wire[29]), .B(address_MW_reg[29]), .S(n2437), 
        .Z(n889) );
  MUX2_X1 U1924 ( .A(n2093), .B(address_MW_reg[28]), .S(n2437), .Z(n890) );
  MUX2_X1 U1925 ( .A(address_EX_wire[27]), .B(address_MW_reg[27]), .S(n2437), 
        .Z(n891) );
  MUX2_X1 U1926 ( .A(address_EX_wire[26]), .B(address_MW_reg[26]), .S(n2437), 
        .Z(n892) );
  MUX2_X1 U1927 ( .A(n2086), .B(address_MW_reg[25]), .S(n2437), .Z(n893) );
  MUX2_X1 U1928 ( .A(n2097), .B(address_MW_reg[24]), .S(n2437), .Z(n894) );
  MUX2_X1 U1929 ( .A(n2098), .B(address_MW_reg[23]), .S(n2437), .Z(n895) );
  MUX2_X1 U1930 ( .A(n2099), .B(address_MW_reg[22]), .S(n2437), .Z(n896) );
  MUX2_X1 U1931 ( .A(n2092), .B(address_MW_reg[21]), .S(n2437), .Z(n897) );
  MUX2_X1 U1932 ( .A(address_EX_wire[20]), .B(address_MW_reg[20]), .S(n2438), 
        .Z(n898) );
  MUX2_X1 U1933 ( .A(n2090), .B(address_MW_reg[19]), .S(n2438), .Z(n899) );
  MUX2_X1 U1934 ( .A(address_EX_wire[18]), .B(address_MW_reg[18]), .S(n2438), 
        .Z(n900) );
  MUX2_X1 U1935 ( .A(address_EX_wire[17]), .B(address_MW_reg[17]), .S(n2438), 
        .Z(n901) );
  MUX2_X1 U1936 ( .A(n2010), .B(address_MW_reg[16]), .S(n2438), .Z(n902) );
  MUX2_X1 U1937 ( .A(address_EX_wire[15]), .B(address_MW_reg[15]), .S(n2438), 
        .Z(n903) );
  MUX2_X1 U1938 ( .A(address_EX_wire[14]), .B(address_MW_reg[14]), .S(n2438), 
        .Z(n904) );
  MUX2_X1 U1939 ( .A(address_EX_wire[13]), .B(address_MW_reg[13]), .S(n2438), 
        .Z(n905) );
  MUX2_X1 U1940 ( .A(address_EX_wire[12]), .B(address_MW_reg[12]), .S(n2438), 
        .Z(n906) );
  MUX2_X1 U1941 ( .A(address_EX_wire[11]), .B(address_MW_reg[11]), .S(n2438), 
        .Z(n907) );
  MUX2_X1 U1942 ( .A(address_EX_wire[10]), .B(address_MW_reg[10]), .S(n2438), 
        .Z(n908) );
  MUX2_X1 U1943 ( .A(address_EX_wire[9]), .B(address_MW_reg[9]), .S(n2438), 
        .Z(n909) );
  MUX2_X1 U1944 ( .A(address_EX_wire[8]), .B(address_MW_reg[8]), .S(n2439), 
        .Z(n910) );
endmodule

